VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top_dac_adc
  CLASS BLOCK ;
  FOREIGN top_dac_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.048500 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 256.000000 ;
    ANTENNADIFFAREA 4.850000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.444000 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN VGND
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1622.984985 ;
    ANTENNADIFFAREA 901.023560 ;
    PORT
      LAYER met4 ;
        RECT 35.920 5.050 37.920 7.050 ;
    END
  END VGND
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1026.025024 ;
    ANTENNADIFFAREA 1187.786011 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1026.025024 ;
    ANTENNADIFFAREA 1187.786011 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1026.025024 ;
    ANTENNADIFFAREA 1187.786011 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1026.025024 ;
    ANTENNADIFFAREA 1187.786011 ;
    PORT
      LAYER met4 ;
        RECT 32.560 5.050 34.560 7.050 ;
    END
  END VDPWR
  OBS
      LAYER nwell ;
        RECT 17.080 219.855 147.180 221.460 ;
      LAYER pwell ;
        RECT 17.275 218.655 18.645 219.465 ;
        RECT 18.655 218.655 24.165 219.465 ;
        RECT 24.175 218.655 29.685 219.465 ;
        RECT 30.165 218.740 30.595 219.525 ;
        RECT 30.615 218.655 36.125 219.465 ;
        RECT 36.135 218.655 41.645 219.465 ;
        RECT 41.655 218.655 43.025 219.465 ;
        RECT 43.045 218.740 43.475 219.525 ;
        RECT 43.495 218.655 49.005 219.465 ;
        RECT 49.015 218.655 54.525 219.465 ;
        RECT 54.535 218.655 55.905 219.465 ;
        RECT 55.925 218.740 56.355 219.525 ;
        RECT 56.375 218.655 60.045 219.465 ;
        RECT 60.515 218.655 63.125 219.565 ;
        RECT 63.275 218.655 68.785 219.465 ;
        RECT 68.805 218.740 69.235 219.525 ;
        RECT 69.255 218.655 74.765 219.465 ;
        RECT 74.775 218.655 78.445 219.465 ;
        RECT 78.455 218.655 79.825 219.465 ;
        RECT 79.835 219.335 81.180 219.565 ;
        RECT 79.835 218.655 81.665 219.335 ;
        RECT 81.685 218.740 82.115 219.525 ;
        RECT 85.555 219.475 86.505 219.565 ;
        RECT 83.055 218.655 84.425 219.435 ;
        RECT 85.555 218.655 87.485 219.475 ;
        RECT 87.655 218.655 89.025 219.435 ;
        RECT 89.035 218.655 90.405 219.465 ;
        RECT 90.425 218.655 91.775 219.565 ;
        RECT 91.795 218.655 94.545 219.465 ;
        RECT 94.565 218.740 94.995 219.525 ;
        RECT 95.935 219.335 97.280 219.565 ;
        RECT 95.935 218.655 97.765 219.335 ;
        RECT 97.775 218.655 103.285 219.465 ;
        RECT 103.295 218.655 106.965 219.465 ;
        RECT 107.445 218.740 107.875 219.525 ;
        RECT 107.895 218.655 113.405 219.465 ;
        RECT 113.415 218.655 118.925 219.465 ;
        RECT 118.935 218.655 120.305 219.465 ;
        RECT 120.325 218.740 120.755 219.525 ;
        RECT 120.775 218.655 126.285 219.465 ;
        RECT 126.295 218.655 131.805 219.465 ;
        RECT 131.815 218.655 133.185 219.465 ;
        RECT 133.205 218.740 133.635 219.525 ;
        RECT 133.655 218.655 139.165 219.465 ;
        RECT 139.175 218.655 144.685 219.465 ;
        RECT 145.615 218.655 146.985 219.465 ;
        RECT 17.415 218.445 17.585 218.655 ;
        RECT 18.795 218.445 18.965 218.655 ;
        RECT 24.315 218.445 24.485 218.655 ;
        RECT 29.835 218.605 30.005 218.635 ;
        RECT 29.830 218.495 30.005 218.605 ;
        RECT 29.835 218.445 30.005 218.495 ;
        RECT 30.755 218.465 30.925 218.655 ;
        RECT 35.355 218.445 35.525 218.635 ;
        RECT 36.275 218.465 36.445 218.655 ;
        RECT 40.875 218.445 41.045 218.635 ;
        RECT 41.795 218.465 41.965 218.655 ;
        RECT 42.710 218.495 42.830 218.605 ;
        RECT 43.635 218.445 43.805 218.655 ;
        RECT 49.155 218.445 49.325 218.655 ;
        RECT 51.910 218.495 52.030 218.605 ;
        RECT 53.750 218.445 53.920 218.635 ;
        RECT 54.675 218.465 54.845 218.655 ;
        RECT 55.590 218.445 55.760 218.635 ;
        RECT 56.065 218.490 56.225 218.600 ;
        RECT 56.515 218.465 56.685 218.655 ;
        RECT 56.975 218.445 57.145 218.635 ;
        RECT 60.190 218.495 60.310 218.605 ;
        RECT 60.660 218.445 60.830 218.655 ;
        RECT 62.035 218.445 62.205 218.635 ;
        RECT 63.415 218.465 63.585 218.655 ;
        RECT 69.395 218.635 69.565 218.655 ;
        RECT 65.715 218.445 65.885 218.635 ;
        RECT 68.475 218.445 68.645 218.635 ;
        RECT 69.395 218.465 69.570 218.635 ;
        RECT 69.400 218.445 69.570 218.465 ;
        RECT 70.775 218.445 70.945 218.635 ;
        RECT 74.915 218.465 75.085 218.655 ;
        RECT 76.295 218.445 76.465 218.635 ;
        RECT 78.595 218.465 78.765 218.655 ;
        RECT 79.985 218.490 80.145 218.600 ;
        RECT 80.895 218.445 81.065 218.635 ;
        RECT 81.355 218.465 81.525 218.655 ;
        RECT 82.285 218.500 82.445 218.610 ;
        RECT 83.205 218.465 83.375 218.655 ;
        RECT 87.335 218.635 87.485 218.655 ;
        RECT 84.575 218.445 84.745 218.635 ;
        RECT 85.955 218.445 86.125 218.635 ;
        RECT 87.335 218.465 87.505 218.635 ;
        RECT 87.805 218.465 87.975 218.655 ;
        RECT 89.175 218.465 89.345 218.655 ;
        RECT 89.640 218.445 89.810 218.635 ;
        RECT 90.555 218.465 90.725 218.655 ;
        RECT 91.935 218.465 92.105 218.655 ;
        RECT 92.850 218.495 92.970 218.605 ;
        RECT 93.310 218.445 93.480 218.635 ;
        RECT 17.275 217.635 18.645 218.445 ;
        RECT 18.655 217.635 24.165 218.445 ;
        RECT 24.175 217.635 29.685 218.445 ;
        RECT 29.695 217.635 35.205 218.445 ;
        RECT 35.215 217.635 40.725 218.445 ;
        RECT 40.735 217.635 42.565 218.445 ;
        RECT 43.045 217.575 43.475 218.360 ;
        RECT 43.495 217.635 49.005 218.445 ;
        RECT 49.015 217.635 51.765 218.445 ;
        RECT 52.295 217.535 54.065 218.445 ;
        RECT 54.135 217.535 55.905 218.445 ;
        RECT 56.945 217.765 60.410 218.445 ;
        RECT 59.490 217.535 60.410 217.765 ;
        RECT 60.515 217.535 61.865 218.445 ;
        RECT 61.895 217.635 65.565 218.445 ;
        RECT 65.575 217.635 66.945 218.445 ;
        RECT 66.955 217.535 68.770 218.445 ;
        RECT 68.805 217.575 69.235 218.360 ;
        RECT 69.255 217.535 70.605 218.445 ;
        RECT 70.635 217.635 76.145 218.445 ;
        RECT 76.155 217.635 79.825 218.445 ;
        RECT 80.865 217.765 84.330 218.445 ;
        RECT 83.410 217.535 84.330 217.765 ;
        RECT 84.435 217.635 85.805 218.445 ;
        RECT 85.925 217.765 89.390 218.445 ;
        RECT 88.470 217.535 89.390 217.765 ;
        RECT 89.495 217.535 92.415 218.445 ;
        RECT 93.195 217.535 94.545 218.445 ;
        RECT 95.160 218.415 95.330 218.635 ;
        RECT 97.455 218.465 97.625 218.655 ;
        RECT 97.915 218.465 98.085 218.655 ;
        RECT 98.385 218.490 98.545 218.600 ;
        RECT 99.295 218.445 99.465 218.635 ;
        RECT 102.515 218.465 102.685 218.635 ;
        RECT 103.435 218.465 103.605 218.655 ;
        RECT 102.520 218.445 102.685 218.465 ;
        RECT 104.815 218.445 104.985 218.635 ;
        RECT 107.110 218.495 107.230 218.605 ;
        RECT 108.035 218.465 108.205 218.655 ;
        RECT 110.335 218.445 110.505 218.635 ;
        RECT 113.555 218.465 113.725 218.655 ;
        RECT 115.855 218.445 116.025 218.635 ;
        RECT 119.075 218.465 119.245 218.655 ;
        RECT 119.545 218.490 119.705 218.600 ;
        RECT 120.915 218.445 121.085 218.655 ;
        RECT 126.435 218.445 126.605 218.655 ;
        RECT 131.955 218.445 132.125 218.655 ;
        RECT 133.795 218.465 133.965 218.655 ;
        RECT 137.475 218.445 137.645 218.635 ;
        RECT 139.315 218.465 139.485 218.655 ;
        RECT 142.995 218.445 143.165 218.635 ;
        RECT 144.845 218.500 145.005 218.610 ;
        RECT 146.675 218.445 146.845 218.655 ;
        RECT 97.290 218.415 98.225 218.445 ;
        RECT 94.565 217.575 94.995 218.360 ;
        RECT 95.160 218.215 98.225 218.415 ;
        RECT 95.015 217.735 98.225 218.215 ;
        RECT 95.015 217.535 95.945 217.735 ;
        RECT 97.275 217.535 98.225 217.735 ;
        RECT 99.255 217.535 102.365 218.445 ;
        RECT 102.520 217.765 104.355 218.445 ;
        RECT 103.425 217.535 104.355 217.765 ;
        RECT 104.675 217.635 110.185 218.445 ;
        RECT 110.195 217.635 115.705 218.445 ;
        RECT 115.715 217.635 119.385 218.445 ;
        RECT 120.325 217.575 120.755 218.360 ;
        RECT 120.775 217.635 126.285 218.445 ;
        RECT 126.295 217.635 131.805 218.445 ;
        RECT 131.815 217.635 137.325 218.445 ;
        RECT 137.335 217.635 142.845 218.445 ;
        RECT 142.855 217.635 145.605 218.445 ;
        RECT 145.615 217.635 146.985 218.445 ;
      LAYER nwell ;
        RECT 17.080 214.415 147.180 217.245 ;
      LAYER pwell ;
        RECT 17.275 213.215 18.645 214.025 ;
        RECT 18.655 213.215 24.165 214.025 ;
        RECT 24.175 213.215 29.685 214.025 ;
        RECT 30.165 213.300 30.595 214.085 ;
        RECT 30.615 213.215 36.125 214.025 ;
        RECT 36.135 213.215 41.645 214.025 ;
        RECT 41.655 213.215 47.165 214.025 ;
        RECT 47.175 213.215 49.005 214.025 ;
        RECT 49.110 213.895 50.030 214.125 ;
        RECT 49.110 213.215 52.575 213.895 ;
        RECT 52.695 213.215 55.805 214.125 ;
        RECT 55.925 213.300 56.355 214.085 ;
        RECT 56.415 213.895 57.765 214.125 ;
        RECT 59.300 213.895 60.210 214.115 ;
        RECT 64.235 213.895 65.585 214.125 ;
        RECT 67.120 213.895 68.030 214.115 ;
        RECT 56.415 213.215 63.725 213.895 ;
        RECT 64.235 213.215 71.545 213.895 ;
        RECT 71.555 213.215 77.065 214.025 ;
        RECT 77.075 213.215 80.745 214.025 ;
        RECT 81.685 213.300 82.115 214.085 ;
        RECT 82.635 213.895 83.985 214.125 ;
        RECT 85.520 213.895 86.430 214.115 ;
        RECT 93.470 213.895 94.380 214.115 ;
        RECT 95.915 213.895 97.265 214.125 ;
        RECT 100.830 213.895 101.740 214.115 ;
        RECT 103.275 213.895 104.625 214.125 ;
        RECT 82.635 213.215 89.945 213.895 ;
        RECT 89.955 213.215 97.265 213.895 ;
        RECT 97.315 213.215 104.625 213.895 ;
        RECT 104.685 213.215 107.425 213.895 ;
        RECT 107.445 213.300 107.875 214.085 ;
        RECT 107.895 213.215 113.405 214.025 ;
        RECT 113.415 213.215 118.925 214.025 ;
        RECT 118.935 213.215 124.445 214.025 ;
        RECT 124.455 213.215 129.965 214.025 ;
        RECT 129.975 213.215 132.725 214.025 ;
        RECT 133.205 213.300 133.635 214.085 ;
        RECT 133.655 213.215 139.165 214.025 ;
        RECT 139.175 213.215 144.685 214.025 ;
        RECT 145.615 213.215 146.985 214.025 ;
        RECT 17.415 213.005 17.585 213.215 ;
        RECT 18.795 213.005 18.965 213.215 ;
        RECT 24.315 213.005 24.485 213.215 ;
        RECT 29.835 213.165 30.005 213.195 ;
        RECT 29.830 213.055 30.005 213.165 ;
        RECT 29.835 213.005 30.005 213.055 ;
        RECT 30.755 213.025 30.925 213.215 ;
        RECT 35.355 213.005 35.525 213.195 ;
        RECT 36.275 213.025 36.445 213.215 ;
        RECT 40.875 213.005 41.045 213.195 ;
        RECT 41.795 213.025 41.965 213.215 ;
        RECT 42.710 213.055 42.830 213.165 ;
        RECT 43.635 213.005 43.805 213.195 ;
        RECT 45.930 213.005 46.100 213.195 ;
        RECT 46.395 213.005 46.565 213.195 ;
        RECT 47.315 213.025 47.485 213.215 ;
        RECT 52.375 213.025 52.545 213.215 ;
        RECT 53.755 213.005 53.925 213.195 ;
        RECT 55.595 213.025 55.765 213.215 ;
        RECT 63.415 213.025 63.585 213.215 ;
        RECT 63.870 213.055 63.990 213.165 ;
        RECT 64.335 213.005 64.505 213.195 ;
        RECT 64.790 213.055 64.910 213.165 ;
        RECT 65.255 213.005 65.425 213.195 ;
        RECT 71.235 213.025 71.405 213.215 ;
        RECT 71.695 213.025 71.865 213.215 ;
        RECT 72.615 213.005 72.785 213.195 ;
        RECT 73.075 213.005 73.245 213.195 ;
        RECT 77.215 213.025 77.385 213.215 ;
        RECT 80.435 213.005 80.605 213.195 ;
        RECT 80.905 213.060 81.065 213.170 ;
        RECT 82.270 213.055 82.390 213.165 ;
        RECT 87.805 213.050 87.965 213.160 ;
        RECT 88.720 213.005 88.890 213.195 ;
        RECT 89.635 213.025 89.805 213.215 ;
        RECT 90.095 213.025 90.265 213.215 ;
        RECT 97.455 213.195 97.625 213.215 ;
        RECT 93.315 213.005 93.485 213.195 ;
        RECT 93.785 213.050 93.945 213.160 ;
        RECT 17.275 212.195 18.645 213.005 ;
        RECT 18.655 212.195 24.165 213.005 ;
        RECT 24.175 212.195 29.685 213.005 ;
        RECT 29.695 212.195 35.205 213.005 ;
        RECT 35.215 212.195 40.725 213.005 ;
        RECT 40.735 212.195 42.565 213.005 ;
        RECT 43.045 212.135 43.475 212.920 ;
        RECT 43.495 212.195 44.865 213.005 ;
        RECT 44.895 212.095 46.245 213.005 ;
        RECT 46.255 212.325 53.565 213.005 ;
        RECT 53.615 212.325 60.925 213.005 ;
        RECT 49.770 212.105 50.680 212.325 ;
        RECT 52.215 212.095 53.565 212.325 ;
        RECT 57.130 212.105 58.040 212.325 ;
        RECT 59.575 212.095 60.925 212.325 ;
        RECT 61.070 212.325 64.535 213.005 ;
        RECT 65.225 212.325 68.690 213.005 ;
        RECT 61.070 212.095 61.990 212.325 ;
        RECT 67.770 212.095 68.690 212.325 ;
        RECT 68.805 212.135 69.235 212.920 ;
        RECT 69.395 212.095 72.845 213.005 ;
        RECT 72.935 212.325 80.245 213.005 ;
        RECT 80.295 212.325 87.605 213.005 ;
        RECT 76.450 212.105 77.360 212.325 ;
        RECT 78.895 212.095 80.245 212.325 ;
        RECT 83.810 212.105 84.720 212.325 ;
        RECT 86.255 212.095 87.605 212.325 ;
        RECT 88.575 212.095 92.230 213.005 ;
        RECT 92.265 212.095 93.615 213.005 ;
        RECT 95.150 212.975 95.320 213.195 ;
        RECT 97.455 213.025 97.630 213.195 ;
        RECT 107.115 213.025 107.285 213.215 ;
        RECT 97.460 213.005 97.630 213.025 ;
        RECT 108.035 213.005 108.205 213.215 ;
        RECT 108.495 213.005 108.665 213.195 ;
        RECT 113.555 213.025 113.725 213.215 ;
        RECT 114.015 213.005 114.185 213.195 ;
        RECT 119.075 213.025 119.245 213.215 ;
        RECT 119.545 213.050 119.705 213.160 ;
        RECT 120.915 213.005 121.085 213.195 ;
        RECT 124.595 213.025 124.765 213.215 ;
        RECT 126.435 213.005 126.605 213.195 ;
        RECT 130.115 213.025 130.285 213.215 ;
        RECT 131.955 213.005 132.125 213.195 ;
        RECT 132.870 213.055 132.990 213.165 ;
        RECT 133.795 213.025 133.965 213.215 ;
        RECT 137.475 213.005 137.645 213.195 ;
        RECT 139.315 213.025 139.485 213.215 ;
        RECT 142.995 213.005 143.165 213.195 ;
        RECT 144.845 213.060 145.005 213.170 ;
        RECT 146.675 213.005 146.845 213.215 ;
        RECT 96.350 212.975 97.305 213.005 ;
        RECT 94.565 212.135 94.995 212.920 ;
        RECT 95.025 212.295 97.305 212.975 ;
        RECT 96.350 212.095 97.305 212.295 ;
        RECT 97.315 212.325 100.900 213.005 ;
        RECT 101.035 212.325 108.345 213.005 ;
        RECT 97.315 212.095 98.235 212.325 ;
        RECT 101.035 212.095 102.385 212.325 ;
        RECT 103.920 212.105 104.830 212.325 ;
        RECT 108.355 212.195 113.865 213.005 ;
        RECT 113.875 212.195 119.385 213.005 ;
        RECT 120.325 212.135 120.755 212.920 ;
        RECT 120.775 212.195 126.285 213.005 ;
        RECT 126.295 212.195 131.805 213.005 ;
        RECT 131.815 212.195 137.325 213.005 ;
        RECT 137.335 212.195 142.845 213.005 ;
        RECT 142.855 212.195 145.605 213.005 ;
        RECT 145.615 212.195 146.985 213.005 ;
      LAYER nwell ;
        RECT 17.080 208.975 147.180 211.805 ;
      LAYER pwell ;
        RECT 17.275 207.775 18.645 208.585 ;
        RECT 18.655 207.775 24.165 208.585 ;
        RECT 24.175 207.775 29.685 208.585 ;
        RECT 30.165 207.860 30.595 208.645 ;
        RECT 30.615 207.775 36.125 208.585 ;
        RECT 36.135 207.775 41.645 208.585 ;
        RECT 41.655 207.775 45.325 208.585 ;
        RECT 49.310 208.455 50.220 208.675 ;
        RECT 51.755 208.455 53.105 208.685 ;
        RECT 45.795 207.775 53.105 208.455 ;
        RECT 54.075 207.775 55.890 208.685 ;
        RECT 55.925 207.860 56.355 208.645 ;
        RECT 58.450 208.455 59.585 208.685 ;
        RECT 56.375 207.775 59.585 208.455 ;
        RECT 60.055 208.455 60.975 208.685 ;
        RECT 60.055 207.775 62.345 208.455 ;
        RECT 62.455 207.775 65.565 208.685 ;
        RECT 69.090 208.455 70.000 208.675 ;
        RECT 71.535 208.455 72.885 208.685 ;
        RECT 74.270 208.485 75.225 208.685 ;
        RECT 65.575 207.775 72.885 208.455 ;
        RECT 72.945 207.805 75.225 208.485 ;
        RECT 17.415 207.565 17.585 207.775 ;
        RECT 18.795 207.565 18.965 207.775 ;
        RECT 24.315 207.565 24.485 207.775 ;
        RECT 29.835 207.725 30.005 207.755 ;
        RECT 29.830 207.615 30.005 207.725 ;
        RECT 29.835 207.565 30.005 207.615 ;
        RECT 30.755 207.585 30.925 207.775 ;
        RECT 35.355 207.565 35.525 207.755 ;
        RECT 36.275 207.585 36.445 207.775 ;
        RECT 40.875 207.565 41.045 207.755 ;
        RECT 41.795 207.585 41.965 207.775 ;
        RECT 42.710 207.615 42.830 207.725 ;
        RECT 43.635 207.565 43.805 207.755 ;
        RECT 45.470 207.615 45.590 207.725 ;
        RECT 45.935 207.585 46.105 207.775 ;
        RECT 49.155 207.565 49.325 207.755 ;
        RECT 50.540 207.565 50.710 207.755 ;
        RECT 51.915 207.565 52.085 207.755 ;
        RECT 53.305 207.620 53.465 207.730 ;
        RECT 54.670 207.615 54.790 207.725 ;
        RECT 55.595 207.585 55.765 207.775 ;
        RECT 56.055 207.565 56.225 207.755 ;
        RECT 56.515 207.565 56.685 207.775 ;
        RECT 59.730 207.615 59.850 207.725 ;
        RECT 62.035 207.565 62.205 207.775 ;
        RECT 62.495 207.585 62.665 207.775 ;
        RECT 65.250 207.565 65.420 207.755 ;
        RECT 65.715 207.585 65.885 207.775 ;
        RECT 68.475 207.565 68.645 207.755 ;
        RECT 70.775 207.565 70.945 207.755 ;
        RECT 71.235 207.565 71.405 207.755 ;
        RECT 73.070 207.585 73.240 207.805 ;
        RECT 74.270 207.775 75.225 207.805 ;
        RECT 75.235 207.775 80.745 208.585 ;
        RECT 81.685 207.860 82.115 208.645 ;
        RECT 82.595 208.455 85.420 208.685 ;
        RECT 86.370 208.455 87.290 208.685 ;
        RECT 89.955 208.485 90.900 208.685 ;
        RECT 92.235 208.485 93.165 208.685 ;
        RECT 82.595 207.775 86.125 208.455 ;
        RECT 86.370 207.775 89.835 208.455 ;
        RECT 89.955 208.005 93.165 208.485 ;
        RECT 94.225 208.455 95.155 208.685 ;
        RECT 89.955 207.805 93.025 208.005 ;
        RECT 89.955 207.775 90.900 207.805 ;
        RECT 75.375 207.585 75.545 207.775 ;
        RECT 85.925 207.755 86.125 207.775 ;
        RECT 76.755 207.565 76.925 207.755 ;
        RECT 80.905 207.620 81.065 207.730 ;
        RECT 82.275 207.725 82.445 207.755 ;
        RECT 82.270 207.615 82.445 207.725 ;
        RECT 85.030 207.615 85.150 207.725 ;
        RECT 82.275 207.565 82.445 207.615 ;
        RECT 85.495 207.565 85.665 207.755 ;
        RECT 85.955 207.585 86.125 207.755 ;
        RECT 88.255 207.565 88.425 207.755 ;
        RECT 89.635 207.585 89.805 207.775 ;
        RECT 92.855 207.585 93.025 207.805 ;
        RECT 93.320 207.775 95.155 208.455 ;
        RECT 95.475 207.775 97.305 208.585 ;
        RECT 97.315 207.775 100.975 208.685 ;
        RECT 100.995 207.775 106.505 208.585 ;
        RECT 107.445 207.860 107.875 208.645 ;
        RECT 107.895 207.775 113.405 208.585 ;
        RECT 113.415 207.775 118.925 208.585 ;
        RECT 118.935 207.775 124.445 208.585 ;
        RECT 124.455 207.775 129.965 208.585 ;
        RECT 129.975 207.775 132.725 208.585 ;
        RECT 133.205 207.860 133.635 208.645 ;
        RECT 133.655 207.775 139.165 208.585 ;
        RECT 139.175 207.775 144.685 208.585 ;
        RECT 145.615 207.775 146.985 208.585 ;
        RECT 93.320 207.755 93.485 207.775 ;
        RECT 93.315 207.585 93.485 207.755 ;
        RECT 93.785 207.610 93.945 207.720 ;
        RECT 95.160 207.565 95.330 207.755 ;
        RECT 95.615 207.585 95.785 207.775 ;
        RECT 96.535 207.565 96.705 207.755 ;
        RECT 100.680 207.585 100.850 207.775 ;
        RECT 101.135 207.585 101.305 207.775 ;
        RECT 102.055 207.565 102.225 207.755 ;
        RECT 106.665 207.620 106.825 207.730 ;
        RECT 107.575 207.565 107.745 207.755 ;
        RECT 108.035 207.585 108.205 207.775 ;
        RECT 110.330 207.615 110.450 207.725 ;
        RECT 110.795 207.565 110.965 207.755 ;
        RECT 113.555 207.585 113.725 207.775 ;
        RECT 114.475 207.565 114.645 207.755 ;
        RECT 119.075 207.585 119.245 207.775 ;
        RECT 119.990 207.615 120.110 207.725 ;
        RECT 120.915 207.565 121.085 207.755 ;
        RECT 124.595 207.585 124.765 207.775 ;
        RECT 126.435 207.565 126.605 207.755 ;
        RECT 130.115 207.585 130.285 207.775 ;
        RECT 131.955 207.565 132.125 207.755 ;
        RECT 132.870 207.615 132.990 207.725 ;
        RECT 133.795 207.585 133.965 207.775 ;
        RECT 137.475 207.565 137.645 207.755 ;
        RECT 139.315 207.585 139.485 207.775 ;
        RECT 142.995 207.565 143.165 207.755 ;
        RECT 144.845 207.620 145.005 207.730 ;
        RECT 146.675 207.565 146.845 207.775 ;
        RECT 17.275 206.755 18.645 207.565 ;
        RECT 18.655 206.755 24.165 207.565 ;
        RECT 24.175 206.755 29.685 207.565 ;
        RECT 29.695 206.755 35.205 207.565 ;
        RECT 35.215 206.755 40.725 207.565 ;
        RECT 40.735 206.755 42.565 207.565 ;
        RECT 43.045 206.695 43.475 207.480 ;
        RECT 43.495 206.755 49.005 207.565 ;
        RECT 49.015 206.755 50.385 207.565 ;
        RECT 50.395 206.655 51.745 207.565 ;
        RECT 51.775 206.755 54.525 207.565 ;
        RECT 55.005 206.655 56.355 207.565 ;
        RECT 56.375 206.755 61.885 207.565 ;
        RECT 61.895 206.755 63.725 207.565 ;
        RECT 63.795 206.655 65.565 207.565 ;
        RECT 66.495 206.885 68.785 207.565 ;
        RECT 66.495 206.655 67.415 206.885 ;
        RECT 68.805 206.695 69.235 207.480 ;
        RECT 69.255 206.885 71.085 207.565 ;
        RECT 69.255 206.655 70.600 206.885 ;
        RECT 71.095 206.755 76.605 207.565 ;
        RECT 76.615 206.755 82.125 207.565 ;
        RECT 82.135 206.755 84.885 207.565 ;
        RECT 85.355 206.655 88.105 207.565 ;
        RECT 88.115 206.755 93.625 207.565 ;
        RECT 94.565 206.695 94.995 207.480 ;
        RECT 95.015 206.655 96.365 207.565 ;
        RECT 96.395 206.755 101.905 207.565 ;
        RECT 101.915 206.755 107.425 207.565 ;
        RECT 107.435 206.755 110.185 207.565 ;
        RECT 110.765 206.885 114.230 207.565 ;
        RECT 113.310 206.655 114.230 206.885 ;
        RECT 114.335 206.755 119.845 207.565 ;
        RECT 120.325 206.695 120.755 207.480 ;
        RECT 120.775 206.755 126.285 207.565 ;
        RECT 126.295 206.755 131.805 207.565 ;
        RECT 131.815 206.755 137.325 207.565 ;
        RECT 137.335 206.755 142.845 207.565 ;
        RECT 142.855 206.755 145.605 207.565 ;
        RECT 145.615 206.755 146.985 207.565 ;
      LAYER nwell ;
        RECT 17.080 203.535 147.180 206.365 ;
      LAYER pwell ;
        RECT 17.275 202.335 18.645 203.145 ;
        RECT 18.655 202.335 24.165 203.145 ;
        RECT 24.175 202.335 26.005 203.145 ;
        RECT 26.015 202.335 27.845 203.245 ;
        RECT 27.855 202.335 29.685 203.145 ;
        RECT 30.165 202.420 30.595 203.205 ;
        RECT 30.615 202.335 36.125 203.145 ;
        RECT 36.135 202.335 38.885 203.145 ;
        RECT 38.895 202.335 40.725 203.015 ;
        RECT 40.735 202.335 46.245 203.145 ;
        RECT 46.255 202.335 51.765 203.145 ;
        RECT 51.775 202.335 53.605 203.145 ;
        RECT 54.665 203.015 55.595 203.245 ;
        RECT 53.760 202.335 55.595 203.015 ;
        RECT 55.925 202.420 56.355 203.205 ;
        RECT 56.375 202.335 59.125 203.245 ;
        RECT 59.150 202.335 60.965 203.245 ;
        RECT 60.975 202.335 66.485 203.145 ;
        RECT 66.495 202.335 72.005 203.145 ;
        RECT 72.015 202.335 77.525 203.145 ;
        RECT 77.535 202.335 79.365 203.145 ;
        RECT 79.835 202.335 81.665 203.245 ;
        RECT 81.685 202.420 82.115 203.205 ;
        RECT 85.650 203.015 86.560 203.235 ;
        RECT 88.095 203.015 89.445 203.245 ;
        RECT 82.135 202.335 89.445 203.015 ;
        RECT 89.590 203.015 90.510 203.245 ;
        RECT 93.175 203.045 94.120 203.245 ;
        RECT 95.455 203.045 96.385 203.245 ;
        RECT 89.590 202.335 93.055 203.015 ;
        RECT 93.175 202.565 96.385 203.045 ;
        RECT 99.910 203.015 100.820 203.235 ;
        RECT 102.355 203.015 103.705 203.245 ;
        RECT 93.175 202.365 96.245 202.565 ;
        RECT 93.175 202.335 94.120 202.365 ;
        RECT 17.415 202.125 17.585 202.335 ;
        RECT 18.795 202.125 18.965 202.335 ;
        RECT 20.175 202.125 20.345 202.315 ;
        RECT 21.555 202.125 21.725 202.315 ;
        RECT 24.315 202.145 24.485 202.335 ;
        RECT 25.235 202.125 25.405 202.315 ;
        RECT 27.530 202.145 27.700 202.335 ;
        RECT 27.995 202.145 28.165 202.335 ;
        RECT 29.830 202.175 29.950 202.285 ;
        RECT 30.755 202.145 30.925 202.335 ;
        RECT 32.595 202.125 32.765 202.315 ;
        RECT 36.275 202.145 36.445 202.335 ;
        RECT 39.035 202.145 39.205 202.335 ;
        RECT 39.960 202.125 40.130 202.315 ;
        RECT 40.875 202.145 41.045 202.335 ;
        RECT 42.715 202.125 42.885 202.315 ;
        RECT 46.395 202.145 46.565 202.335 ;
        RECT 49.155 202.125 49.325 202.315 ;
        RECT 49.615 202.125 49.785 202.315 ;
        RECT 50.995 202.125 51.165 202.315 ;
        RECT 51.915 202.145 52.085 202.335 ;
        RECT 53.760 202.315 53.925 202.335 ;
        RECT 53.755 202.125 53.925 202.315 ;
        RECT 17.275 201.315 18.645 202.125 ;
        RECT 18.655 201.345 20.025 202.125 ;
        RECT 20.035 201.315 21.405 202.125 ;
        RECT 21.415 201.445 24.165 202.125 ;
        RECT 25.095 201.445 32.405 202.125 ;
        RECT 32.455 201.445 39.765 202.125 ;
        RECT 23.235 201.215 24.165 201.445 ;
        RECT 28.610 201.225 29.520 201.445 ;
        RECT 31.055 201.215 32.405 201.445 ;
        RECT 35.970 201.225 36.880 201.445 ;
        RECT 38.415 201.215 39.765 201.445 ;
        RECT 39.815 201.215 41.165 202.125 ;
        RECT 41.195 201.445 43.025 202.125 ;
        RECT 41.195 201.215 42.540 201.445 ;
        RECT 43.045 201.255 43.475 202.040 ;
        RECT 43.645 201.215 49.465 202.125 ;
        RECT 49.475 201.315 50.845 202.125 ;
        RECT 50.855 201.215 53.260 202.125 ;
        RECT 53.615 201.445 56.825 202.125 ;
        RECT 56.980 202.095 57.150 202.315 ;
        RECT 58.815 202.145 58.985 202.335 ;
        RECT 59.275 202.145 59.445 202.335 ;
        RECT 60.655 202.125 60.825 202.315 ;
        RECT 61.115 202.145 61.285 202.335 ;
        RECT 64.335 202.125 64.505 202.315 ;
        RECT 64.795 202.125 64.965 202.315 ;
        RECT 66.635 202.145 66.805 202.335 ;
        RECT 68.470 202.175 68.590 202.285 ;
        RECT 69.390 202.175 69.510 202.285 ;
        RECT 72.155 202.145 72.325 202.335 ;
        RECT 73.075 202.125 73.245 202.315 ;
        RECT 75.375 202.145 75.545 202.315 ;
        RECT 75.830 202.175 75.950 202.285 ;
        RECT 77.675 202.145 77.845 202.335 ;
        RECT 79.510 202.175 79.630 202.285 ;
        RECT 79.980 202.145 80.150 202.335 ;
        RECT 75.375 202.125 75.525 202.145 ;
        RECT 80.895 202.125 81.065 202.315 ;
        RECT 82.275 202.125 82.445 202.335 ;
        RECT 82.735 202.125 82.905 202.315 ;
        RECT 86.425 202.170 86.585 202.280 ;
        RECT 87.335 202.125 87.505 202.315 ;
        RECT 92.855 202.145 93.025 202.335 ;
        RECT 95.430 202.125 95.600 202.315 ;
        RECT 96.075 202.145 96.245 202.365 ;
        RECT 96.395 202.335 103.705 203.015 ;
        RECT 103.850 203.015 104.770 203.245 ;
        RECT 103.850 202.335 107.315 203.015 ;
        RECT 107.445 202.420 107.875 203.205 ;
        RECT 108.395 203.015 109.745 203.245 ;
        RECT 111.280 203.015 112.190 203.235 ;
        RECT 108.395 202.335 115.705 203.015 ;
        RECT 115.715 202.335 121.225 203.145 ;
        RECT 121.235 202.335 126.745 203.145 ;
        RECT 126.755 202.335 132.265 203.145 ;
        RECT 133.205 202.420 133.635 203.205 ;
        RECT 133.655 202.335 139.165 203.145 ;
        RECT 139.175 202.335 144.685 203.145 ;
        RECT 145.615 202.335 146.985 203.145 ;
        RECT 96.535 202.145 96.705 202.335 ;
        RECT 99.290 202.145 99.460 202.315 ;
        RECT 99.325 202.125 99.460 202.145 ;
        RECT 102.980 202.125 103.150 202.315 ;
        RECT 106.195 202.125 106.365 202.315 ;
        RECT 107.115 202.145 107.285 202.335 ;
        RECT 107.575 202.125 107.745 202.315 ;
        RECT 108.030 202.175 108.150 202.285 ;
        RECT 114.660 202.125 114.830 202.315 ;
        RECT 115.395 202.125 115.565 202.335 ;
        RECT 115.855 202.145 116.025 202.335 ;
        RECT 119.075 202.125 119.245 202.315 ;
        RECT 120.915 202.125 121.085 202.315 ;
        RECT 121.375 202.145 121.545 202.335 ;
        RECT 126.435 202.125 126.605 202.315 ;
        RECT 126.895 202.145 127.065 202.335 ;
        RECT 131.955 202.125 132.125 202.315 ;
        RECT 132.425 202.180 132.585 202.290 ;
        RECT 133.795 202.145 133.965 202.335 ;
        RECT 137.475 202.125 137.645 202.315 ;
        RECT 139.315 202.145 139.485 202.335 ;
        RECT 142.995 202.125 143.165 202.315 ;
        RECT 144.845 202.180 145.005 202.290 ;
        RECT 146.675 202.125 146.845 202.335 ;
        RECT 59.555 202.095 60.505 202.125 ;
        RECT 55.690 201.215 56.825 201.445 ;
        RECT 56.835 201.415 60.505 202.095 ;
        RECT 59.555 201.215 60.505 201.415 ;
        RECT 60.515 201.215 63.265 202.125 ;
        RECT 63.285 201.215 64.635 202.125 ;
        RECT 64.655 201.315 68.325 202.125 ;
        RECT 68.805 201.255 69.235 202.040 ;
        RECT 69.810 201.445 73.275 202.125 ;
        RECT 69.810 201.215 70.730 201.445 ;
        RECT 73.595 201.305 75.525 202.125 ;
        RECT 76.390 201.445 81.205 202.125 ;
        RECT 73.595 201.215 74.545 201.305 ;
        RECT 81.225 201.215 82.575 202.125 ;
        RECT 82.705 201.445 86.170 202.125 ;
        RECT 87.195 201.445 94.505 202.125 ;
        RECT 85.250 201.215 86.170 201.445 ;
        RECT 90.710 201.225 91.620 201.445 ;
        RECT 93.155 201.215 94.505 201.445 ;
        RECT 94.565 201.255 94.995 202.040 ;
        RECT 95.015 201.445 98.915 202.125 ;
        RECT 95.015 201.215 95.945 201.445 ;
        RECT 99.325 201.215 102.825 202.125 ;
        RECT 102.835 201.215 105.755 202.125 ;
        RECT 106.065 201.215 107.415 202.125 ;
        RECT 107.435 201.315 111.105 202.125 ;
        RECT 111.345 201.445 115.245 202.125 ;
        RECT 114.315 201.215 115.245 201.445 ;
        RECT 115.255 201.315 118.925 202.125 ;
        RECT 118.935 201.315 120.305 202.125 ;
        RECT 120.325 201.255 120.755 202.040 ;
        RECT 120.775 201.315 126.285 202.125 ;
        RECT 126.295 201.315 131.805 202.125 ;
        RECT 131.815 201.315 137.325 202.125 ;
        RECT 137.335 201.315 142.845 202.125 ;
        RECT 142.855 201.315 145.605 202.125 ;
        RECT 145.615 201.315 146.985 202.125 ;
      LAYER nwell ;
        RECT 17.080 198.095 147.180 200.925 ;
      LAYER pwell ;
        RECT 17.275 196.895 18.645 197.705 ;
        RECT 18.655 196.895 21.405 197.705 ;
        RECT 24.930 197.575 25.840 197.795 ;
        RECT 27.375 197.575 28.725 197.805 ;
        RECT 21.415 196.895 28.725 197.575 ;
        RECT 28.795 196.895 30.145 197.805 ;
        RECT 30.165 196.980 30.595 197.765 ;
        RECT 30.625 196.895 33.355 197.805 ;
        RECT 34.425 197.575 35.355 197.805 ;
        RECT 33.520 196.895 35.355 197.575 ;
        RECT 35.675 197.575 36.595 197.805 ;
        RECT 35.675 196.895 37.965 197.575 ;
        RECT 38.895 196.895 41.505 197.805 ;
        RECT 42.115 197.125 45.315 197.805 ;
        RECT 46.385 197.575 47.315 197.805 ;
        RECT 42.260 196.895 45.315 197.125 ;
        RECT 45.480 196.895 47.315 197.575 ;
        RECT 48.570 196.895 50.385 197.805 ;
        RECT 51.535 197.715 52.485 197.805 ;
        RECT 50.555 196.895 52.485 197.715 ;
        RECT 52.985 196.895 55.905 197.805 ;
        RECT 55.925 196.980 56.355 197.765 ;
        RECT 56.385 196.895 57.735 197.805 ;
        RECT 59.335 197.575 62.335 197.805 ;
        RECT 57.755 197.485 62.335 197.575 ;
        RECT 62.355 197.605 63.300 197.805 ;
        RECT 64.635 197.605 65.565 197.805 ;
        RECT 57.755 197.125 62.345 197.485 ;
        RECT 57.755 196.895 59.325 197.125 ;
        RECT 61.415 196.935 62.345 197.125 ;
        RECT 62.355 197.125 65.565 197.605 ;
        RECT 61.415 196.895 62.335 196.935 ;
        RECT 62.355 196.925 65.425 197.125 ;
        RECT 62.355 196.895 63.300 196.925 ;
        RECT 17.415 196.685 17.585 196.895 ;
        RECT 18.795 196.845 18.965 196.895 ;
        RECT 18.790 196.735 18.965 196.845 ;
        RECT 18.795 196.705 18.965 196.735 ;
        RECT 21.555 196.705 21.725 196.895 ;
        RECT 26.155 196.685 26.325 196.875 ;
        RECT 28.910 196.705 29.080 196.895 ;
        RECT 29.375 196.685 29.545 196.875 ;
        RECT 29.840 196.685 30.010 196.875 ;
        RECT 30.755 196.705 30.925 196.895 ;
        RECT 33.520 196.875 33.685 196.895 ;
        RECT 33.050 196.735 33.170 196.845 ;
        RECT 33.510 196.705 33.685 196.875 ;
        RECT 37.655 196.705 37.825 196.895 ;
        RECT 39.040 196.875 39.210 196.895 ;
        RECT 38.125 196.740 38.285 196.850 ;
        RECT 17.275 195.875 18.645 196.685 ;
        RECT 19.155 196.005 26.465 196.685 ;
        RECT 26.475 196.005 29.685 196.685 ;
        RECT 19.155 195.775 20.505 196.005 ;
        RECT 22.040 195.785 22.950 196.005 ;
        RECT 26.475 195.775 27.610 196.005 ;
        RECT 29.695 195.775 32.615 196.685 ;
        RECT 33.510 196.655 33.680 196.705 ;
        RECT 38.575 196.685 38.745 196.875 ;
        RECT 39.035 196.705 39.210 196.875 ;
        RECT 41.790 196.735 41.910 196.845 ;
        RECT 42.260 196.705 42.430 196.895 ;
        RECT 45.480 196.875 45.645 196.895 ;
        RECT 39.035 196.685 39.205 196.705 ;
        RECT 43.640 196.685 43.810 196.875 ;
        RECT 45.475 196.705 45.645 196.875 ;
        RECT 47.315 196.685 47.485 196.875 ;
        RECT 47.775 196.685 47.945 196.875 ;
        RECT 48.695 196.705 48.865 196.895 ;
        RECT 50.555 196.875 50.705 196.895 ;
        RECT 50.535 196.845 50.705 196.875 ;
        RECT 50.530 196.735 50.705 196.845 ;
        RECT 50.535 196.705 50.705 196.735 ;
        RECT 50.990 196.685 51.160 196.875 ;
        RECT 34.710 196.655 35.665 196.685 ;
        RECT 33.385 195.975 35.665 196.655 ;
        RECT 34.710 195.775 35.665 195.975 ;
        RECT 35.675 195.775 38.885 196.685 ;
        RECT 38.895 195.775 42.105 196.685 ;
        RECT 43.045 195.815 43.475 196.600 ;
        RECT 43.640 196.455 45.330 196.685 ;
        RECT 43.495 195.775 45.330 196.455 ;
        RECT 45.795 196.005 47.625 196.685 ;
        RECT 47.635 195.875 50.385 196.685 ;
        RECT 50.875 195.775 52.225 196.685 ;
        RECT 52.370 196.655 52.540 196.875 ;
        RECT 54.675 196.685 54.845 196.875 ;
        RECT 55.590 196.705 55.760 196.895 ;
        RECT 57.435 196.705 57.605 196.895 ;
        RECT 57.895 196.705 58.065 196.895 ;
        RECT 61.110 196.685 61.280 196.875 ;
        RECT 63.875 196.685 64.045 196.875 ;
        RECT 64.335 196.685 64.505 196.875 ;
        RECT 65.255 196.705 65.425 196.925 ;
        RECT 65.575 196.895 67.405 197.805 ;
        RECT 67.415 196.895 68.785 197.705 ;
        RECT 68.795 196.895 70.145 197.805 ;
        RECT 73.690 197.575 74.600 197.795 ;
        RECT 76.135 197.575 77.485 197.805 ;
        RECT 70.175 196.895 77.485 197.575 ;
        RECT 78.000 196.895 79.365 197.575 ;
        RECT 79.375 196.895 81.205 197.705 ;
        RECT 81.685 196.980 82.115 197.765 ;
        RECT 82.135 196.895 83.965 197.705 ;
        RECT 83.985 196.895 86.715 197.805 ;
        RECT 86.735 196.895 88.565 197.705 ;
        RECT 89.035 196.895 90.385 197.805 ;
        RECT 90.435 196.895 91.785 197.805 ;
        RECT 91.805 196.895 93.155 197.805 ;
        RECT 93.185 196.895 95.915 197.805 ;
        RECT 95.935 196.895 99.605 197.805 ;
        RECT 99.925 197.575 100.855 197.805 ;
        RECT 99.925 196.895 101.760 197.575 ;
        RECT 101.930 196.895 105.585 197.805 ;
        RECT 105.605 196.895 106.955 197.805 ;
        RECT 107.445 196.980 107.875 197.765 ;
        RECT 107.895 196.895 109.245 197.805 ;
        RECT 110.195 197.575 111.125 197.805 ;
        RECT 114.430 197.575 115.350 197.805 ;
        RECT 110.195 196.895 114.095 197.575 ;
        RECT 114.430 196.895 117.895 197.575 ;
        RECT 118.015 196.895 121.685 197.705 ;
        RECT 122.155 196.895 125.365 197.805 ;
        RECT 125.375 196.895 130.885 197.705 ;
        RECT 130.895 196.895 132.725 197.705 ;
        RECT 133.205 196.980 133.635 197.765 ;
        RECT 133.655 196.895 139.165 197.705 ;
        RECT 139.175 196.895 144.685 197.705 ;
        RECT 145.615 196.895 146.985 197.705 ;
        RECT 65.720 196.705 65.890 196.895 ;
        RECT 67.555 196.705 67.725 196.895 ;
        RECT 68.025 196.730 68.185 196.840 ;
        RECT 68.940 196.705 69.110 196.895 ;
        RECT 69.395 196.685 69.565 196.875 ;
        RECT 70.315 196.705 70.485 196.895 ;
        RECT 71.240 196.685 71.410 196.875 ;
        RECT 77.675 196.705 77.845 196.875 ;
        RECT 79.515 196.705 79.685 196.895 ;
        RECT 79.975 196.685 80.145 196.875 ;
        RECT 80.430 196.735 80.550 196.845 ;
        RECT 80.895 196.685 81.065 196.875 ;
        RECT 81.350 196.735 81.470 196.845 ;
        RECT 82.275 196.705 82.445 196.895 ;
        RECT 84.115 196.705 84.285 196.895 ;
        RECT 86.875 196.705 87.045 196.895 ;
        RECT 88.255 196.685 88.425 196.875 ;
        RECT 88.710 196.735 88.830 196.845 ;
        RECT 90.100 196.705 90.270 196.895 ;
        RECT 91.470 196.705 91.640 196.895 ;
        RECT 92.855 196.705 93.025 196.895 ;
        RECT 93.785 196.730 93.945 196.840 ;
        RECT 95.155 196.685 95.325 196.875 ;
        RECT 95.615 196.705 95.785 196.895 ;
        RECT 96.075 196.705 96.245 196.895 ;
        RECT 101.595 196.875 101.760 196.895 ;
        RECT 97.915 196.685 98.085 196.875 ;
        RECT 101.130 196.735 101.250 196.845 ;
        RECT 101.595 196.705 101.765 196.875 ;
        RECT 104.350 196.685 104.520 196.875 ;
        RECT 104.815 196.685 104.985 196.875 ;
        RECT 105.270 196.705 105.440 196.895 ;
        RECT 105.735 196.705 105.905 196.895 ;
        RECT 106.195 196.685 106.365 196.875 ;
        RECT 107.110 196.735 107.230 196.845 ;
        RECT 107.575 196.685 107.745 196.875 ;
        RECT 108.040 196.705 108.210 196.895 ;
        RECT 109.425 196.740 109.585 196.850 ;
        RECT 110.610 196.705 110.780 196.895 ;
        RECT 114.935 196.685 115.105 196.875 ;
        RECT 117.695 196.705 117.865 196.895 ;
        RECT 118.155 196.705 118.325 196.895 ;
        RECT 121.190 196.685 121.360 196.875 ;
        RECT 121.830 196.735 121.950 196.845 ;
        RECT 125.055 196.705 125.225 196.895 ;
        RECT 125.515 196.705 125.685 196.895 ;
        RECT 131.035 196.705 131.205 196.895 ;
        RECT 132.875 196.845 133.045 196.875 ;
        RECT 132.870 196.735 133.045 196.845 ;
        RECT 132.875 196.685 133.045 196.735 ;
        RECT 133.795 196.705 133.965 196.895 ;
        RECT 134.715 196.685 134.885 196.875 ;
        RECT 135.175 196.685 135.345 196.875 ;
        RECT 139.315 196.705 139.485 196.895 ;
        RECT 140.695 196.685 140.865 196.875 ;
        RECT 144.375 196.685 144.545 196.875 ;
        RECT 144.845 196.740 145.005 196.850 ;
        RECT 146.675 196.685 146.845 196.895 ;
        RECT 53.570 196.655 54.525 196.685 ;
        RECT 52.245 195.975 54.525 196.655 ;
        RECT 53.570 195.775 54.525 195.975 ;
        RECT 54.535 195.775 57.745 196.685 ;
        RECT 57.950 195.775 61.425 196.685 ;
        RECT 61.445 195.775 64.175 196.685 ;
        RECT 64.195 195.875 67.865 196.685 ;
        RECT 68.805 195.815 69.235 196.600 ;
        RECT 69.255 195.875 71.085 196.685 ;
        RECT 71.095 195.775 72.865 196.685 ;
        RECT 72.975 196.005 80.285 196.685 ;
        RECT 80.755 196.005 88.065 196.685 ;
        RECT 72.975 195.775 74.325 196.005 ;
        RECT 75.860 195.785 76.770 196.005 ;
        RECT 84.270 195.785 85.180 196.005 ;
        RECT 86.715 195.775 88.065 196.005 ;
        RECT 88.115 195.875 93.625 196.685 ;
        RECT 94.565 195.815 94.995 196.600 ;
        RECT 95.015 195.875 97.765 196.685 ;
        RECT 97.775 195.775 100.985 196.685 ;
        RECT 101.745 195.775 104.665 196.685 ;
        RECT 104.685 195.775 106.035 196.685 ;
        RECT 106.055 195.875 107.425 196.685 ;
        RECT 107.435 196.005 114.745 196.685 ;
        RECT 110.950 195.785 111.860 196.005 ;
        RECT 113.395 195.775 114.745 196.005 ;
        RECT 114.795 195.875 120.305 196.685 ;
        RECT 120.325 195.815 120.755 196.600 ;
        RECT 120.775 196.005 124.675 196.685 ;
        RECT 125.875 196.005 133.185 196.685 ;
        RECT 133.195 196.005 135.025 196.685 ;
        RECT 120.775 195.775 121.705 196.005 ;
        RECT 125.875 195.775 127.225 196.005 ;
        RECT 128.760 195.785 129.670 196.005 ;
        RECT 135.035 195.875 140.545 196.685 ;
        RECT 140.555 195.875 144.225 196.685 ;
        RECT 144.235 195.875 145.605 196.685 ;
        RECT 145.615 195.875 146.985 196.685 ;
      LAYER nwell ;
        RECT 17.080 192.655 147.180 195.485 ;
      LAYER pwell ;
        RECT 17.275 191.455 18.645 192.265 ;
        RECT 18.655 191.455 22.325 192.265 ;
        RECT 22.795 192.135 23.715 192.365 ;
        RECT 26.015 192.135 26.935 192.365 ;
        RECT 22.795 191.455 25.085 192.135 ;
        RECT 26.015 191.455 28.305 192.135 ;
        RECT 28.325 191.455 29.675 192.365 ;
        RECT 30.165 191.540 30.595 192.325 ;
        RECT 30.615 191.455 36.125 192.265 ;
        RECT 36.135 191.455 37.505 192.265 ;
        RECT 37.515 191.455 40.265 192.365 ;
        RECT 40.295 191.455 41.645 192.365 ;
        RECT 41.855 192.275 42.805 192.365 ;
        RECT 41.855 191.455 43.785 192.275 ;
        RECT 44.010 191.455 54.030 192.365 ;
        RECT 54.075 191.455 55.905 192.265 ;
        RECT 55.925 191.540 56.355 192.325 ;
        RECT 56.375 191.455 59.585 192.365 ;
        RECT 59.795 192.275 60.745 192.365 ;
        RECT 59.795 191.455 61.725 192.275 ;
        RECT 61.895 191.455 67.405 192.265 ;
        RECT 67.415 191.455 71.085 192.265 ;
        RECT 71.095 191.455 72.465 192.265 ;
        RECT 72.575 191.455 75.685 192.365 ;
        RECT 76.850 191.455 81.665 192.135 ;
        RECT 81.685 191.540 82.115 192.325 ;
        RECT 82.135 191.455 87.645 192.265 ;
        RECT 87.655 191.455 91.325 192.265 ;
        RECT 91.430 192.135 92.350 192.365 ;
        RECT 98.530 192.135 99.440 192.355 ;
        RECT 100.975 192.135 102.325 192.365 ;
        RECT 91.430 191.455 94.895 192.135 ;
        RECT 95.015 191.455 102.325 192.135 ;
        RECT 102.375 192.135 103.305 192.365 ;
        RECT 102.375 191.455 106.275 192.135 ;
        RECT 107.445 191.540 107.875 192.325 ;
        RECT 111.410 192.135 112.320 192.355 ;
        RECT 113.855 192.135 115.205 192.365 ;
        RECT 107.895 191.455 115.205 192.135 ;
        RECT 115.255 191.455 118.005 192.265 ;
        RECT 118.015 192.135 118.945 192.365 ;
        RECT 124.810 192.135 125.730 192.365 ;
        RECT 118.015 191.455 121.915 192.135 ;
        RECT 122.265 191.455 125.730 192.135 ;
        RECT 125.835 191.455 127.205 192.265 ;
        RECT 129.870 192.135 130.790 192.365 ;
        RECT 131.380 192.135 132.725 192.365 ;
        RECT 127.325 191.455 130.790 192.135 ;
        RECT 130.895 191.455 132.725 192.135 ;
        RECT 133.205 191.540 133.635 192.325 ;
        RECT 133.655 191.455 136.865 192.365 ;
        RECT 136.875 191.455 142.385 192.265 ;
        RECT 142.395 191.455 145.145 192.265 ;
        RECT 145.615 191.455 146.985 192.265 ;
        RECT 17.415 191.245 17.585 191.455 ;
        RECT 18.795 191.245 18.965 191.455 ;
        RECT 24.775 191.435 24.945 191.455 ;
        RECT 22.470 191.295 22.590 191.405 ;
        RECT 24.310 191.295 24.430 191.405 ;
        RECT 24.770 191.265 24.945 191.435 ;
        RECT 25.245 191.300 25.405 191.410 ;
        RECT 24.770 191.245 24.940 191.265 ;
        RECT 26.155 191.245 26.325 191.435 ;
        RECT 27.995 191.265 28.165 191.455 ;
        RECT 28.455 191.265 28.625 191.455 ;
        RECT 29.830 191.295 29.950 191.405 ;
        RECT 30.755 191.265 30.925 191.455 ;
        RECT 31.675 191.245 31.845 191.435 ;
        RECT 36.275 191.265 36.445 191.455 ;
        RECT 37.660 191.265 37.830 191.455 ;
        RECT 38.570 191.245 38.740 191.435 ;
        RECT 40.410 191.265 40.580 191.455 ;
        RECT 43.635 191.435 43.785 191.455 ;
        RECT 42.250 191.245 42.420 191.435 ;
        RECT 42.710 191.295 42.830 191.405 ;
        RECT 43.635 191.245 43.805 191.435 ;
        RECT 44.095 191.265 44.265 191.455 ;
        RECT 48.695 191.245 48.865 191.435 ;
        RECT 54.215 191.245 54.385 191.455 ;
        RECT 54.675 191.245 54.845 191.435 ;
        RECT 56.515 191.245 56.685 191.455 ;
        RECT 61.575 191.435 61.725 191.455 ;
        RECT 59.730 191.245 59.900 191.435 ;
        RECT 60.190 191.295 60.310 191.405 ;
        RECT 17.275 190.435 18.645 191.245 ;
        RECT 18.655 190.435 24.165 191.245 ;
        RECT 24.655 190.335 26.005 191.245 ;
        RECT 26.015 190.435 31.525 191.245 ;
        RECT 31.535 190.435 35.205 191.245 ;
        RECT 35.410 190.335 38.885 191.245 ;
        RECT 39.090 190.335 42.565 191.245 ;
        RECT 43.045 190.375 43.475 191.160 ;
        RECT 43.495 190.565 48.310 191.245 ;
        RECT 48.605 190.335 51.765 191.245 ;
        RECT 52.435 190.435 54.525 191.245 ;
        RECT 54.535 190.435 56.365 191.245 ;
        RECT 56.385 190.335 57.735 191.245 ;
        RECT 57.770 190.565 60.045 191.245 ;
        RECT 60.660 191.215 60.830 191.435 ;
        RECT 61.575 191.265 61.745 191.435 ;
        RECT 62.035 191.265 62.205 191.455 ;
        RECT 63.415 191.245 63.585 191.435 ;
        RECT 66.635 191.265 66.805 191.435 ;
        RECT 67.555 191.265 67.725 191.455 ;
        RECT 66.640 191.245 66.805 191.265 ;
        RECT 70.775 191.245 70.945 191.435 ;
        RECT 71.235 191.245 71.405 191.455 ;
        RECT 72.615 191.265 72.785 191.455 ;
        RECT 75.845 191.300 76.005 191.410 ;
        RECT 76.755 191.245 76.925 191.435 ;
        RECT 77.210 191.295 77.330 191.405 ;
        RECT 77.675 191.265 77.845 191.435 ;
        RECT 80.900 191.245 81.070 191.435 ;
        RECT 81.355 191.265 81.525 191.455 ;
        RECT 82.275 191.245 82.445 191.455 ;
        RECT 87.795 191.265 87.965 191.455 ;
        RECT 88.990 191.245 89.160 191.435 ;
        RECT 92.855 191.245 93.025 191.435 ;
        RECT 94.695 191.265 94.865 191.455 ;
        RECT 95.155 191.405 95.325 191.455 ;
        RECT 95.150 191.295 95.325 191.405 ;
        RECT 95.155 191.265 95.325 191.295 ;
        RECT 95.890 191.245 96.060 191.435 ;
        RECT 99.755 191.245 99.925 191.435 ;
        RECT 102.790 191.265 102.960 191.455 ;
        RECT 103.435 191.245 103.605 191.435 ;
        RECT 106.665 191.300 106.825 191.410 ;
        RECT 107.115 191.245 107.285 191.435 ;
        RECT 108.035 191.265 108.205 191.455 ;
        RECT 108.770 191.245 108.940 191.435 ;
        RECT 115.395 191.265 115.565 191.455 ;
        RECT 115.855 191.245 116.025 191.435 ;
        RECT 116.590 191.245 116.760 191.435 ;
        RECT 118.430 191.265 118.600 191.455 ;
        RECT 120.915 191.245 121.085 191.435 ;
        RECT 122.295 191.265 122.465 191.455 ;
        RECT 125.975 191.265 126.145 191.455 ;
        RECT 127.355 191.265 127.525 191.455 ;
        RECT 131.035 191.265 131.205 191.455 ;
        RECT 131.495 191.245 131.665 191.435 ;
        RECT 131.955 191.265 132.125 191.435 ;
        RECT 132.870 191.295 132.990 191.405 ;
        RECT 136.555 191.265 136.725 191.455 ;
        RECT 137.015 191.265 137.185 191.455 ;
        RECT 131.960 191.245 132.125 191.265 ;
        RECT 141.155 191.245 141.325 191.435 ;
        RECT 141.615 191.245 141.785 191.435 ;
        RECT 142.535 191.265 142.705 191.455 ;
        RECT 145.290 191.295 145.410 191.405 ;
        RECT 146.675 191.245 146.845 191.455 ;
        RECT 62.320 191.215 63.265 191.245 ;
        RECT 57.770 190.335 59.140 190.565 ;
        RECT 60.515 190.535 63.265 191.215 ;
        RECT 62.320 190.335 63.265 190.535 ;
        RECT 63.275 190.335 66.485 191.245 ;
        RECT 66.640 190.565 68.475 191.245 ;
        RECT 67.545 190.335 68.475 190.565 ;
        RECT 68.805 190.375 69.235 191.160 ;
        RECT 69.255 190.335 71.070 191.245 ;
        RECT 71.095 190.565 73.385 191.245 ;
        RECT 72.465 190.335 73.385 190.565 ;
        RECT 73.490 190.565 76.955 191.245 ;
        RECT 77.940 190.565 80.365 191.245 ;
        RECT 73.490 190.335 74.410 190.565 ;
        RECT 80.755 190.335 82.105 191.245 ;
        RECT 82.135 190.435 87.645 191.245 ;
        RECT 88.575 190.565 92.475 191.245 ;
        RECT 88.575 190.335 89.505 190.565 ;
        RECT 92.715 190.435 94.545 191.245 ;
        RECT 94.565 190.375 94.995 191.160 ;
        RECT 95.475 190.565 99.375 191.245 ;
        RECT 99.725 190.565 103.190 191.245 ;
        RECT 103.405 190.565 106.870 191.245 ;
        RECT 95.475 190.335 96.405 190.565 ;
        RECT 102.270 190.335 103.190 190.565 ;
        RECT 105.950 190.335 106.870 190.565 ;
        RECT 106.975 190.435 108.345 191.245 ;
        RECT 108.355 190.565 112.255 191.245 ;
        RECT 112.590 190.565 116.055 191.245 ;
        RECT 116.175 190.565 120.075 191.245 ;
        RECT 108.355 190.335 109.285 190.565 ;
        RECT 112.590 190.335 113.510 190.565 ;
        RECT 116.175 190.335 117.105 190.565 ;
        RECT 120.325 190.375 120.755 191.160 ;
        RECT 120.775 190.565 128.085 191.245 ;
        RECT 124.290 190.345 125.200 190.565 ;
        RECT 126.735 190.335 128.085 190.565 ;
        RECT 128.230 190.565 131.695 191.245 ;
        RECT 131.960 190.565 133.795 191.245 ;
        RECT 128.230 190.335 129.150 190.565 ;
        RECT 132.865 190.335 133.795 190.565 ;
        RECT 134.155 190.565 141.465 191.245 ;
        RECT 134.155 190.335 135.505 190.565 ;
        RECT 137.040 190.345 137.950 190.565 ;
        RECT 141.475 190.435 145.145 191.245 ;
        RECT 145.615 190.435 146.985 191.245 ;
      LAYER nwell ;
        RECT 17.080 187.215 147.180 190.045 ;
      LAYER pwell ;
        RECT 17.275 186.015 18.645 186.825 ;
        RECT 18.655 186.015 22.325 186.825 ;
        RECT 22.335 186.695 23.255 186.925 ;
        RECT 25.685 186.695 26.615 186.925 ;
        RECT 22.335 186.015 24.625 186.695 ;
        RECT 24.780 186.015 26.615 186.695 ;
        RECT 26.945 186.015 28.295 186.925 ;
        RECT 28.315 186.015 29.665 186.925 ;
        RECT 30.165 186.100 30.595 186.885 ;
        RECT 30.615 186.015 34.285 186.825 ;
        RECT 34.950 186.015 38.425 186.925 ;
        RECT 38.455 186.015 39.805 186.925 ;
        RECT 39.815 186.725 40.745 186.925 ;
        RECT 42.080 186.725 43.025 186.925 ;
        RECT 39.815 186.245 43.025 186.725 ;
        RECT 39.955 186.045 43.025 186.245 ;
        RECT 17.415 185.805 17.585 186.015 ;
        RECT 18.795 185.825 18.965 186.015 ;
        RECT 19.715 185.805 19.885 185.995 ;
        RECT 24.315 185.825 24.485 186.015 ;
        RECT 24.780 185.995 24.945 186.015 ;
        RECT 24.775 185.825 24.945 185.995 ;
        RECT 27.075 185.805 27.245 186.015 ;
        RECT 29.380 185.825 29.550 186.015 ;
        RECT 29.830 185.855 29.950 185.965 ;
        RECT 30.755 185.825 30.925 186.015 ;
        RECT 31.215 185.805 31.385 185.995 ;
        RECT 31.675 185.805 31.845 185.995 ;
        RECT 33.055 185.805 33.225 185.995 ;
        RECT 34.430 185.855 34.550 185.965 ;
        RECT 36.730 185.855 36.850 185.965 ;
        RECT 37.195 185.825 37.365 185.995 ;
        RECT 38.110 185.825 38.280 186.015 ;
        RECT 38.570 185.825 38.740 186.015 ;
        RECT 39.955 185.825 40.125 186.045 ;
        RECT 42.080 186.015 43.025 186.045 ;
        RECT 43.270 186.015 48.085 186.695 ;
        RECT 48.095 186.015 53.605 186.825 ;
        RECT 53.615 186.015 55.445 186.825 ;
        RECT 55.925 186.100 56.355 186.885 ;
        RECT 56.835 186.015 58.665 186.925 ;
        RECT 58.675 186.015 61.080 186.925 ;
        RECT 61.435 186.015 65.095 186.925 ;
        RECT 65.115 186.015 70.625 186.825 ;
        RECT 70.635 186.015 72.005 186.825 ;
        RECT 72.015 186.015 73.785 186.925 ;
        RECT 73.895 186.695 75.245 186.925 ;
        RECT 76.780 186.695 77.690 186.915 ;
        RECT 73.895 186.015 81.205 186.695 ;
        RECT 81.685 186.100 82.115 186.885 ;
        RECT 82.135 186.015 83.965 186.825 ;
        RECT 87.950 186.695 88.860 186.915 ;
        RECT 90.395 186.695 91.745 186.925 ;
        RECT 84.435 186.015 91.745 186.695 ;
        RECT 92.755 186.695 94.105 186.925 ;
        RECT 95.640 186.695 96.550 186.915 ;
        RECT 100.075 186.695 101.005 186.925 ;
        RECT 92.755 186.015 100.065 186.695 ;
        RECT 100.075 186.015 103.975 186.695 ;
        RECT 104.215 186.015 106.965 186.825 ;
        RECT 107.445 186.100 107.875 186.885 ;
        RECT 107.895 186.015 111.105 186.925 ;
        RECT 111.115 186.015 116.625 186.825 ;
        RECT 116.675 186.695 118.025 186.925 ;
        RECT 119.560 186.695 120.470 186.915 ;
        RECT 116.675 186.015 123.985 186.695 ;
        RECT 123.995 186.015 127.205 186.925 ;
        RECT 127.215 186.725 128.170 186.925 ;
        RECT 127.215 186.045 129.495 186.725 ;
        RECT 127.215 186.015 128.170 186.045 ;
        RECT 37.205 185.805 37.365 185.825 ;
        RECT 41.340 185.805 41.510 185.995 ;
        RECT 42.710 185.855 42.830 185.965 ;
        RECT 43.635 185.805 43.805 185.995 ;
        RECT 46.855 185.805 47.025 185.995 ;
        RECT 47.775 185.825 47.945 186.015 ;
        RECT 48.235 185.825 48.405 186.015 ;
        RECT 52.375 185.805 52.545 185.995 ;
        RECT 53.755 185.825 53.925 186.015 ;
        RECT 55.590 185.855 55.710 185.965 ;
        RECT 56.510 185.855 56.630 185.965 ;
        RECT 56.980 185.825 57.150 186.015 ;
        RECT 57.895 185.805 58.065 185.995 ;
        RECT 58.815 185.825 58.985 186.015 ;
        RECT 60.650 185.855 60.770 185.965 ;
        RECT 61.120 185.805 61.290 185.995 ;
        RECT 62.490 185.855 62.610 185.965 ;
        RECT 62.945 185.805 63.115 185.995 ;
        RECT 64.800 185.825 64.970 186.015 ;
        RECT 65.255 185.825 65.425 186.015 ;
        RECT 66.175 185.805 66.345 185.995 ;
        RECT 69.395 185.805 69.565 185.995 ;
        RECT 70.775 185.825 70.945 186.015 ;
        RECT 72.160 185.825 72.330 186.015 ;
        RECT 73.075 185.805 73.245 185.995 ;
        RECT 74.455 185.805 74.625 185.995 ;
        RECT 78.140 185.805 78.310 185.995 ;
        RECT 79.515 185.805 79.685 185.995 ;
        RECT 80.895 185.825 81.065 186.015 ;
        RECT 81.350 185.855 81.470 185.965 ;
        RECT 82.275 185.825 82.445 186.015 ;
        RECT 84.110 185.855 84.230 185.965 ;
        RECT 84.575 185.825 84.745 186.015 ;
        RECT 85.035 185.805 85.205 185.995 ;
        RECT 86.870 185.855 86.990 185.965 ;
        RECT 87.335 185.805 87.505 185.995 ;
        RECT 91.945 185.860 92.105 185.970 ;
        RECT 98.375 185.805 98.545 185.995 ;
        RECT 99.755 185.825 99.925 186.015 ;
        RECT 100.490 185.825 100.660 186.015 ;
        RECT 102.055 185.805 102.225 185.995 ;
        RECT 104.355 185.825 104.525 186.015 ;
        RECT 105.735 185.805 105.905 185.995 ;
        RECT 106.195 185.825 106.365 185.995 ;
        RECT 107.110 185.855 107.230 185.965 ;
        RECT 110.795 185.825 110.965 186.015 ;
        RECT 111.255 185.825 111.425 186.015 ;
        RECT 112.175 185.805 112.345 185.995 ;
        RECT 112.635 185.805 112.805 185.995 ;
        RECT 118.155 185.805 118.325 185.995 ;
        RECT 119.990 185.855 120.110 185.965 ;
        RECT 120.915 185.805 121.085 185.995 ;
        RECT 123.675 185.965 123.845 186.015 ;
        RECT 123.670 185.855 123.845 185.965 ;
        RECT 123.675 185.825 123.845 185.855 ;
        RECT 125.975 185.825 126.145 185.995 ;
        RECT 125.975 185.805 126.140 185.825 ;
        RECT 126.435 185.805 126.605 185.995 ;
        RECT 126.895 185.825 127.065 186.015 ;
        RECT 129.200 185.825 129.370 186.045 ;
        RECT 129.515 186.015 133.185 186.925 ;
        RECT 133.205 186.100 133.635 186.885 ;
        RECT 137.170 186.695 138.080 186.915 ;
        RECT 139.615 186.695 140.965 186.925 ;
        RECT 133.655 186.015 140.965 186.695 ;
        RECT 141.015 186.015 144.225 186.925 ;
        RECT 144.235 186.015 145.605 186.825 ;
        RECT 145.615 186.015 146.985 186.825 ;
        RECT 129.650 185.805 129.820 185.995 ;
        RECT 130.125 185.850 130.285 185.960 ;
        RECT 131.030 185.805 131.200 185.995 ;
        RECT 132.870 185.825 133.040 186.015 ;
        RECT 133.795 185.825 133.965 186.015 ;
        RECT 135.170 185.805 135.340 185.995 ;
        RECT 137.015 185.805 137.185 185.995 ;
        RECT 137.475 185.805 137.645 185.995 ;
        RECT 143.915 185.825 144.085 186.015 ;
        RECT 144.375 185.825 144.545 186.015 ;
        RECT 144.845 185.850 145.005 185.960 ;
        RECT 146.675 185.805 146.845 186.015 ;
        RECT 17.275 184.995 18.645 185.805 ;
        RECT 19.575 185.125 26.885 185.805 ;
        RECT 26.935 185.125 29.225 185.805 ;
        RECT 23.090 184.905 24.000 185.125 ;
        RECT 25.535 184.895 26.885 185.125 ;
        RECT 28.305 184.895 29.225 185.125 ;
        RECT 29.235 185.125 31.525 185.805 ;
        RECT 29.235 184.895 30.155 185.125 ;
        RECT 31.545 184.895 32.895 185.805 ;
        RECT 32.915 184.995 36.585 185.805 ;
        RECT 37.205 184.895 40.860 185.805 ;
        RECT 41.195 184.895 42.545 185.805 ;
        RECT 43.045 184.935 43.475 185.720 ;
        RECT 43.575 184.895 46.575 185.805 ;
        RECT 46.715 184.995 52.225 185.805 ;
        RECT 52.235 184.995 57.745 185.805 ;
        RECT 57.755 184.995 60.505 185.805 ;
        RECT 60.975 184.895 62.325 185.805 ;
        RECT 62.815 184.895 66.025 185.805 ;
        RECT 66.035 184.995 68.785 185.805 ;
        RECT 68.805 184.935 69.235 185.720 ;
        RECT 69.255 184.995 72.925 185.805 ;
        RECT 72.935 184.995 74.305 185.805 ;
        RECT 74.425 185.125 77.890 185.805 ;
        RECT 76.970 184.895 77.890 185.125 ;
        RECT 77.995 184.895 79.345 185.805 ;
        RECT 79.375 184.995 84.885 185.805 ;
        RECT 84.895 184.995 86.725 185.805 ;
        RECT 87.195 185.125 94.505 185.805 ;
        RECT 90.710 184.905 91.620 185.125 ;
        RECT 93.155 184.895 94.505 185.125 ;
        RECT 94.565 184.935 94.995 185.720 ;
        RECT 95.110 185.125 98.575 185.805 ;
        RECT 98.790 185.125 102.255 185.805 ;
        RECT 102.470 185.125 105.935 185.805 ;
        RECT 106.460 185.125 108.885 185.805 ;
        RECT 109.275 185.125 112.485 185.805 ;
        RECT 95.110 184.895 96.030 185.125 ;
        RECT 98.790 184.895 99.710 185.125 ;
        RECT 102.470 184.895 103.390 185.125 ;
        RECT 109.275 184.895 110.410 185.125 ;
        RECT 112.495 184.995 118.005 185.805 ;
        RECT 118.015 184.995 119.845 185.805 ;
        RECT 120.325 184.935 120.755 185.720 ;
        RECT 120.775 184.995 123.525 185.805 ;
        RECT 124.305 185.125 126.140 185.805 ;
        RECT 126.295 185.125 128.585 185.805 ;
        RECT 124.305 184.895 125.235 185.125 ;
        RECT 127.665 184.895 128.585 185.125 ;
        RECT 128.615 184.895 129.965 185.805 ;
        RECT 130.915 184.895 132.265 185.805 ;
        RECT 132.565 184.895 135.485 185.805 ;
        RECT 135.495 185.125 137.325 185.805 ;
        RECT 137.335 185.125 144.645 185.805 ;
        RECT 140.850 184.905 141.760 185.125 ;
        RECT 143.295 184.895 144.645 185.125 ;
        RECT 145.615 184.995 146.985 185.805 ;
      LAYER nwell ;
        RECT 17.080 181.775 147.180 184.605 ;
      LAYER pwell ;
        RECT 17.275 180.575 18.645 181.385 ;
        RECT 18.655 180.575 21.405 181.385 ;
        RECT 21.915 181.255 23.265 181.485 ;
        RECT 24.800 181.255 25.710 181.475 ;
        RECT 21.915 180.575 29.225 181.255 ;
        RECT 30.165 180.660 30.595 181.445 ;
        RECT 30.615 180.575 36.125 181.385 ;
        RECT 36.135 180.575 37.505 181.385 ;
        RECT 37.645 180.575 40.645 181.485 ;
        RECT 40.735 181.255 41.655 181.485 ;
        RECT 40.735 180.575 44.320 181.255 ;
        RECT 44.435 180.575 45.785 181.485 ;
        RECT 46.295 181.255 47.645 181.485 ;
        RECT 49.180 181.255 50.090 181.475 ;
        RECT 46.295 180.575 53.605 181.255 ;
        RECT 53.615 180.575 55.445 181.385 ;
        RECT 55.925 180.660 56.355 181.445 ;
        RECT 56.375 180.575 61.885 181.385 ;
        RECT 61.895 180.575 63.725 181.385 ;
        RECT 64.195 181.255 65.115 181.485 ;
        RECT 64.195 180.575 66.485 181.255 ;
        RECT 66.495 180.575 68.310 181.485 ;
        RECT 68.335 180.575 69.685 181.485 ;
        RECT 71.775 181.395 72.725 181.485 ;
        RECT 70.795 180.575 72.725 181.395 ;
        RECT 72.975 181.255 74.325 181.485 ;
        RECT 75.860 181.255 76.770 181.475 ;
        RECT 72.975 180.575 80.285 181.255 ;
        RECT 80.295 180.575 81.665 181.385 ;
        RECT 81.685 180.660 82.115 181.445 ;
        RECT 82.135 180.575 85.805 181.385 ;
        RECT 89.790 181.255 90.700 181.475 ;
        RECT 92.235 181.255 93.585 181.485 ;
        RECT 86.275 180.575 93.585 181.255 ;
        RECT 93.635 181.255 94.565 181.485 ;
        RECT 93.635 180.575 97.535 181.255 ;
        RECT 97.775 180.575 100.525 181.385 ;
        RECT 100.535 181.255 101.465 181.485 ;
        RECT 100.535 180.575 104.435 181.255 ;
        RECT 105.615 180.575 106.965 181.485 ;
        RECT 107.445 180.660 107.875 181.445 ;
        RECT 111.410 181.255 112.320 181.475 ;
        RECT 113.855 181.255 115.205 181.485 ;
        RECT 107.895 180.575 115.205 181.255 ;
        RECT 115.255 180.575 120.765 181.385 ;
        RECT 120.775 180.575 122.605 181.385 ;
        RECT 123.095 180.575 124.445 181.485 ;
        RECT 124.455 180.575 129.965 181.385 ;
        RECT 130.455 180.575 131.805 181.485 ;
        RECT 131.835 180.575 133.185 181.485 ;
        RECT 133.205 180.660 133.635 181.445 ;
        RECT 133.655 180.575 135.005 181.485 ;
        RECT 135.955 180.575 139.165 181.485 ;
        RECT 139.185 180.575 140.535 181.485 ;
        RECT 140.555 180.575 141.905 181.485 ;
        RECT 141.935 180.575 145.605 181.385 ;
        RECT 145.615 180.575 146.985 181.385 ;
        RECT 17.415 180.365 17.585 180.575 ;
        RECT 18.795 180.365 18.965 180.575 ;
        RECT 21.550 180.415 21.670 180.525 ;
        RECT 24.315 180.365 24.485 180.555 ;
        RECT 28.915 180.385 29.085 180.575 ;
        RECT 29.385 180.420 29.545 180.530 ;
        RECT 29.835 180.365 30.005 180.555 ;
        RECT 30.755 180.385 30.925 180.575 ;
        RECT 33.515 180.365 33.685 180.555 ;
        RECT 36.275 180.385 36.445 180.575 ;
        RECT 38.110 180.365 38.280 180.555 ;
        RECT 38.575 180.385 38.745 180.555 ;
        RECT 40.415 180.385 40.585 180.575 ;
        RECT 40.880 180.555 41.050 180.575 ;
        RECT 40.875 180.385 41.050 180.555 ;
        RECT 42.710 180.415 42.830 180.525 ;
        RECT 38.580 180.365 38.745 180.385 ;
        RECT 40.875 180.365 41.045 180.385 ;
        RECT 43.640 180.365 43.810 180.555 ;
        RECT 44.550 180.385 44.720 180.575 ;
        RECT 45.930 180.415 46.050 180.525 ;
        RECT 47.315 180.365 47.485 180.555 ;
        RECT 50.535 180.385 50.705 180.555 ;
        RECT 50.555 180.365 50.705 180.385 ;
        RECT 52.835 180.365 53.005 180.555 ;
        RECT 53.295 180.385 53.465 180.575 ;
        RECT 53.755 180.385 53.925 180.575 ;
        RECT 56.515 180.525 56.685 180.575 ;
        RECT 55.590 180.415 55.710 180.525 ;
        RECT 56.510 180.415 56.685 180.525 ;
        RECT 56.515 180.385 56.685 180.415 ;
        RECT 58.350 180.365 58.520 180.555 ;
        RECT 61.575 180.365 61.745 180.555 ;
        RECT 62.035 180.365 62.205 180.575 ;
        RECT 63.870 180.415 63.990 180.525 ;
        RECT 66.175 180.385 66.345 180.575 ;
        RECT 68.015 180.385 68.185 180.575 ;
        RECT 68.480 180.555 68.650 180.575 ;
        RECT 70.795 180.555 70.945 180.575 ;
        RECT 68.475 180.385 68.650 180.555 ;
        RECT 69.865 180.420 70.025 180.530 ;
        RECT 70.775 180.385 70.945 180.555 ;
        RECT 68.475 180.365 68.645 180.385 ;
        RECT 72.615 180.365 72.785 180.555 ;
        RECT 74.450 180.365 74.620 180.555 ;
        RECT 74.915 180.365 75.085 180.555 ;
        RECT 77.675 180.365 77.845 180.555 ;
        RECT 79.975 180.385 80.145 180.575 ;
        RECT 80.435 180.385 80.605 180.575 ;
        RECT 82.275 180.385 82.445 180.575 ;
        RECT 85.035 180.365 85.205 180.555 ;
        RECT 85.950 180.415 86.070 180.525 ;
        RECT 86.415 180.385 86.585 180.575 ;
        RECT 90.555 180.365 90.725 180.555 ;
        RECT 94.050 180.385 94.220 180.575 ;
        RECT 94.230 180.415 94.350 180.525 ;
        RECT 95.430 180.365 95.600 180.555 ;
        RECT 97.915 180.385 98.085 180.575 ;
        RECT 99.295 180.365 99.465 180.555 ;
        RECT 100.950 180.385 101.120 180.575 ;
        RECT 101.135 180.365 101.305 180.555 ;
        RECT 104.825 180.420 104.985 180.530 ;
        RECT 106.195 180.365 106.365 180.555 ;
        RECT 106.650 180.385 106.820 180.575 ;
        RECT 107.110 180.415 107.230 180.525 ;
        RECT 108.035 180.365 108.205 180.575 ;
        RECT 115.395 180.385 115.565 180.575 ;
        RECT 116.315 180.385 116.485 180.555 ;
        RECT 119.990 180.415 120.110 180.525 ;
        RECT 116.315 180.365 116.515 180.385 ;
        RECT 120.915 180.365 121.085 180.575 ;
        RECT 122.750 180.415 122.870 180.525 ;
        RECT 123.210 180.385 123.380 180.575 ;
        RECT 124.595 180.385 124.765 180.575 ;
        RECT 126.435 180.365 126.605 180.555 ;
        RECT 128.280 180.365 128.450 180.555 ;
        RECT 129.655 180.365 129.825 180.555 ;
        RECT 130.110 180.415 130.230 180.525 ;
        RECT 131.490 180.385 131.660 180.575 ;
        RECT 132.870 180.385 133.040 180.575 ;
        RECT 133.800 180.385 133.970 180.575 ;
        RECT 135.185 180.420 135.345 180.530 ;
        RECT 135.640 180.365 135.810 180.555 ;
        RECT 136.095 180.385 136.265 180.575 ;
        RECT 137.935 180.385 138.105 180.555 ;
        RECT 137.935 180.365 138.085 180.385 ;
        RECT 138.400 180.365 138.570 180.555 ;
        RECT 139.775 180.365 139.945 180.555 ;
        RECT 140.235 180.385 140.405 180.575 ;
        RECT 141.620 180.385 141.790 180.575 ;
        RECT 142.075 180.385 142.245 180.575 ;
        RECT 145.290 180.415 145.410 180.525 ;
        RECT 146.675 180.365 146.845 180.575 ;
        RECT 17.275 179.555 18.645 180.365 ;
        RECT 18.655 179.555 24.165 180.365 ;
        RECT 24.175 179.555 29.685 180.365 ;
        RECT 29.695 179.555 33.365 180.365 ;
        RECT 33.375 179.555 34.745 180.365 ;
        RECT 34.755 179.685 38.425 180.365 ;
        RECT 38.580 179.685 40.415 180.365 ;
        RECT 37.500 179.455 38.425 179.685 ;
        RECT 39.485 179.455 40.415 179.685 ;
        RECT 40.735 179.555 42.565 180.365 ;
        RECT 43.045 179.495 43.475 180.280 ;
        RECT 43.495 179.685 47.080 180.365 ;
        RECT 43.495 179.455 44.415 179.685 ;
        RECT 47.215 179.455 50.385 180.365 ;
        RECT 50.555 179.545 52.485 180.365 ;
        RECT 52.695 179.555 56.365 180.365 ;
        RECT 51.535 179.455 52.485 179.545 ;
        RECT 56.895 179.455 58.665 180.365 ;
        RECT 58.675 179.455 61.785 180.365 ;
        RECT 61.995 179.455 65.105 180.365 ;
        RECT 65.210 179.685 68.675 180.365 ;
        RECT 65.210 179.455 66.130 179.685 ;
        RECT 68.805 179.495 69.235 180.280 ;
        RECT 69.350 179.685 72.815 180.365 ;
        RECT 69.350 179.455 70.270 179.685 ;
        RECT 72.995 179.455 74.765 180.365 ;
        RECT 74.775 179.555 77.525 180.365 ;
        RECT 77.535 179.685 84.845 180.365 ;
        RECT 81.050 179.465 81.960 179.685 ;
        RECT 83.495 179.455 84.845 179.685 ;
        RECT 84.895 179.555 90.405 180.365 ;
        RECT 90.415 179.555 94.085 180.365 ;
        RECT 94.565 179.495 94.995 180.280 ;
        RECT 95.015 179.685 98.915 180.365 ;
        RECT 95.015 179.455 95.945 179.685 ;
        RECT 99.155 179.555 100.985 180.365 ;
        RECT 100.995 179.685 105.810 180.365 ;
        RECT 106.055 179.555 107.885 180.365 ;
        RECT 107.895 179.685 115.205 180.365 ;
        RECT 116.315 179.685 119.845 180.365 ;
        RECT 111.410 179.465 112.320 179.685 ;
        RECT 113.855 179.455 115.205 179.685 ;
        RECT 117.020 179.455 119.845 179.685 ;
        RECT 120.325 179.495 120.755 180.280 ;
        RECT 120.775 179.555 126.285 180.365 ;
        RECT 126.310 179.455 128.125 180.365 ;
        RECT 128.135 179.455 129.485 180.365 ;
        RECT 129.515 179.555 132.265 180.365 ;
        RECT 132.275 179.455 135.935 180.365 ;
        RECT 136.155 179.545 138.085 180.365 ;
        RECT 136.155 179.455 137.105 179.545 ;
        RECT 138.255 179.455 139.605 180.365 ;
        RECT 139.635 179.555 145.145 180.365 ;
        RECT 145.615 179.555 146.985 180.365 ;
      LAYER nwell ;
        RECT 17.080 176.335 147.180 179.165 ;
      LAYER pwell ;
        RECT 17.275 175.135 18.645 175.945 ;
        RECT 18.655 175.135 22.325 175.945 ;
        RECT 22.335 175.135 23.705 175.945 ;
        RECT 23.725 175.135 25.075 176.045 ;
        RECT 25.755 175.955 26.705 176.045 ;
        RECT 25.755 175.135 27.685 175.955 ;
        RECT 27.855 175.135 29.685 175.945 ;
        RECT 30.165 175.220 30.595 176.005 ;
        RECT 30.615 175.135 33.825 176.045 ;
        RECT 33.835 175.135 36.125 176.045 ;
        RECT 36.135 175.135 37.485 176.045 ;
        RECT 37.515 175.135 43.025 175.945 ;
        RECT 45.300 175.845 46.245 176.045 ;
        RECT 43.495 175.165 46.245 175.845 ;
        RECT 47.625 175.815 48.545 176.045 ;
        RECT 17.415 174.925 17.585 175.135 ;
        RECT 18.795 174.925 18.965 175.135 ;
        RECT 22.475 174.945 22.645 175.135 ;
        RECT 22.475 174.925 22.640 174.945 ;
        RECT 24.775 174.925 24.945 175.135 ;
        RECT 27.535 175.115 27.685 175.135 ;
        RECT 25.230 174.975 25.350 175.085 ;
        RECT 27.075 174.945 27.245 175.115 ;
        RECT 27.535 175.085 27.705 175.115 ;
        RECT 27.530 174.975 27.705 175.085 ;
        RECT 27.535 174.945 27.705 174.975 ;
        RECT 27.995 174.945 28.165 175.135 ;
        RECT 30.755 175.115 30.925 175.135 ;
        RECT 29.830 174.975 29.950 175.085 ;
        RECT 30.750 174.945 30.925 175.115 ;
        RECT 27.075 174.925 27.240 174.945 ;
        RECT 30.750 174.925 30.920 174.945 ;
        RECT 32.135 174.925 32.305 175.115 ;
        RECT 32.595 174.925 32.765 175.115 ;
        RECT 35.815 174.945 35.985 175.135 ;
        RECT 36.270 174.975 36.390 175.085 ;
        RECT 37.200 174.945 37.370 175.135 ;
        RECT 37.655 174.945 37.825 175.135 ;
        RECT 38.575 174.945 38.745 175.115 ;
        RECT 38.575 174.925 38.740 174.945 ;
        RECT 39.955 174.925 40.125 175.115 ;
        RECT 40.415 174.925 40.585 175.115 ;
        RECT 42.710 174.925 42.880 175.115 ;
        RECT 43.170 174.975 43.290 175.085 ;
        RECT 43.640 174.945 43.810 175.165 ;
        RECT 45.300 175.135 46.245 175.165 ;
        RECT 46.255 175.135 48.545 175.815 ;
        RECT 48.565 175.135 49.915 176.045 ;
        RECT 49.935 175.135 52.685 175.945 ;
        RECT 53.165 175.135 54.515 176.045 ;
        RECT 54.535 175.135 55.905 175.945 ;
        RECT 55.925 175.220 56.355 176.005 ;
        RECT 56.855 175.135 58.205 176.045 ;
        RECT 61.730 175.815 62.640 176.035 ;
        RECT 64.175 175.815 65.525 176.045 ;
        RECT 58.215 175.135 65.525 175.815 ;
        RECT 65.615 175.815 66.965 176.045 ;
        RECT 68.500 175.815 69.410 176.035 ;
        RECT 65.615 175.135 72.925 175.815 ;
        RECT 72.935 175.135 78.445 175.945 ;
        RECT 78.455 175.135 81.205 175.945 ;
        RECT 81.685 175.220 82.115 176.005 ;
        RECT 82.135 175.135 83.965 175.945 ;
        RECT 87.090 175.815 88.010 176.045 ;
        RECT 84.545 175.135 88.010 175.815 ;
        RECT 88.115 175.135 91.785 175.945 ;
        RECT 91.795 175.135 93.165 175.945 ;
        RECT 96.690 175.815 97.600 176.035 ;
        RECT 99.135 175.815 100.485 176.045 ;
        RECT 93.175 175.135 100.485 175.815 ;
        RECT 100.535 175.815 101.465 176.045 ;
        RECT 100.535 175.135 104.435 175.815 ;
        RECT 105.595 175.135 107.410 176.045 ;
        RECT 107.445 175.220 107.875 176.005 ;
        RECT 107.905 175.135 109.255 176.045 ;
        RECT 109.275 175.815 113.205 176.045 ;
        RECT 113.875 175.845 114.825 176.045 ;
        RECT 118.695 175.955 119.645 176.045 ;
        RECT 109.275 175.135 113.690 175.815 ;
        RECT 113.875 175.165 117.545 175.845 ;
        RECT 113.875 175.135 114.825 175.165 ;
        RECT 46.395 174.925 46.565 175.135 ;
        RECT 47.780 174.925 47.950 175.115 ;
        RECT 48.230 174.975 48.350 175.085 ;
        RECT 48.695 174.945 48.865 175.135 ;
        RECT 50.075 174.945 50.245 175.135 ;
        RECT 52.830 174.975 52.950 175.085 ;
        RECT 53.295 174.945 53.465 175.135 ;
        RECT 54.675 174.945 54.845 175.135 ;
        RECT 55.595 174.925 55.765 175.115 ;
        RECT 56.055 174.925 56.225 175.115 ;
        RECT 56.510 174.975 56.630 175.085 ;
        RECT 57.890 174.945 58.060 175.135 ;
        RECT 58.355 174.945 58.525 175.135 ;
        RECT 61.575 174.925 61.745 175.115 ;
        RECT 69.395 174.925 69.565 175.115 ;
        RECT 72.615 174.945 72.785 175.135 ;
        RECT 73.075 174.945 73.245 175.135 ;
        RECT 74.915 174.925 75.085 175.115 ;
        RECT 78.595 174.945 78.765 175.135 ;
        RECT 81.350 174.975 81.470 175.085 ;
        RECT 82.275 174.945 82.445 175.135 ;
        RECT 83.655 174.925 83.825 175.115 ;
        RECT 84.120 175.085 84.290 175.115 ;
        RECT 84.110 174.975 84.290 175.085 ;
        RECT 84.120 174.925 84.290 174.975 ;
        RECT 84.575 174.945 84.745 175.135 ;
        RECT 87.800 174.925 87.970 175.115 ;
        RECT 88.255 174.945 88.425 175.135 ;
        RECT 91.015 174.925 91.185 175.115 ;
        RECT 91.935 174.945 92.105 175.135 ;
        RECT 93.315 174.945 93.485 175.135 ;
        RECT 95.155 174.925 95.325 175.115 ;
        RECT 98.830 174.925 99.000 175.115 ;
        RECT 100.950 174.945 101.120 175.135 ;
        RECT 104.825 174.980 104.985 175.090 ;
        RECT 107.115 174.925 107.285 175.135 ;
        RECT 108.035 174.945 108.205 175.135 ;
        RECT 113.580 175.115 113.690 175.135 ;
        RECT 110.795 174.925 110.965 175.115 ;
        RECT 111.255 174.945 111.425 175.115 ;
        RECT 113.580 174.945 113.750 175.115 ;
        RECT 111.255 174.925 111.455 174.945 ;
        RECT 17.275 174.115 18.645 174.925 ;
        RECT 18.655 174.115 20.485 174.925 ;
        RECT 20.805 174.245 22.640 174.925 ;
        RECT 22.795 174.245 25.085 174.925 ;
        RECT 25.405 174.245 27.240 174.925 ;
        RECT 20.805 174.015 21.735 174.245 ;
        RECT 22.795 174.015 23.715 174.245 ;
        RECT 25.405 174.015 26.335 174.245 ;
        RECT 28.145 174.015 31.065 174.925 ;
        RECT 31.085 174.015 32.435 174.925 ;
        RECT 32.455 174.115 36.125 174.925 ;
        RECT 36.905 174.245 38.740 174.925 ;
        RECT 36.905 174.015 37.835 174.245 ;
        RECT 38.905 174.015 40.255 174.925 ;
        RECT 40.275 174.115 41.645 174.925 ;
        RECT 41.675 174.015 43.025 174.925 ;
        RECT 43.045 174.055 43.475 174.840 ;
        RECT 43.495 174.015 46.705 174.925 ;
        RECT 46.715 174.015 48.065 174.925 ;
        RECT 48.595 174.245 55.905 174.925 ;
        RECT 48.595 174.015 49.945 174.245 ;
        RECT 51.480 174.025 52.390 174.245 ;
        RECT 55.915 174.115 61.425 174.925 ;
        RECT 61.435 174.245 68.745 174.925 ;
        RECT 64.950 174.025 65.860 174.245 ;
        RECT 67.395 174.015 68.745 174.245 ;
        RECT 68.805 174.055 69.235 174.840 ;
        RECT 69.255 174.115 74.765 174.925 ;
        RECT 74.775 174.115 76.605 174.925 ;
        RECT 76.655 174.245 83.965 174.925 ;
        RECT 83.975 174.245 87.560 174.925 ;
        RECT 76.655 174.015 78.005 174.245 ;
        RECT 79.540 174.025 80.450 174.245 ;
        RECT 83.975 174.015 84.895 174.245 ;
        RECT 87.655 174.015 90.770 174.925 ;
        RECT 90.875 174.115 94.545 174.925 ;
        RECT 94.565 174.055 94.995 174.840 ;
        RECT 95.015 174.115 98.685 174.925 ;
        RECT 98.715 174.015 100.065 174.925 ;
        RECT 100.115 174.245 107.425 174.925 ;
        RECT 107.530 174.245 110.995 174.925 ;
        RECT 111.255 174.245 114.785 174.925 ;
        RECT 114.940 174.895 115.110 175.115 ;
        RECT 117.230 174.945 117.400 175.165 ;
        RECT 117.715 175.135 119.645 175.955 ;
        RECT 119.875 175.135 121.225 176.045 ;
        RECT 121.235 175.135 122.605 175.945 ;
        RECT 122.615 175.845 123.560 176.045 ;
        RECT 124.895 175.845 125.825 176.045 ;
        RECT 122.615 175.365 125.825 175.845 ;
        RECT 127.655 175.815 128.585 176.045 ;
        RECT 122.615 175.165 125.685 175.365 ;
        RECT 122.615 175.135 123.560 175.165 ;
        RECT 117.715 175.115 117.865 175.135 ;
        RECT 117.695 174.945 117.865 175.115 ;
        RECT 118.615 174.925 118.785 175.115 ;
        RECT 119.990 174.945 120.160 175.135 ;
        RECT 121.375 174.945 121.545 175.135 ;
        RECT 122.755 174.925 122.925 175.115 ;
        RECT 123.215 174.925 123.385 175.115 ;
        RECT 125.515 174.945 125.685 175.165 ;
        RECT 125.835 175.135 128.585 175.815 ;
        RECT 128.595 175.135 130.410 176.045 ;
        RECT 130.455 175.135 131.805 176.045 ;
        RECT 131.815 175.135 133.185 175.945 ;
        RECT 133.205 175.220 133.635 176.005 ;
        RECT 134.990 175.845 135.945 176.045 ;
        RECT 133.665 175.165 135.945 175.845 ;
        RECT 125.975 174.945 126.145 175.135 ;
        RECT 128.285 174.970 128.445 175.080 ;
        RECT 129.195 174.945 129.365 175.115 ;
        RECT 130.115 174.945 130.285 175.135 ;
        RECT 131.490 174.945 131.660 175.135 ;
        RECT 131.955 174.945 132.125 175.135 ;
        RECT 133.330 174.975 133.450 175.085 ;
        RECT 133.790 174.945 133.960 175.165 ;
        RECT 134.990 175.135 135.945 175.165 ;
        RECT 135.955 175.135 137.305 176.045 ;
        RECT 137.335 175.135 142.845 175.945 ;
        RECT 143.775 175.815 145.120 176.045 ;
        RECT 143.775 175.135 145.605 175.815 ;
        RECT 145.615 175.135 146.985 175.945 ;
        RECT 135.635 174.945 135.805 175.115 ;
        RECT 136.090 174.975 136.210 175.085 ;
        RECT 129.205 174.925 129.365 174.945 ;
        RECT 135.635 174.925 135.800 174.945 ;
        RECT 136.555 174.925 136.725 175.115 ;
        RECT 137.020 174.945 137.190 175.135 ;
        RECT 137.475 174.945 137.645 175.135 ;
        RECT 143.005 174.980 143.165 175.090 ;
        RECT 143.915 174.925 144.085 175.115 ;
        RECT 145.295 174.945 145.465 175.135 ;
        RECT 146.675 174.925 146.845 175.135 ;
        RECT 117.515 174.895 118.465 174.925 ;
        RECT 100.115 174.015 101.465 174.245 ;
        RECT 103.000 174.025 103.910 174.245 ;
        RECT 107.530 174.015 108.450 174.245 ;
        RECT 111.960 174.015 114.785 174.245 ;
        RECT 114.795 174.215 118.465 174.895 ;
        RECT 117.515 174.015 118.465 174.215 ;
        RECT 118.475 174.115 120.305 174.925 ;
        RECT 120.325 174.055 120.755 174.840 ;
        RECT 120.775 174.245 123.065 174.925 ;
        RECT 123.075 174.245 127.890 174.925 ;
        RECT 120.775 174.015 121.695 174.245 ;
        RECT 129.205 174.015 132.860 174.925 ;
        RECT 133.965 174.245 135.800 174.925 ;
        RECT 136.415 174.245 143.725 174.925 ;
        RECT 143.775 174.245 145.605 174.925 ;
        RECT 133.965 174.015 134.895 174.245 ;
        RECT 139.930 174.025 140.840 174.245 ;
        RECT 142.375 174.015 143.725 174.245 ;
        RECT 144.260 174.015 145.605 174.245 ;
        RECT 145.615 174.115 146.985 174.925 ;
      LAYER nwell ;
        RECT 17.080 170.895 147.180 173.725 ;
      LAYER pwell ;
        RECT 17.275 169.695 18.645 170.505 ;
        RECT 22.630 170.375 23.540 170.595 ;
        RECT 25.075 170.375 26.425 170.605 ;
        RECT 19.115 169.695 26.425 170.375 ;
        RECT 26.475 169.695 27.825 170.605 ;
        RECT 29.225 170.375 30.145 170.605 ;
        RECT 27.855 169.695 30.145 170.375 ;
        RECT 30.165 169.780 30.595 170.565 ;
        RECT 34.130 170.375 35.040 170.595 ;
        RECT 36.575 170.375 37.925 170.605 ;
        RECT 39.115 170.515 40.065 170.605 ;
        RECT 30.615 169.695 37.925 170.375 ;
        RECT 38.135 169.695 40.065 170.515 ;
        RECT 43.165 170.375 44.095 170.605 ;
        RECT 45.785 170.375 46.705 170.605 ;
        RECT 40.275 169.695 42.105 170.375 ;
        RECT 42.260 169.695 44.095 170.375 ;
        RECT 44.415 169.695 46.705 170.375 ;
        RECT 46.815 169.695 49.925 170.605 ;
        RECT 51.075 170.515 52.025 170.605 ;
        RECT 50.095 169.695 52.025 170.515 ;
        RECT 52.235 169.695 55.905 170.505 ;
        RECT 55.925 169.780 56.355 170.565 ;
        RECT 56.375 169.695 61.885 170.505 ;
        RECT 61.895 169.695 67.405 170.505 ;
        RECT 67.415 169.695 72.925 170.505 ;
        RECT 72.935 169.695 78.445 170.505 ;
        RECT 78.455 169.695 81.205 170.505 ;
        RECT 81.685 169.780 82.115 170.565 ;
        RECT 82.595 169.925 85.345 170.605 ;
        RECT 85.355 170.405 86.285 170.605 ;
        RECT 87.615 170.405 88.565 170.605 ;
        RECT 85.355 169.925 88.565 170.405 ;
        RECT 82.735 169.695 85.345 169.925 ;
        RECT 85.500 169.725 88.565 169.925 ;
        RECT 17.415 169.485 17.585 169.695 ;
        RECT 18.795 169.645 18.965 169.675 ;
        RECT 18.790 169.535 18.965 169.645 ;
        RECT 18.795 169.485 18.965 169.535 ;
        RECT 19.255 169.505 19.425 169.695 ;
        RECT 22.015 169.485 22.185 169.675 ;
        RECT 22.475 169.485 22.645 169.675 ;
        RECT 27.540 169.505 27.710 169.695 ;
        RECT 27.995 169.505 28.165 169.695 ;
        RECT 29.835 169.485 30.005 169.675 ;
        RECT 30.755 169.505 30.925 169.695 ;
        RECT 38.135 169.675 38.285 169.695 ;
        RECT 32.135 169.485 32.305 169.675 ;
        RECT 34.890 169.535 35.010 169.645 ;
        RECT 35.355 169.485 35.525 169.675 ;
        RECT 38.115 169.505 38.285 169.675 ;
        RECT 41.795 169.505 41.965 169.695 ;
        RECT 42.260 169.675 42.425 169.695 ;
        RECT 42.255 169.505 42.425 169.675 ;
        RECT 42.710 169.535 42.830 169.645 ;
        RECT 43.635 169.485 43.805 169.675 ;
        RECT 44.555 169.505 44.725 169.695 ;
        RECT 46.855 169.505 47.025 169.695 ;
        RECT 50.095 169.675 50.245 169.695 ;
        RECT 50.075 169.505 50.245 169.675 ;
        RECT 51.915 169.485 52.085 169.675 ;
        RECT 52.375 169.485 52.545 169.695 ;
        RECT 56.515 169.505 56.685 169.695 ;
        RECT 57.895 169.485 58.065 169.675 ;
        RECT 61.570 169.535 61.690 169.645 ;
        RECT 62.035 169.505 62.205 169.695 ;
        RECT 62.955 169.485 63.125 169.675 ;
        RECT 63.425 169.530 63.585 169.640 ;
        RECT 67.555 169.485 67.725 169.695 ;
        RECT 68.025 169.530 68.185 169.640 ;
        RECT 69.395 169.485 69.565 169.675 ;
        RECT 73.075 169.505 73.245 169.695 ;
        RECT 74.915 169.485 75.085 169.675 ;
        RECT 78.595 169.505 78.765 169.695 ;
        RECT 79.515 169.485 79.685 169.675 ;
        RECT 81.350 169.535 81.470 169.645 ;
        RECT 82.270 169.535 82.390 169.645 ;
        RECT 82.735 169.505 82.905 169.695 ;
        RECT 83.195 169.485 83.365 169.675 ;
        RECT 85.500 169.505 85.670 169.725 ;
        RECT 87.630 169.695 88.565 169.725 ;
        RECT 88.575 169.695 89.925 170.605 ;
        RECT 93.930 170.375 94.840 170.595 ;
        RECT 96.375 170.375 97.725 170.605 ;
        RECT 102.930 170.375 103.850 170.605 ;
        RECT 90.415 169.695 97.725 170.375 ;
        RECT 98.010 169.695 102.825 170.375 ;
        RECT 102.930 169.695 106.395 170.375 ;
        RECT 107.445 169.780 107.875 170.565 ;
        RECT 107.945 169.695 111.105 170.605 ;
        RECT 111.115 170.405 112.045 170.605 ;
        RECT 113.375 170.405 114.325 170.605 ;
        RECT 111.115 169.925 114.325 170.405 ;
        RECT 111.260 169.725 114.325 169.925 ;
        RECT 89.640 169.675 89.810 169.695 ;
        RECT 89.635 169.505 89.810 169.675 ;
        RECT 90.555 169.675 90.725 169.695 ;
        RECT 90.090 169.535 90.210 169.645 ;
        RECT 90.555 169.505 90.730 169.675 ;
        RECT 95.155 169.505 95.325 169.675 ;
        RECT 97.450 169.535 97.570 169.645 ;
        RECT 89.635 169.485 89.805 169.505 ;
        RECT 90.560 169.485 90.730 169.505 ;
        RECT 95.160 169.485 95.325 169.505 ;
        RECT 101.595 169.485 101.765 169.675 ;
        RECT 102.515 169.505 102.685 169.695 ;
        RECT 105.275 169.485 105.445 169.675 ;
        RECT 106.195 169.505 106.365 169.695 ;
        RECT 106.665 169.540 106.825 169.650 ;
        RECT 108.035 169.505 108.205 169.695 ;
        RECT 108.495 169.485 108.665 169.675 ;
        RECT 108.965 169.530 109.125 169.640 ;
        RECT 111.260 169.505 111.430 169.725 ;
        RECT 113.390 169.695 114.325 169.725 ;
        RECT 114.415 169.695 116.625 170.605 ;
        RECT 117.565 169.695 120.295 170.605 ;
        RECT 120.785 169.695 123.515 170.605 ;
        RECT 124.195 169.695 126.285 170.505 ;
        RECT 126.445 169.695 130.100 170.605 ;
        RECT 130.745 170.375 131.675 170.605 ;
        RECT 130.745 169.695 132.580 170.375 ;
        RECT 133.205 169.780 133.635 170.565 ;
        RECT 134.990 170.405 135.945 170.605 ;
        RECT 133.665 169.725 135.945 170.405 ;
        RECT 115.390 169.485 115.560 169.675 ;
        RECT 115.855 169.485 116.025 169.675 ;
        RECT 116.310 169.505 116.480 169.695 ;
        RECT 116.785 169.540 116.945 169.650 ;
        RECT 117.695 169.505 117.865 169.695 ;
        RECT 120.915 169.675 121.085 169.695 ;
        RECT 118.160 169.485 118.330 169.675 ;
        RECT 118.610 169.535 118.730 169.645 ;
        RECT 119.070 169.485 119.240 169.675 ;
        RECT 120.450 169.535 120.570 169.645 ;
        RECT 120.910 169.505 121.085 169.675 ;
        RECT 17.275 168.675 18.645 169.485 ;
        RECT 18.655 168.675 20.025 169.485 ;
        RECT 20.035 168.805 22.325 169.485 ;
        RECT 22.335 168.805 29.645 169.485 ;
        RECT 29.695 168.805 31.985 169.485 ;
        RECT 20.035 168.575 20.955 168.805 ;
        RECT 25.850 168.585 26.760 168.805 ;
        RECT 28.295 168.575 29.645 168.805 ;
        RECT 31.065 168.575 31.985 168.805 ;
        RECT 31.995 168.675 34.745 169.485 ;
        RECT 35.215 168.805 42.525 169.485 ;
        RECT 38.730 168.585 39.640 168.805 ;
        RECT 41.175 168.575 42.525 168.805 ;
        RECT 43.045 168.615 43.475 169.400 ;
        RECT 43.495 168.675 44.865 169.485 ;
        RECT 44.915 168.805 52.225 169.485 ;
        RECT 44.915 168.575 46.265 168.805 ;
        RECT 47.800 168.585 48.710 168.805 ;
        RECT 52.235 168.675 57.745 169.485 ;
        RECT 57.755 168.675 61.425 169.485 ;
        RECT 61.905 168.575 63.255 169.485 ;
        RECT 64.290 168.805 67.755 169.485 ;
        RECT 64.290 168.575 65.210 168.805 ;
        RECT 68.805 168.615 69.235 169.400 ;
        RECT 69.255 168.675 74.765 169.485 ;
        RECT 74.775 168.675 78.445 169.485 ;
        RECT 79.485 168.805 82.950 169.485 ;
        RECT 82.030 168.575 82.950 168.805 ;
        RECT 83.055 168.675 86.725 169.485 ;
        RECT 88.105 169.455 89.945 169.485 ;
        RECT 86.780 168.805 89.945 169.455 ;
        RECT 86.780 168.775 89.460 168.805 ;
        RECT 88.105 168.575 89.460 168.775 ;
        RECT 90.415 168.575 94.305 169.485 ;
        RECT 94.565 168.615 94.995 169.400 ;
        RECT 95.160 168.805 96.995 169.485 ;
        RECT 96.065 168.575 96.995 168.805 ;
        RECT 97.775 168.575 101.905 169.485 ;
        RECT 102.010 168.805 105.475 169.485 ;
        RECT 102.010 168.575 102.930 168.805 ;
        RECT 105.595 168.575 108.805 169.485 ;
        RECT 109.995 168.575 115.705 169.485 ;
        RECT 115.725 168.575 117.075 169.485 ;
        RECT 117.095 168.575 118.445 169.485 ;
        RECT 118.955 168.575 120.305 169.485 ;
        RECT 120.910 169.455 121.080 169.505 ;
        RECT 123.215 169.485 123.385 169.675 ;
        RECT 125.975 169.505 126.145 169.695 ;
        RECT 126.445 169.675 126.605 169.695 ;
        RECT 132.415 169.675 132.580 169.695 ;
        RECT 126.435 169.505 126.605 169.675 ;
        RECT 131.490 169.485 131.660 169.675 ;
        RECT 131.955 169.485 132.125 169.675 ;
        RECT 132.415 169.505 132.585 169.675 ;
        RECT 132.870 169.535 132.990 169.645 ;
        RECT 133.790 169.505 133.960 169.725 ;
        RECT 134.990 169.695 135.945 169.725 ;
        RECT 135.955 169.695 137.325 170.505 ;
        RECT 137.335 170.375 138.265 170.605 ;
        RECT 141.570 170.375 142.490 170.605 ;
        RECT 137.335 169.695 141.235 170.375 ;
        RECT 141.570 169.695 145.035 170.375 ;
        RECT 145.615 169.695 146.985 170.505 ;
        RECT 135.170 169.535 135.290 169.645 ;
        RECT 135.635 169.485 135.805 169.675 ;
        RECT 136.095 169.505 136.265 169.695 ;
        RECT 137.750 169.505 137.920 169.695 ;
        RECT 143.005 169.530 143.165 169.640 ;
        RECT 143.915 169.485 144.085 169.675 ;
        RECT 144.835 169.505 145.005 169.695 ;
        RECT 145.290 169.535 145.410 169.645 ;
        RECT 146.675 169.485 146.845 169.695 ;
        RECT 122.110 169.455 123.065 169.485 ;
        RECT 120.325 168.615 120.755 169.400 ;
        RECT 120.785 168.775 123.065 169.455 ;
        RECT 123.075 168.805 127.890 169.485 ;
        RECT 122.110 168.575 123.065 168.775 ;
        RECT 128.330 168.575 131.805 169.485 ;
        RECT 131.815 168.575 135.025 169.485 ;
        RECT 135.495 168.805 142.805 169.485 ;
        RECT 143.775 168.805 145.605 169.485 ;
        RECT 139.010 168.585 139.920 168.805 ;
        RECT 141.455 168.575 142.805 168.805 ;
        RECT 144.260 168.575 145.605 168.805 ;
        RECT 145.615 168.675 146.985 169.485 ;
      LAYER nwell ;
        RECT 17.080 165.455 147.180 168.285 ;
      LAYER pwell ;
        RECT 17.275 164.255 18.645 165.065 ;
        RECT 18.655 164.255 24.165 165.065 ;
        RECT 24.175 164.255 29.685 165.065 ;
        RECT 30.165 164.340 30.595 165.125 ;
        RECT 30.615 164.255 36.125 165.065 ;
        RECT 36.595 164.935 37.515 165.165 ;
        RECT 36.595 164.255 38.885 164.935 ;
        RECT 38.895 164.255 44.405 165.065 ;
        RECT 44.415 164.255 49.925 165.065 ;
        RECT 49.935 164.255 55.445 165.065 ;
        RECT 55.925 164.340 56.355 165.125 ;
        RECT 56.375 164.255 58.205 165.065 ;
        RECT 61.330 164.935 62.250 165.165 ;
        RECT 58.785 164.255 62.250 164.935 ;
        RECT 62.365 164.255 65.095 165.165 ;
        RECT 66.345 164.935 67.275 165.165 ;
        RECT 66.345 164.255 68.180 164.935 ;
        RECT 68.335 164.255 70.165 164.935 ;
        RECT 70.175 164.255 71.525 165.165 ;
        RECT 75.070 164.935 75.980 165.155 ;
        RECT 77.515 164.935 78.865 165.165 ;
        RECT 71.555 164.255 78.865 164.935 ;
        RECT 78.915 164.935 79.835 165.165 ;
        RECT 78.915 164.255 81.205 164.935 ;
        RECT 81.685 164.340 82.115 165.125 ;
        RECT 82.135 164.255 87.645 165.065 ;
        RECT 87.655 164.255 93.165 165.065 ;
        RECT 93.175 164.255 96.845 165.065 ;
        RECT 97.315 164.255 98.665 165.165 ;
        RECT 98.695 164.255 104.205 165.065 ;
        RECT 104.215 164.255 106.965 165.065 ;
        RECT 107.445 164.340 107.875 165.125 ;
        RECT 107.895 164.255 111.565 165.065 ;
        RECT 114.690 164.935 115.610 165.165 ;
        RECT 112.145 164.255 115.610 164.935 ;
        RECT 115.715 164.255 119.215 165.165 ;
        RECT 119.395 164.255 121.225 165.065 ;
        RECT 121.715 164.255 123.065 165.165 ;
        RECT 127.805 164.935 128.735 165.165 ;
        RECT 123.480 164.255 125.905 164.935 ;
        RECT 126.900 164.255 128.735 164.935 ;
        RECT 129.055 164.255 131.805 165.165 ;
        RECT 131.815 164.255 133.185 165.065 ;
        RECT 133.205 164.340 133.635 165.125 ;
        RECT 133.655 164.255 135.485 165.165 ;
        RECT 135.495 164.255 136.865 165.035 ;
        RECT 136.875 164.935 137.805 165.165 ;
        RECT 141.110 164.935 142.030 165.165 ;
        RECT 136.875 164.255 140.775 164.935 ;
        RECT 141.110 164.255 144.575 164.935 ;
        RECT 145.615 164.255 146.985 165.065 ;
        RECT 17.415 164.045 17.585 164.255 ;
        RECT 18.795 164.045 18.965 164.255 ;
        RECT 20.635 164.045 20.805 164.235 ;
        RECT 24.315 164.065 24.485 164.255 ;
        RECT 26.155 164.045 26.325 164.235 ;
        RECT 29.830 164.095 29.950 164.205 ;
        RECT 30.755 164.065 30.925 164.255 ;
        RECT 31.675 164.045 31.845 164.235 ;
        RECT 36.270 164.095 36.390 164.205 ;
        RECT 37.195 164.045 37.365 164.235 ;
        RECT 38.575 164.065 38.745 164.255 ;
        RECT 39.035 164.065 39.205 164.255 ;
        RECT 42.710 164.095 42.830 164.205 ;
        RECT 43.635 164.045 43.805 164.235 ;
        RECT 44.555 164.065 44.725 164.255 ;
        RECT 49.155 164.045 49.325 164.235 ;
        RECT 50.075 164.065 50.245 164.255 ;
        RECT 54.675 164.045 54.845 164.235 ;
        RECT 55.590 164.095 55.710 164.205 ;
        RECT 56.055 164.065 56.225 164.235 ;
        RECT 56.515 164.065 56.685 164.255 ;
        RECT 58.350 164.095 58.470 164.205 ;
        RECT 56.205 164.045 56.225 164.065 ;
        RECT 58.815 164.045 58.985 164.255 ;
        RECT 62.495 164.065 62.665 164.255 ;
        RECT 68.015 164.235 68.180 164.255 ;
        RECT 65.265 164.100 65.425 164.210 ;
        RECT 66.175 164.045 66.345 164.235 ;
        RECT 68.015 164.065 68.185 164.235 ;
        RECT 69.855 164.065 70.025 164.255 ;
        RECT 70.320 164.065 70.490 164.255 ;
        RECT 71.695 164.045 71.865 164.255 ;
        RECT 72.155 164.045 72.325 164.235 ;
        RECT 75.835 164.045 76.005 164.235 ;
        RECT 80.895 164.065 81.065 164.255 ;
        RECT 81.350 164.095 81.470 164.205 ;
        RECT 82.275 164.065 82.445 164.255 ;
        RECT 86.415 164.045 86.585 164.235 ;
        RECT 86.880 164.045 87.050 164.235 ;
        RECT 87.795 164.065 87.965 164.255 ;
        RECT 89.185 164.090 89.345 164.200 ;
        RECT 90.095 164.065 90.265 164.235 ;
        RECT 93.315 164.045 93.485 164.255 ;
        RECT 95.155 164.045 95.325 164.235 ;
        RECT 96.990 164.095 97.110 164.205 ;
        RECT 97.460 164.065 97.630 164.255 ;
        RECT 98.835 164.065 99.005 164.255 ;
        RECT 100.675 164.045 100.845 164.235 ;
        RECT 102.510 164.095 102.630 164.205 ;
        RECT 102.975 164.045 103.145 164.235 ;
        RECT 104.355 164.065 104.525 164.255 ;
        RECT 107.110 164.095 107.230 164.205 ;
        RECT 108.035 164.065 108.205 164.255 ;
        RECT 110.345 164.090 110.505 164.200 ;
        RECT 111.710 164.095 111.830 164.205 ;
        RECT 112.175 164.065 112.345 164.255 ;
        RECT 119.080 164.235 119.215 164.255 ;
        RECT 114.015 164.045 114.185 164.235 ;
        RECT 17.275 163.235 18.645 164.045 ;
        RECT 18.655 163.365 20.485 164.045 ;
        RECT 19.140 163.135 20.485 163.365 ;
        RECT 20.495 163.235 26.005 164.045 ;
        RECT 26.015 163.235 31.525 164.045 ;
        RECT 31.535 163.235 37.045 164.045 ;
        RECT 37.055 163.235 42.565 164.045 ;
        RECT 43.045 163.175 43.475 163.960 ;
        RECT 43.495 163.235 49.005 164.045 ;
        RECT 49.015 163.235 54.525 164.045 ;
        RECT 54.535 163.235 55.905 164.045 ;
        RECT 56.205 163.365 58.655 164.045 ;
        RECT 58.675 163.365 65.985 164.045 ;
        RECT 66.035 163.365 68.785 164.045 ;
        RECT 56.695 163.135 58.655 163.365 ;
        RECT 62.190 163.145 63.100 163.365 ;
        RECT 64.635 163.135 65.985 163.365 ;
        RECT 67.855 163.135 68.785 163.365 ;
        RECT 68.805 163.175 69.235 163.960 ;
        RECT 69.255 163.135 72.005 164.045 ;
        RECT 72.125 163.365 75.590 164.045 ;
        RECT 75.695 163.365 83.005 164.045 ;
        RECT 74.670 163.135 75.590 163.365 ;
        RECT 79.210 163.145 80.120 163.365 ;
        RECT 81.655 163.135 83.005 163.365 ;
        RECT 83.150 163.365 86.615 164.045 ;
        RECT 86.735 163.365 89.010 164.045 ;
        RECT 90.360 163.365 92.785 164.045 ;
        RECT 83.150 163.135 84.070 163.365 ;
        RECT 87.640 163.135 89.010 163.365 ;
        RECT 93.175 163.235 94.545 164.045 ;
        RECT 94.565 163.175 94.995 163.960 ;
        RECT 95.015 163.235 100.525 164.045 ;
        RECT 100.535 163.235 102.365 164.045 ;
        RECT 102.835 163.365 110.145 164.045 ;
        RECT 106.350 163.145 107.260 163.365 ;
        RECT 108.795 163.135 110.145 163.365 ;
        RECT 111.115 163.135 114.325 164.045 ;
        RECT 114.335 164.015 115.290 164.045 ;
        RECT 116.320 164.015 116.490 164.235 ;
        RECT 116.775 164.045 116.945 164.235 ;
        RECT 118.155 164.065 118.325 164.235 ;
        RECT 119.080 164.065 119.250 164.235 ;
        RECT 119.535 164.065 119.705 164.255 ;
        RECT 118.160 164.045 118.325 164.065 ;
        RECT 120.915 164.045 121.085 164.235 ;
        RECT 121.370 164.095 121.490 164.205 ;
        RECT 122.750 164.065 122.920 164.255 ;
        RECT 126.900 164.235 127.065 164.255 ;
        RECT 123.215 164.065 123.385 164.235 ;
        RECT 124.135 164.045 124.305 164.235 ;
        RECT 126.430 164.095 126.550 164.205 ;
        RECT 126.895 164.065 127.065 164.235 ;
        RECT 129.655 164.045 129.825 164.235 ;
        RECT 131.495 164.065 131.665 164.255 ;
        RECT 131.955 164.065 132.125 164.255 ;
        RECT 132.415 164.045 132.585 164.235 ;
        RECT 134.255 164.045 134.425 164.235 ;
        RECT 134.990 164.045 135.160 164.235 ;
        RECT 135.170 164.065 135.340 164.255 ;
        RECT 135.635 164.065 135.805 164.255 ;
        RECT 137.290 164.065 137.460 164.255 ;
        RECT 142.075 164.045 142.245 164.235 ;
        RECT 142.535 164.045 142.705 164.235 ;
        RECT 143.915 164.045 144.085 164.235 ;
        RECT 144.375 164.065 144.545 164.255 ;
        RECT 144.845 164.100 145.005 164.210 ;
        RECT 146.675 164.045 146.845 164.255 ;
        RECT 114.335 163.335 116.615 164.015 ;
        RECT 114.335 163.135 115.290 163.335 ;
        RECT 116.645 163.135 117.995 164.045 ;
        RECT 118.160 163.365 119.995 164.045 ;
        RECT 119.065 163.135 119.995 163.365 ;
        RECT 120.325 163.175 120.755 163.960 ;
        RECT 120.775 163.135 123.985 164.045 ;
        RECT 123.995 163.235 129.505 164.045 ;
        RECT 129.515 163.265 130.885 164.045 ;
        RECT 130.895 163.365 132.725 164.045 ;
        RECT 132.735 163.365 134.565 164.045 ;
        RECT 134.575 163.365 138.475 164.045 ;
        RECT 138.810 163.365 142.275 164.045 ;
        RECT 130.895 163.135 132.240 163.365 ;
        RECT 132.735 163.135 134.080 163.365 ;
        RECT 134.575 163.135 135.505 163.365 ;
        RECT 138.810 163.135 139.730 163.365 ;
        RECT 142.395 163.265 143.765 164.045 ;
        RECT 143.775 163.365 145.605 164.045 ;
        RECT 144.260 163.135 145.605 163.365 ;
        RECT 145.615 163.235 146.985 164.045 ;
      LAYER nwell ;
        RECT 17.080 160.015 147.180 162.845 ;
      LAYER pwell ;
        RECT 17.275 158.815 18.645 159.625 ;
        RECT 18.655 158.815 24.165 159.625 ;
        RECT 24.175 158.815 29.685 159.625 ;
        RECT 30.165 158.900 30.595 159.685 ;
        RECT 30.615 158.815 33.365 159.625 ;
        RECT 34.145 159.495 35.075 159.725 ;
        RECT 36.135 159.495 37.055 159.725 ;
        RECT 34.145 158.815 35.980 159.495 ;
        RECT 36.135 158.815 38.425 159.495 ;
        RECT 38.435 158.815 40.265 159.725 ;
        RECT 40.275 158.815 43.025 159.725 ;
        RECT 43.035 158.815 46.705 159.625 ;
        RECT 48.085 159.495 49.005 159.725 ;
        RECT 46.715 158.815 49.005 159.495 ;
        RECT 49.015 158.815 54.525 159.625 ;
        RECT 54.535 158.815 55.885 159.725 ;
        RECT 55.925 158.900 56.355 159.685 ;
        RECT 57.745 159.495 58.665 159.725 ;
        RECT 62.190 159.495 63.100 159.715 ;
        RECT 64.635 159.495 65.985 159.725 ;
        RECT 56.375 158.815 58.665 159.495 ;
        RECT 58.675 158.815 65.985 159.495 ;
        RECT 66.045 158.815 68.775 159.725 ;
        RECT 68.795 158.815 70.145 159.725 ;
        RECT 70.730 159.495 71.650 159.725 ;
        RECT 77.830 159.495 78.740 159.715 ;
        RECT 80.275 159.495 81.625 159.725 ;
        RECT 70.730 158.815 74.195 159.495 ;
        RECT 74.315 158.815 81.625 159.495 ;
        RECT 81.685 158.900 82.115 159.685 ;
        RECT 82.135 158.815 83.485 159.725 ;
        RECT 83.515 158.815 85.345 159.625 ;
        RECT 85.370 158.815 87.185 159.725 ;
        RECT 87.685 159.525 89.065 159.725 ;
        RECT 87.685 158.845 90.390 159.525 ;
        RECT 93.930 159.495 94.840 159.715 ;
        RECT 96.375 159.495 97.725 159.725 ;
        RECT 87.685 158.815 89.065 158.845 ;
        RECT 17.415 158.605 17.585 158.815 ;
        RECT 18.795 158.605 18.965 158.815 ;
        RECT 24.315 158.605 24.485 158.815 ;
        RECT 29.830 158.760 29.950 158.765 ;
        RECT 29.830 158.655 30.005 158.760 ;
        RECT 29.845 158.650 30.005 158.655 ;
        RECT 30.755 158.625 30.925 158.815 ;
        RECT 35.815 158.795 35.980 158.815 ;
        RECT 31.680 158.605 31.850 158.795 ;
        RECT 32.135 158.605 32.305 158.795 ;
        RECT 33.510 158.655 33.630 158.765 ;
        RECT 34.435 158.605 34.605 158.795 ;
        RECT 35.815 158.625 35.985 158.795 ;
        RECT 38.115 158.625 38.285 158.815 ;
        RECT 39.950 158.625 40.120 158.815 ;
        RECT 41.795 158.605 41.965 158.795 ;
        RECT 42.715 158.625 42.885 158.815 ;
        RECT 43.175 158.625 43.345 158.815 ;
        RECT 43.635 158.605 43.805 158.795 ;
        RECT 45.475 158.605 45.645 158.795 ;
        RECT 46.855 158.625 47.025 158.815 ;
        RECT 48.695 158.605 48.865 158.795 ;
        RECT 49.155 158.625 49.325 158.815 ;
        RECT 50.080 158.605 50.250 158.795 ;
        RECT 54.680 158.625 54.850 158.815 ;
        RECT 56.515 158.795 56.685 158.815 ;
        RECT 55.135 158.605 55.305 158.795 ;
        RECT 55.605 158.650 55.765 158.760 ;
        RECT 56.515 158.625 56.690 158.795 ;
        RECT 58.815 158.625 58.985 158.815 ;
        RECT 60.205 158.650 60.365 158.760 ;
        RECT 56.520 158.605 56.690 158.625 ;
        RECT 61.115 158.605 61.285 158.795 ;
        RECT 66.175 158.625 66.345 158.815 ;
        RECT 69.860 158.795 70.030 158.815 ;
        RECT 66.175 158.605 66.340 158.625 ;
        RECT 66.635 158.605 66.805 158.795 ;
        RECT 68.470 158.655 68.590 158.765 ;
        RECT 69.390 158.655 69.510 158.765 ;
        RECT 69.855 158.625 70.030 158.795 ;
        RECT 70.310 158.655 70.430 158.765 ;
        RECT 73.995 158.625 74.165 158.815 ;
        RECT 74.455 158.625 74.625 158.815 ;
        RECT 69.855 158.605 70.025 158.625 ;
        RECT 77.215 158.605 77.385 158.795 ;
        RECT 79.970 158.655 80.090 158.765 ;
        RECT 80.435 158.605 80.605 158.795 ;
        RECT 82.280 158.625 82.450 158.815 ;
        RECT 83.655 158.625 83.825 158.815 ;
        RECT 85.495 158.625 85.665 158.815 ;
        RECT 87.330 158.655 87.450 158.765 ;
        RECT 89.635 158.605 89.805 158.795 ;
        RECT 90.095 158.625 90.265 158.845 ;
        RECT 90.415 158.815 97.725 159.495 ;
        RECT 98.735 159.495 100.085 159.725 ;
        RECT 101.620 159.495 102.530 159.715 ;
        RECT 98.735 158.815 106.045 159.495 ;
        RECT 106.055 158.815 107.425 159.625 ;
        RECT 107.445 158.900 107.875 159.685 ;
        RECT 107.895 159.495 108.825 159.725 ;
        RECT 107.895 158.815 111.795 159.495 ;
        RECT 112.035 158.815 113.385 159.725 ;
        RECT 113.415 158.815 118.925 159.625 ;
        RECT 118.955 158.815 120.305 159.725 ;
        RECT 120.315 158.815 122.145 159.625 ;
        RECT 122.625 158.815 123.975 159.725 ;
        RECT 125.205 158.815 128.125 159.725 ;
        RECT 128.135 158.815 129.485 159.725 ;
        RECT 129.515 158.815 133.185 159.625 ;
        RECT 133.205 158.900 133.635 159.685 ;
        RECT 137.170 159.495 138.080 159.715 ;
        RECT 139.615 159.495 140.965 159.725 ;
        RECT 133.655 158.815 140.965 159.495 ;
        RECT 141.015 159.495 141.945 159.725 ;
        RECT 141.015 158.815 144.915 159.495 ;
        RECT 145.615 158.815 146.985 159.625 ;
        RECT 90.555 158.625 90.725 158.815 ;
        RECT 93.315 158.605 93.485 158.795 ;
        RECT 95.430 158.605 95.600 158.795 ;
        RECT 97.925 158.660 98.085 158.770 ;
        RECT 99.570 158.605 99.740 158.795 ;
        RECT 104.355 158.605 104.525 158.795 ;
        RECT 105.090 158.605 105.260 158.795 ;
        RECT 105.735 158.625 105.905 158.815 ;
        RECT 106.195 158.625 106.365 158.815 ;
        RECT 108.310 158.625 108.480 158.815 ;
        RECT 108.955 158.605 109.125 158.795 ;
        RECT 110.795 158.605 110.965 158.795 ;
        RECT 112.180 158.625 112.350 158.815 ;
        RECT 113.555 158.625 113.725 158.815 ;
        RECT 114.480 158.605 114.650 158.795 ;
        RECT 117.690 158.605 117.860 158.795 ;
        RECT 118.160 158.605 118.330 158.795 ;
        RECT 119.070 158.625 119.240 158.815 ;
        RECT 119.990 158.655 120.110 158.765 ;
        RECT 120.455 158.625 120.625 158.815 ;
        RECT 120.910 158.655 121.030 158.765 ;
        RECT 122.290 158.655 122.410 158.765 ;
        RECT 122.755 158.625 122.925 158.815 ;
        RECT 124.130 158.770 124.300 158.795 ;
        RECT 124.130 158.660 124.305 158.770 ;
        RECT 124.130 158.605 124.300 158.660 ;
        RECT 124.590 158.605 124.760 158.795 ;
        RECT 125.985 158.650 126.145 158.760 ;
        RECT 126.895 158.625 127.065 158.795 ;
        RECT 127.810 158.625 127.980 158.815 ;
        RECT 129.200 158.795 129.370 158.815 ;
        RECT 129.195 158.625 129.370 158.795 ;
        RECT 129.655 158.625 129.825 158.815 ;
        RECT 126.900 158.605 127.065 158.625 ;
        RECT 129.195 158.605 129.365 158.625 ;
        RECT 132.415 158.605 132.585 158.795 ;
        RECT 133.795 158.625 133.965 158.815 ;
        RECT 134.255 158.605 134.425 158.795 ;
        RECT 141.430 158.625 141.600 158.815 ;
        RECT 141.890 158.605 142.060 158.795 ;
        RECT 145.290 158.655 145.410 158.765 ;
        RECT 146.675 158.605 146.845 158.815 ;
        RECT 17.275 157.795 18.645 158.605 ;
        RECT 18.655 157.795 24.165 158.605 ;
        RECT 24.175 157.795 29.685 158.605 ;
        RECT 30.615 157.695 31.965 158.605 ;
        RECT 31.995 157.925 34.285 158.605 ;
        RECT 34.295 157.925 41.605 158.605 ;
        RECT 33.365 157.695 34.285 157.925 ;
        RECT 37.810 157.705 38.720 157.925 ;
        RECT 40.255 157.695 41.605 157.925 ;
        RECT 41.655 157.795 43.025 158.605 ;
        RECT 43.045 157.735 43.475 158.520 ;
        RECT 43.495 157.795 45.325 158.605 ;
        RECT 45.335 157.695 48.545 158.605 ;
        RECT 48.555 157.795 49.925 158.605 ;
        RECT 49.935 157.695 53.590 158.605 ;
        RECT 53.615 157.695 55.430 158.605 ;
        RECT 56.375 157.695 60.030 158.605 ;
        RECT 60.975 157.695 64.185 158.605 ;
        RECT 64.505 157.925 66.340 158.605 ;
        RECT 64.505 157.695 65.435 157.925 ;
        RECT 66.495 157.795 68.325 158.605 ;
        RECT 68.805 157.735 69.235 158.520 ;
        RECT 69.715 157.925 77.025 158.605 ;
        RECT 73.230 157.705 74.140 157.925 ;
        RECT 75.675 157.695 77.025 157.925 ;
        RECT 77.075 157.795 79.825 158.605 ;
        RECT 80.295 157.925 89.400 158.605 ;
        RECT 89.605 157.925 93.070 158.605 ;
        RECT 92.150 157.695 93.070 157.925 ;
        RECT 93.175 157.795 94.545 158.605 ;
        RECT 94.565 157.735 94.995 158.520 ;
        RECT 95.015 157.925 98.915 158.605 ;
        RECT 99.155 157.925 103.055 158.605 ;
        RECT 95.015 157.695 95.945 157.925 ;
        RECT 99.155 157.695 100.085 157.925 ;
        RECT 103.305 157.695 104.655 158.605 ;
        RECT 104.675 157.925 108.575 158.605 ;
        RECT 104.675 157.695 105.605 157.925 ;
        RECT 108.815 157.795 110.645 158.605 ;
        RECT 110.765 157.925 114.230 158.605 ;
        RECT 113.310 157.695 114.230 157.925 ;
        RECT 114.335 157.695 116.165 158.605 ;
        RECT 116.175 157.695 118.005 158.605 ;
        RECT 118.015 157.695 119.845 158.605 ;
        RECT 120.325 157.735 120.755 158.520 ;
        RECT 121.525 157.695 124.445 158.605 ;
        RECT 124.475 157.695 125.825 158.605 ;
        RECT 126.900 157.925 128.735 158.605 ;
        RECT 127.805 157.695 128.735 157.925 ;
        RECT 129.055 157.695 132.265 158.605 ;
        RECT 132.275 157.795 134.105 158.605 ;
        RECT 134.115 157.925 141.425 158.605 ;
        RECT 137.630 157.705 138.540 157.925 ;
        RECT 140.075 157.695 141.425 157.925 ;
        RECT 141.475 157.925 145.375 158.605 ;
        RECT 141.475 157.695 142.405 157.925 ;
        RECT 145.615 157.795 146.985 158.605 ;
      LAYER nwell ;
        RECT 17.080 154.575 147.180 157.405 ;
      LAYER pwell ;
        RECT 17.275 153.375 18.645 154.185 ;
        RECT 18.655 153.375 24.165 154.185 ;
        RECT 24.175 153.375 29.685 154.185 ;
        RECT 30.165 153.460 30.595 154.245 ;
        RECT 31.115 154.055 32.465 154.285 ;
        RECT 34.000 154.055 34.910 154.275 ;
        RECT 31.115 153.375 38.425 154.055 ;
        RECT 38.435 153.375 41.355 154.285 ;
        RECT 42.115 153.375 45.325 154.285 ;
        RECT 45.345 153.375 48.075 154.285 ;
        RECT 48.095 153.375 53.605 154.185 ;
        RECT 53.615 153.375 55.445 154.185 ;
        RECT 55.925 153.460 56.355 154.245 ;
        RECT 58.435 154.195 59.385 154.285 ;
        RECT 57.455 153.375 59.385 154.195 ;
        RECT 59.595 154.085 60.525 154.285 ;
        RECT 61.855 154.085 62.805 154.285 ;
        RECT 59.595 153.605 62.805 154.085 ;
        RECT 59.740 153.405 62.805 153.605 ;
        RECT 17.415 153.165 17.585 153.375 ;
        RECT 18.795 153.165 18.965 153.375 ;
        RECT 24.315 153.165 24.485 153.375 ;
        RECT 29.835 153.325 30.005 153.355 ;
        RECT 29.830 153.215 30.005 153.325 ;
        RECT 30.750 153.215 30.870 153.325 ;
        RECT 31.670 153.215 31.790 153.325 ;
        RECT 29.835 153.165 30.005 153.215 ;
        RECT 32.135 153.165 32.305 153.355 ;
        RECT 34.905 153.210 35.065 153.320 ;
        RECT 38.115 153.165 38.285 153.375 ;
        RECT 38.580 153.185 38.750 153.375 ;
        RECT 41.335 153.165 41.505 153.355 ;
        RECT 41.795 153.325 41.965 153.355 ;
        RECT 41.790 153.215 41.965 153.325 ;
        RECT 41.795 153.165 41.965 153.215 ;
        RECT 43.635 153.165 43.805 153.355 ;
        RECT 45.025 153.185 45.195 153.375 ;
        RECT 47.775 153.185 47.945 153.375 ;
        RECT 48.235 153.185 48.405 153.375 ;
        RECT 49.155 153.165 49.325 153.355 ;
        RECT 53.755 153.185 53.925 153.375 ;
        RECT 57.455 153.355 57.605 153.375 ;
        RECT 55.600 153.325 55.770 153.355 ;
        RECT 55.590 153.215 55.770 153.325 ;
        RECT 56.050 153.215 56.170 153.325 ;
        RECT 55.600 153.165 55.770 153.215 ;
        RECT 17.275 152.355 18.645 153.165 ;
        RECT 18.655 152.355 24.165 153.165 ;
        RECT 24.175 152.355 29.685 153.165 ;
        RECT 29.695 152.355 31.525 153.165 ;
        RECT 31.995 152.485 34.745 153.165 ;
        RECT 33.815 152.255 34.745 152.485 ;
        RECT 35.685 152.255 38.415 153.165 ;
        RECT 38.435 152.485 41.645 153.165 ;
        RECT 38.435 152.255 39.570 152.485 ;
        RECT 41.655 152.355 43.025 153.165 ;
        RECT 43.045 152.295 43.475 153.080 ;
        RECT 43.495 152.355 49.005 153.165 ;
        RECT 49.015 152.355 54.525 153.165 ;
        RECT 54.535 152.255 55.885 153.165 ;
        RECT 56.520 153.135 56.690 153.355 ;
        RECT 57.435 153.185 57.605 153.355 ;
        RECT 59.740 153.325 59.910 153.405 ;
        RECT 61.870 153.375 62.805 153.405 ;
        RECT 63.125 154.055 64.055 154.285 ;
        RECT 63.125 153.375 64.960 154.055 ;
        RECT 65.115 153.375 70.625 154.185 ;
        RECT 70.635 153.375 76.145 154.185 ;
        RECT 76.925 154.055 77.855 154.285 ;
        RECT 76.925 153.375 78.760 154.055 ;
        RECT 78.925 153.375 80.275 154.285 ;
        RECT 80.295 153.375 81.665 154.185 ;
        RECT 81.685 153.460 82.115 154.245 ;
        RECT 82.135 153.375 85.805 154.185 ;
        RECT 85.815 153.375 87.185 154.185 ;
        RECT 87.235 154.055 88.585 154.285 ;
        RECT 90.120 154.055 91.030 154.275 ;
        RECT 98.070 154.055 98.980 154.275 ;
        RECT 100.515 154.055 101.865 154.285 ;
        RECT 105.490 154.055 106.410 154.285 ;
        RECT 87.235 153.375 94.545 154.055 ;
        RECT 94.555 153.375 101.865 154.055 ;
        RECT 102.945 153.375 106.410 154.055 ;
        RECT 107.445 153.460 107.875 154.245 ;
        RECT 107.935 154.055 109.285 154.285 ;
        RECT 110.820 154.055 111.730 154.275 ;
        RECT 115.255 154.055 116.185 154.285 ;
        RECT 122.050 154.055 122.970 154.285 ;
        RECT 107.935 153.375 115.245 154.055 ;
        RECT 115.255 153.375 119.155 154.055 ;
        RECT 119.505 153.375 122.970 154.055 ;
        RECT 123.075 153.375 124.905 154.285 ;
        RECT 124.915 154.055 125.845 154.285 ;
        RECT 129.150 154.055 130.070 154.285 ;
        RECT 124.915 153.375 128.815 154.055 ;
        RECT 129.150 153.375 132.615 154.055 ;
        RECT 133.205 153.460 133.635 154.245 ;
        RECT 137.630 154.055 138.540 154.275 ;
        RECT 140.075 154.055 141.425 154.285 ;
        RECT 144.590 154.055 145.510 154.285 ;
        RECT 134.115 153.375 141.425 154.055 ;
        RECT 142.045 153.375 145.510 154.055 ;
        RECT 145.615 153.375 146.985 154.185 ;
        RECT 64.795 153.355 64.960 153.375 ;
        RECT 59.730 153.215 59.910 153.325 ;
        RECT 59.740 153.185 59.910 153.215 ;
        RECT 60.195 153.165 60.365 153.355 ;
        RECT 64.795 153.185 64.965 153.355 ;
        RECT 65.255 153.185 65.425 153.375 ;
        RECT 67.555 153.165 67.725 153.355 ;
        RECT 69.395 153.165 69.565 153.355 ;
        RECT 70.775 153.185 70.945 153.375 ;
        RECT 78.595 153.355 78.760 153.375 ;
        RECT 72.150 153.165 72.320 153.355 ;
        RECT 73.535 153.165 73.705 153.355 ;
        RECT 76.290 153.215 76.410 153.325 ;
        RECT 77.030 153.165 77.200 153.355 ;
        RECT 78.595 153.185 78.765 153.355 ;
        RECT 79.975 153.185 80.145 153.375 ;
        RECT 80.435 153.185 80.605 153.375 ;
        RECT 80.890 153.215 81.010 153.325 ;
        RECT 82.275 153.185 82.445 153.375 ;
        RECT 85.955 153.185 86.125 153.375 ;
        RECT 88.715 153.165 88.885 153.355 ;
        RECT 89.175 153.165 89.345 153.355 ;
        RECT 91.935 153.165 92.105 153.355 ;
        RECT 94.235 153.185 94.405 153.375 ;
        RECT 94.695 153.185 94.865 153.375 ;
        RECT 98.375 153.165 98.545 153.355 ;
        RECT 98.835 153.165 99.005 153.355 ;
        RECT 100.215 153.165 100.385 153.355 ;
        RECT 102.065 153.220 102.225 153.330 ;
        RECT 102.975 153.185 103.145 153.375 ;
        RECT 103.895 153.165 104.065 153.355 ;
        RECT 106.655 153.165 106.825 153.355 ;
        RECT 112.175 153.165 112.345 153.355 ;
        RECT 114.935 153.185 115.105 153.375 ;
        RECT 115.670 153.185 115.840 153.375 ;
        RECT 119.535 153.185 119.705 153.375 ;
        RECT 120.915 153.165 121.085 153.355 ;
        RECT 124.135 153.165 124.305 153.355 ;
        RECT 124.590 153.185 124.760 153.375 ;
        RECT 125.330 153.185 125.500 153.375 ;
        RECT 131.495 153.165 131.665 153.355 ;
        RECT 132.415 153.185 132.585 153.375 ;
        RECT 132.870 153.215 132.990 153.325 ;
        RECT 133.790 153.215 133.910 153.325 ;
        RECT 134.255 153.185 134.425 153.375 ;
        RECT 137.010 153.215 137.130 153.325 ;
        RECT 137.475 153.165 137.645 153.355 ;
        RECT 139.775 153.165 139.945 153.355 ;
        RECT 140.235 153.165 140.405 153.355 ;
        RECT 141.610 153.215 141.730 153.325 ;
        RECT 142.075 153.165 142.245 153.375 ;
        RECT 146.675 153.165 146.845 153.375 ;
        RECT 58.650 153.135 59.585 153.165 ;
        RECT 56.520 152.935 59.585 153.135 ;
        RECT 56.375 152.455 59.585 152.935 ;
        RECT 60.055 152.485 67.365 153.165 ;
        RECT 56.375 152.255 57.305 152.455 ;
        RECT 58.635 152.255 59.585 152.455 ;
        RECT 63.570 152.265 64.480 152.485 ;
        RECT 66.015 152.255 67.365 152.485 ;
        RECT 67.415 152.355 68.785 153.165 ;
        RECT 68.805 152.295 69.235 153.080 ;
        RECT 69.255 152.355 72.005 153.165 ;
        RECT 72.035 152.255 73.385 153.165 ;
        RECT 73.395 152.255 76.145 153.165 ;
        RECT 76.615 152.485 80.515 153.165 ;
        RECT 81.295 152.485 89.025 153.165 ;
        RECT 76.615 152.255 77.545 152.485 ;
        RECT 81.295 152.255 83.065 152.485 ;
        RECT 84.600 152.265 85.510 152.485 ;
        RECT 89.035 152.355 91.785 153.165 ;
        RECT 91.795 152.255 94.545 153.165 ;
        RECT 94.565 152.295 94.995 153.080 ;
        RECT 95.110 152.485 98.575 153.165 ;
        RECT 95.110 152.255 96.030 152.485 ;
        RECT 98.695 152.355 100.065 153.165 ;
        RECT 100.185 152.485 103.650 153.165 ;
        RECT 102.730 152.255 103.650 152.485 ;
        RECT 103.755 152.255 106.505 153.165 ;
        RECT 106.515 152.355 112.025 153.165 ;
        RECT 112.035 152.485 119.345 153.165 ;
        RECT 115.550 152.265 116.460 152.485 ;
        RECT 117.995 152.255 119.345 152.485 ;
        RECT 120.325 152.295 120.755 153.080 ;
        RECT 120.775 152.255 123.985 153.165 ;
        RECT 123.995 152.485 131.305 153.165 ;
        RECT 127.510 152.265 128.420 152.485 ;
        RECT 129.955 152.255 131.305 152.485 ;
        RECT 131.355 152.355 136.865 153.165 ;
        RECT 137.335 152.385 138.705 153.165 ;
        RECT 138.715 152.385 140.085 153.165 ;
        RECT 140.095 152.485 141.925 153.165 ;
        RECT 142.045 152.485 145.510 153.165 ;
        RECT 140.580 152.255 141.925 152.485 ;
        RECT 144.590 152.255 145.510 152.485 ;
        RECT 145.615 152.355 146.985 153.165 ;
      LAYER nwell ;
        RECT 17.080 149.135 147.180 151.965 ;
      LAYER pwell ;
        RECT 17.275 147.935 18.645 148.745 ;
        RECT 18.655 147.935 24.165 148.745 ;
        RECT 24.175 147.935 29.685 148.745 ;
        RECT 30.165 148.020 30.595 148.805 ;
        RECT 30.615 147.935 32.445 148.745 ;
        RECT 32.455 148.645 33.385 148.845 ;
        RECT 34.715 148.645 35.665 148.845 ;
        RECT 32.455 148.165 35.665 148.645 ;
        RECT 39.190 148.615 40.100 148.835 ;
        RECT 41.635 148.615 42.985 148.845 ;
        RECT 32.600 147.965 35.665 148.165 ;
        RECT 17.415 147.725 17.585 147.935 ;
        RECT 18.795 147.745 18.965 147.935 ;
        RECT 20.175 147.725 20.345 147.915 ;
        RECT 20.635 147.725 20.805 147.915 ;
        RECT 24.315 147.745 24.485 147.935 ;
        RECT 26.155 147.725 26.325 147.915 ;
        RECT 28.910 147.775 29.030 147.885 ;
        RECT 29.830 147.775 29.950 147.885 ;
        RECT 30.755 147.745 30.925 147.935 ;
        RECT 32.600 147.745 32.770 147.965 ;
        RECT 34.730 147.935 35.665 147.965 ;
        RECT 35.675 147.935 42.985 148.615 ;
        RECT 43.035 147.935 44.405 148.745 ;
        RECT 44.650 147.935 49.465 148.615 ;
        RECT 49.475 147.935 52.225 148.745 ;
        RECT 52.695 147.935 55.615 148.845 ;
        RECT 55.925 148.020 56.355 148.805 ;
        RECT 56.375 147.935 57.745 148.745 ;
        RECT 57.755 147.935 62.570 148.615 ;
        RECT 62.910 147.935 66.780 148.845 ;
        RECT 66.955 148.615 67.875 148.845 ;
        RECT 66.955 147.935 69.245 148.615 ;
        RECT 69.255 147.935 71.085 148.845 ;
        RECT 74.610 148.615 75.520 148.835 ;
        RECT 77.055 148.615 78.405 148.845 ;
        RECT 80.530 148.615 81.665 148.845 ;
        RECT 71.095 147.935 78.405 148.615 ;
        RECT 78.455 147.935 81.665 148.615 ;
        RECT 81.685 148.020 82.115 148.805 ;
        RECT 85.335 148.615 86.265 148.845 ;
        RECT 82.365 147.935 86.265 148.615 ;
        RECT 86.285 147.935 89.015 148.845 ;
        RECT 89.035 147.935 90.405 148.745 ;
        RECT 93.930 148.615 94.840 148.835 ;
        RECT 96.375 148.615 97.725 148.845 ;
        RECT 101.455 148.615 102.385 148.845 ;
        RECT 106.035 148.615 106.965 148.845 ;
        RECT 90.415 147.935 97.725 148.615 ;
        RECT 97.775 147.935 100.515 148.615 ;
        RECT 101.455 147.935 104.205 148.615 ;
        RECT 104.215 147.935 106.965 148.615 ;
        RECT 107.445 148.020 107.875 148.805 ;
        RECT 107.895 147.935 113.405 148.745 ;
        RECT 113.415 147.935 118.925 148.745 ;
        RECT 118.935 147.935 120.305 148.745 ;
        RECT 120.315 147.935 123.525 148.845 ;
        RECT 123.555 147.935 124.905 148.845 ;
        RECT 124.915 147.935 128.585 148.745 ;
        RECT 128.595 147.935 129.965 148.745 ;
        RECT 129.975 147.935 133.185 148.845 ;
        RECT 133.205 148.020 133.635 148.805 ;
        RECT 134.575 148.615 135.505 148.845 ;
        RECT 138.810 148.615 139.730 148.845 ;
        RECT 134.575 147.935 138.475 148.615 ;
        RECT 138.810 147.935 142.275 148.615 ;
        RECT 142.395 147.935 143.765 148.715 ;
        RECT 144.260 148.615 145.605 148.845 ;
        RECT 143.775 147.935 145.605 148.615 ;
        RECT 145.615 147.935 146.985 148.745 ;
        RECT 35.815 147.745 35.985 147.935 ;
        RECT 36.275 147.725 36.445 147.915 ;
        RECT 36.735 147.725 36.905 147.915 ;
        RECT 39.955 147.745 40.125 147.915 ;
        RECT 39.955 147.725 40.120 147.745 ;
        RECT 40.415 147.725 40.585 147.915 ;
        RECT 43.175 147.745 43.345 147.935 ;
        RECT 43.645 147.770 43.805 147.880 ;
        RECT 44.555 147.745 44.725 147.915 ;
        RECT 48.690 147.775 48.810 147.885 ;
        RECT 49.155 147.745 49.325 147.935 ;
        RECT 49.615 147.745 49.785 147.935 ;
        RECT 44.580 147.725 44.725 147.745 ;
        RECT 49.175 147.725 49.325 147.745 ;
        RECT 17.275 146.915 18.645 147.725 ;
        RECT 18.655 147.045 20.485 147.725 ;
        RECT 18.655 146.815 20.000 147.045 ;
        RECT 20.495 146.915 26.005 147.725 ;
        RECT 26.015 146.915 28.765 147.725 ;
        RECT 29.275 147.045 36.585 147.725 ;
        RECT 29.275 146.815 30.625 147.045 ;
        RECT 32.160 146.825 33.070 147.045 ;
        RECT 36.595 146.915 37.965 147.725 ;
        RECT 38.285 147.045 40.120 147.725 ;
        RECT 38.285 146.815 39.215 147.045 ;
        RECT 40.285 146.815 43.015 147.725 ;
        RECT 43.045 146.855 43.475 147.640 ;
        RECT 44.580 146.815 48.450 147.725 ;
        RECT 49.175 146.905 51.105 147.725 ;
        RECT 51.460 147.695 51.630 147.915 ;
        RECT 52.370 147.775 52.490 147.885 ;
        RECT 52.840 147.745 53.010 147.935 ;
        RECT 54.685 147.770 54.845 147.880 ;
        RECT 56.515 147.745 56.685 147.935 ;
        RECT 57.895 147.745 58.065 147.935 ;
        RECT 66.635 147.915 66.780 147.935 ;
        RECT 62.495 147.725 62.665 147.915 ;
        RECT 64.795 147.745 64.965 147.915 ;
        RECT 64.795 147.725 64.960 147.745 ;
        RECT 65.255 147.725 65.425 147.915 ;
        RECT 66.635 147.745 66.805 147.915 ;
        RECT 68.935 147.745 69.105 147.935 ;
        RECT 69.400 147.745 69.570 147.935 ;
        RECT 70.315 147.725 70.485 147.915 ;
        RECT 71.235 147.745 71.405 147.935 ;
        RECT 77.685 147.770 77.845 147.880 ;
        RECT 78.595 147.725 78.765 147.935 ;
        RECT 82.275 147.725 82.445 147.915 ;
        RECT 85.680 147.745 85.850 147.935 ;
        RECT 53.590 147.695 54.525 147.725 ;
        RECT 51.460 147.495 54.525 147.695 ;
        RECT 50.155 146.815 51.105 146.905 ;
        RECT 51.315 147.015 54.525 147.495 ;
        RECT 51.315 146.815 52.245 147.015 ;
        RECT 53.575 146.815 54.525 147.015 ;
        RECT 55.495 147.045 62.805 147.725 ;
        RECT 63.125 147.045 64.960 147.725 ;
        RECT 55.495 146.815 56.845 147.045 ;
        RECT 58.380 146.825 59.290 147.045 ;
        RECT 63.125 146.815 64.055 147.045 ;
        RECT 65.115 146.915 68.785 147.725 ;
        RECT 68.805 146.855 69.235 147.640 ;
        RECT 70.175 147.045 77.485 147.725 ;
        RECT 78.565 147.045 82.030 147.725 ;
        RECT 82.245 147.045 85.710 147.725 ;
        RECT 85.955 147.695 86.125 147.915 ;
        RECT 88.715 147.725 88.885 147.935 ;
        RECT 89.175 147.745 89.345 147.935 ;
        RECT 90.555 147.745 90.725 147.935 ;
        RECT 94.230 147.775 94.350 147.885 ;
        RECT 95.155 147.725 95.325 147.915 ;
        RECT 97.915 147.745 98.085 147.935 ;
        RECT 100.685 147.725 100.855 147.915 ;
        RECT 101.145 147.770 101.305 147.880 ;
        RECT 102.055 147.725 102.225 147.915 ;
        RECT 103.895 147.745 104.065 147.935 ;
        RECT 104.355 147.745 104.525 147.935 ;
        RECT 107.110 147.775 107.230 147.885 ;
        RECT 108.035 147.745 108.205 147.935 ;
        RECT 109.415 147.725 109.585 147.915 ;
        RECT 113.555 147.745 113.725 147.935 ;
        RECT 116.775 147.725 116.945 147.915 ;
        RECT 119.075 147.745 119.245 147.935 ;
        RECT 120.455 147.745 120.625 147.935 ;
        RECT 123.670 147.745 123.840 147.935 ;
        RECT 124.135 147.725 124.305 147.915 ;
        RECT 124.595 147.725 124.765 147.915 ;
        RECT 125.055 147.745 125.225 147.935 ;
        RECT 128.275 147.725 128.445 147.915 ;
        RECT 128.735 147.745 128.905 147.935 ;
        RECT 129.655 147.725 129.825 147.915 ;
        RECT 130.115 147.745 130.285 147.935 ;
        RECT 132.870 147.775 132.990 147.885 ;
        RECT 133.335 147.725 133.505 147.915 ;
        RECT 133.805 147.780 133.965 147.890 ;
        RECT 134.990 147.745 135.160 147.935 ;
        RECT 140.695 147.725 140.865 147.915 ;
        RECT 142.075 147.725 142.245 147.935 ;
        RECT 143.455 147.745 143.625 147.935 ;
        RECT 143.915 147.725 144.085 147.935 ;
        RECT 146.675 147.725 146.845 147.935 ;
        RECT 87.155 147.695 88.535 147.725 ;
        RECT 73.690 146.825 74.600 147.045 ;
        RECT 76.135 146.815 77.485 147.045 ;
        RECT 81.110 146.815 82.030 147.045 ;
        RECT 84.790 146.815 85.710 147.045 ;
        RECT 85.830 147.015 88.535 147.695 ;
        RECT 87.155 146.815 88.535 147.015 ;
        RECT 88.575 146.915 94.085 147.725 ;
        RECT 94.565 146.855 94.995 147.640 ;
        RECT 95.015 146.915 97.765 147.725 ;
        RECT 97.775 146.815 100.985 147.725 ;
        RECT 101.915 147.045 109.225 147.725 ;
        RECT 109.275 147.045 116.585 147.725 ;
        RECT 105.430 146.825 106.340 147.045 ;
        RECT 107.875 146.815 109.225 147.045 ;
        RECT 112.790 146.825 113.700 147.045 ;
        RECT 115.235 146.815 116.585 147.045 ;
        RECT 116.635 146.915 120.305 147.725 ;
        RECT 120.325 146.855 120.755 147.640 ;
        RECT 120.870 147.045 124.335 147.725 ;
        RECT 120.870 146.815 121.790 147.045 ;
        RECT 124.455 146.915 128.125 147.725 ;
        RECT 128.135 146.915 129.505 147.725 ;
        RECT 129.515 146.815 132.725 147.725 ;
        RECT 133.195 147.045 140.505 147.725 ;
        RECT 136.710 146.825 137.620 147.045 ;
        RECT 139.155 146.815 140.505 147.045 ;
        RECT 140.555 146.945 141.925 147.725 ;
        RECT 141.935 147.045 143.765 147.725 ;
        RECT 143.775 147.045 145.605 147.725 ;
        RECT 142.420 146.815 143.765 147.045 ;
        RECT 144.260 146.815 145.605 147.045 ;
        RECT 145.615 146.915 146.985 147.725 ;
      LAYER nwell ;
        RECT 17.080 143.695 147.180 146.525 ;
      LAYER pwell ;
        RECT 17.275 142.495 18.645 143.305 ;
        RECT 18.655 143.175 20.000 143.405 ;
        RECT 18.655 142.495 20.485 143.175 ;
        RECT 20.495 142.495 26.005 143.305 ;
        RECT 26.015 142.495 29.685 143.305 ;
        RECT 30.165 142.580 30.595 143.365 ;
        RECT 30.615 142.495 34.285 143.305 ;
        RECT 36.585 143.175 37.505 143.405 ;
        RECT 35.215 142.495 37.505 143.175 ;
        RECT 37.515 143.205 38.445 143.405 ;
        RECT 39.775 143.205 40.725 143.405 ;
        RECT 37.515 142.725 40.725 143.205 ;
        RECT 44.250 143.175 45.160 143.395 ;
        RECT 46.695 143.175 48.045 143.405 ;
        RECT 49.465 143.175 50.385 143.405 ;
        RECT 52.365 143.175 53.295 143.405 ;
        RECT 54.985 143.175 55.905 143.405 ;
        RECT 37.660 142.525 40.725 142.725 ;
        RECT 17.415 142.285 17.585 142.495 ;
        RECT 18.790 142.335 18.910 142.445 ;
        RECT 19.255 142.285 19.425 142.475 ;
        RECT 20.175 142.305 20.345 142.495 ;
        RECT 20.635 142.305 20.805 142.495 ;
        RECT 26.155 142.305 26.325 142.495 ;
        RECT 26.625 142.330 26.785 142.440 ;
        RECT 27.535 142.305 27.705 142.475 ;
        RECT 29.835 142.445 30.005 142.475 ;
        RECT 29.830 142.335 30.005 142.445 ;
        RECT 27.540 142.285 27.705 142.305 ;
        RECT 29.835 142.285 30.005 142.335 ;
        RECT 30.755 142.305 30.925 142.495 ;
        RECT 34.445 142.340 34.605 142.450 ;
        RECT 35.355 142.445 35.525 142.495 ;
        RECT 35.350 142.335 35.525 142.445 ;
        RECT 35.355 142.305 35.525 142.335 ;
        RECT 35.815 142.285 35.985 142.475 ;
        RECT 37.660 142.305 37.830 142.525 ;
        RECT 39.790 142.495 40.725 142.525 ;
        RECT 40.735 142.495 48.045 143.175 ;
        RECT 48.095 142.495 50.385 143.175 ;
        RECT 51.460 142.495 53.295 143.175 ;
        RECT 53.615 142.495 55.905 143.175 ;
        RECT 55.925 142.580 56.355 143.365 ;
        RECT 59.890 143.175 60.800 143.395 ;
        RECT 62.335 143.175 63.685 143.405 ;
        RECT 56.375 142.495 63.685 143.175 ;
        RECT 63.735 142.495 69.245 143.305 ;
        RECT 69.255 142.495 72.005 143.305 ;
        RECT 75.530 143.175 76.440 143.395 ;
        RECT 77.975 143.175 79.325 143.405 ;
        RECT 72.015 142.495 79.325 143.175 ;
        RECT 79.375 142.495 81.205 143.405 ;
        RECT 81.685 142.580 82.115 143.365 ;
        RECT 82.230 143.175 83.150 143.405 ;
        RECT 82.230 142.495 85.695 143.175 ;
        RECT 85.835 142.495 87.185 143.405 ;
        RECT 91.630 143.175 92.540 143.395 ;
        RECT 94.075 143.175 95.425 143.405 ;
        RECT 88.115 142.495 95.425 143.175 ;
        RECT 95.475 142.495 96.845 143.305 ;
        RECT 96.855 142.495 100.065 143.405 ;
        RECT 100.075 142.495 102.825 143.305 ;
        RECT 103.295 143.175 104.225 143.405 ;
        RECT 103.295 142.495 107.195 143.175 ;
        RECT 107.445 142.580 107.875 143.365 ;
        RECT 107.895 143.175 108.825 143.405 ;
        RECT 107.895 142.495 111.795 143.175 ;
        RECT 112.035 142.495 117.545 143.305 ;
        RECT 118.515 143.175 119.865 143.405 ;
        RECT 121.400 143.175 122.310 143.395 ;
        RECT 128.490 143.175 129.410 143.405 ;
        RECT 118.515 142.495 125.825 143.175 ;
        RECT 125.945 142.495 129.410 143.175 ;
        RECT 129.515 142.495 133.185 143.305 ;
        RECT 133.205 142.580 133.635 143.365 ;
        RECT 137.170 143.175 138.080 143.395 ;
        RECT 139.615 143.175 140.965 143.405 ;
        RECT 133.655 142.495 140.965 143.175 ;
        RECT 141.110 143.175 142.030 143.405 ;
        RECT 141.110 142.495 144.575 143.175 ;
        RECT 145.615 142.495 146.985 143.305 ;
        RECT 40.875 142.305 41.045 142.495 ;
        RECT 44.560 142.285 44.730 142.475 ;
        RECT 45.015 142.285 45.185 142.475 ;
        RECT 48.235 142.305 48.405 142.495 ;
        RECT 51.460 142.475 51.625 142.495 ;
        RECT 50.545 142.330 50.705 142.450 ;
        RECT 51.455 142.305 51.625 142.475 ;
        RECT 53.755 142.305 53.925 142.495 ;
        RECT 56.515 142.305 56.685 142.495 ;
        RECT 58.355 142.285 58.525 142.475 ;
        RECT 58.815 142.285 58.985 142.475 ;
        RECT 63.875 142.305 64.045 142.495 ;
        RECT 64.335 142.285 64.505 142.475 ;
        RECT 65.715 142.285 65.885 142.475 ;
        RECT 69.395 142.285 69.565 142.495 ;
        RECT 72.155 142.305 72.325 142.495 ;
        RECT 74.455 142.285 74.625 142.475 ;
        RECT 77.220 142.285 77.390 142.475 ;
        RECT 79.055 142.285 79.225 142.475 ;
        RECT 79.520 142.305 79.690 142.495 ;
        RECT 81.350 142.335 81.470 142.445 ;
        RECT 84.570 142.335 84.690 142.445 ;
        RECT 85.035 142.285 85.205 142.475 ;
        RECT 85.495 142.305 85.665 142.495 ;
        RECT 85.950 142.305 86.120 142.495 ;
        RECT 86.415 142.285 86.585 142.475 ;
        RECT 87.345 142.340 87.505 142.450 ;
        RECT 88.255 142.305 88.425 142.495 ;
        RECT 88.710 142.335 88.830 142.445 ;
        RECT 89.450 142.285 89.620 142.475 ;
        RECT 93.315 142.285 93.485 142.475 ;
        RECT 95.155 142.285 95.325 142.475 ;
        RECT 95.615 142.305 95.785 142.495 ;
        RECT 96.985 142.305 97.155 142.495 ;
        RECT 100.215 142.305 100.385 142.495 ;
        RECT 100.675 142.285 100.845 142.475 ;
        RECT 102.515 142.285 102.685 142.475 ;
        RECT 102.970 142.335 103.090 142.445 ;
        RECT 103.710 142.305 103.880 142.495 ;
        RECT 106.195 142.285 106.365 142.475 ;
        RECT 108.035 142.285 108.205 142.475 ;
        RECT 108.310 142.305 108.480 142.495 ;
        RECT 112.175 142.305 112.345 142.495 ;
        RECT 113.095 142.285 113.265 142.475 ;
        RECT 113.555 142.285 113.725 142.475 ;
        RECT 117.230 142.335 117.350 142.445 ;
        RECT 117.705 142.340 117.865 142.450 ;
        RECT 119.995 142.285 120.165 142.475 ;
        RECT 125.515 142.305 125.685 142.495 ;
        RECT 125.975 142.305 126.145 142.495 ;
        RECT 127.815 142.285 127.985 142.475 ;
        RECT 128.275 142.285 128.445 142.475 ;
        RECT 129.655 142.305 129.825 142.495 ;
        RECT 131.035 142.285 131.205 142.475 ;
        RECT 133.795 142.305 133.965 142.495 ;
        RECT 134.070 142.285 134.240 142.475 ;
        RECT 138.210 142.285 138.380 142.475 ;
        RECT 142.075 142.285 142.245 142.475 ;
        RECT 143.450 142.335 143.570 142.445 ;
        RECT 143.915 142.285 144.085 142.475 ;
        RECT 144.375 142.305 144.545 142.495 ;
        RECT 144.845 142.340 145.005 142.450 ;
        RECT 146.675 142.285 146.845 142.495 ;
        RECT 17.275 141.475 18.645 142.285 ;
        RECT 19.115 141.605 26.425 142.285 ;
        RECT 27.540 141.605 29.375 142.285 ;
        RECT 22.630 141.385 23.540 141.605 ;
        RECT 25.075 141.375 26.425 141.605 ;
        RECT 28.445 141.375 29.375 141.605 ;
        RECT 29.695 141.475 35.205 142.285 ;
        RECT 35.675 141.605 42.985 142.285 ;
        RECT 39.190 141.385 40.100 141.605 ;
        RECT 41.635 141.375 42.985 141.605 ;
        RECT 43.045 141.415 43.475 142.200 ;
        RECT 43.495 141.375 44.845 142.285 ;
        RECT 44.875 141.475 50.385 142.285 ;
        RECT 51.355 141.605 58.665 142.285 ;
        RECT 51.355 141.375 52.705 141.605 ;
        RECT 54.240 141.385 55.150 141.605 ;
        RECT 58.675 141.475 64.185 142.285 ;
        RECT 64.195 141.475 65.565 142.285 ;
        RECT 65.625 141.375 68.785 142.285 ;
        RECT 68.805 141.415 69.235 142.200 ;
        RECT 69.255 141.605 74.070 142.285 ;
        RECT 74.315 141.475 77.065 142.285 ;
        RECT 77.075 141.375 78.905 142.285 ;
        RECT 78.915 141.475 84.425 142.285 ;
        RECT 84.905 141.375 86.255 142.285 ;
        RECT 86.275 141.605 88.565 142.285 ;
        RECT 87.645 141.375 88.565 141.605 ;
        RECT 89.035 141.605 92.935 142.285 ;
        RECT 89.035 141.375 89.965 141.605 ;
        RECT 93.175 141.475 94.545 142.285 ;
        RECT 94.565 141.415 94.995 142.200 ;
        RECT 95.015 141.475 100.525 142.285 ;
        RECT 100.535 141.475 102.365 142.285 ;
        RECT 102.485 141.605 105.950 142.285 ;
        RECT 105.030 141.375 105.950 141.605 ;
        RECT 106.055 141.475 107.885 142.285 ;
        RECT 107.895 141.375 110.645 142.285 ;
        RECT 110.665 141.605 113.405 142.285 ;
        RECT 113.415 141.475 117.085 142.285 ;
        RECT 117.555 141.375 120.305 142.285 ;
        RECT 120.325 141.415 120.755 142.200 ;
        RECT 120.815 141.605 128.125 142.285 ;
        RECT 120.815 141.375 122.165 141.605 ;
        RECT 123.700 141.385 124.610 141.605 ;
        RECT 128.135 141.375 130.885 142.285 ;
        RECT 130.895 141.475 133.645 142.285 ;
        RECT 133.655 141.605 137.555 142.285 ;
        RECT 137.795 141.605 141.695 142.285 ;
        RECT 133.655 141.375 134.585 141.605 ;
        RECT 137.795 141.375 138.725 141.605 ;
        RECT 141.935 141.505 143.305 142.285 ;
        RECT 143.775 141.605 145.605 142.285 ;
        RECT 144.260 141.375 145.605 141.605 ;
        RECT 145.615 141.475 146.985 142.285 ;
      LAYER nwell ;
        RECT 17.080 138.255 147.180 141.085 ;
      LAYER pwell ;
        RECT 17.275 137.055 18.645 137.865 ;
        RECT 18.655 137.735 19.585 137.965 ;
        RECT 22.835 137.735 24.185 137.965 ;
        RECT 25.720 137.735 26.630 137.955 ;
        RECT 18.655 137.055 22.555 137.735 ;
        RECT 22.835 137.055 30.145 137.735 ;
        RECT 30.165 137.140 30.595 137.925 ;
        RECT 30.695 137.055 33.695 137.965 ;
        RECT 33.835 137.055 39.345 137.865 ;
        RECT 39.355 137.055 44.865 137.865 ;
        RECT 44.875 137.055 50.385 137.865 ;
        RECT 50.395 137.055 55.905 137.865 ;
        RECT 55.925 137.140 56.355 137.925 ;
        RECT 56.375 137.055 61.885 137.865 ;
        RECT 61.895 137.055 67.405 137.865 ;
        RECT 67.415 137.055 68.785 137.865 ;
        RECT 68.835 137.055 72.005 137.965 ;
        RECT 72.015 137.765 72.965 137.965 ;
        RECT 74.295 137.765 75.225 137.965 ;
        RECT 72.015 137.285 75.225 137.765 ;
        RECT 72.015 137.085 75.080 137.285 ;
        RECT 72.015 137.055 72.950 137.085 ;
        RECT 17.415 136.845 17.585 137.055 ;
        RECT 19.070 136.865 19.240 137.055 ;
        RECT 20.175 136.845 20.345 137.035 ;
        RECT 20.645 136.845 20.815 137.035 ;
        RECT 22.015 136.845 22.185 137.035 ;
        RECT 24.775 136.845 24.945 137.035 ;
        RECT 29.835 136.865 30.005 137.055 ;
        RECT 30.755 136.865 30.925 137.055 ;
        RECT 32.135 136.845 32.305 137.035 ;
        RECT 33.515 136.845 33.685 137.035 ;
        RECT 33.975 136.865 34.145 137.055 ;
        RECT 39.035 136.845 39.205 137.035 ;
        RECT 39.495 136.865 39.665 137.055 ;
        RECT 42.710 136.895 42.830 137.005 ;
        RECT 43.635 136.845 43.805 137.035 ;
        RECT 45.015 136.865 45.185 137.055 ;
        RECT 49.155 136.845 49.325 137.035 ;
        RECT 50.535 136.865 50.705 137.055 ;
        RECT 54.675 136.845 54.845 137.035 ;
        RECT 56.515 136.865 56.685 137.055 ;
        RECT 60.195 136.845 60.365 137.035 ;
        RECT 62.035 136.865 62.205 137.055 ;
        RECT 63.875 136.845 64.045 137.035 ;
        RECT 66.170 136.845 66.340 137.035 ;
        RECT 67.555 136.865 67.725 137.055 ;
        RECT 68.475 136.865 68.645 137.035 ;
        RECT 68.935 136.865 69.105 137.055 ;
        RECT 68.475 136.845 68.640 136.865 ;
        RECT 69.395 136.845 69.565 137.035 ;
        RECT 74.910 136.865 75.080 137.085 ;
        RECT 75.235 137.055 80.745 137.865 ;
        RECT 81.685 137.140 82.115 137.925 ;
        RECT 83.930 137.765 84.885 137.965 ;
        RECT 82.605 137.085 84.885 137.765 ;
        RECT 84.895 137.765 85.825 137.965 ;
        RECT 87.160 137.765 88.105 137.965 ;
        RECT 84.895 137.285 88.105 137.765 ;
        RECT 75.375 136.865 75.545 137.055 ;
        RECT 82.730 137.035 82.900 137.085 ;
        RECT 83.930 137.055 84.885 137.085 ;
        RECT 85.035 137.085 88.105 137.285 ;
        RECT 77.680 136.845 77.850 137.035 ;
        RECT 78.135 136.845 78.305 137.035 ;
        RECT 17.275 136.035 18.645 136.845 ;
        RECT 18.655 136.165 20.485 136.845 ;
        RECT 18.655 135.935 20.000 136.165 ;
        RECT 20.495 136.065 21.865 136.845 ;
        RECT 21.875 136.035 24.625 136.845 ;
        RECT 24.635 136.165 31.945 136.845 ;
        RECT 28.150 135.945 29.060 136.165 ;
        RECT 30.595 135.935 31.945 136.165 ;
        RECT 32.005 135.935 33.355 136.845 ;
        RECT 33.375 136.035 38.885 136.845 ;
        RECT 38.895 136.035 42.565 136.845 ;
        RECT 43.045 135.975 43.475 136.760 ;
        RECT 43.495 136.035 49.005 136.845 ;
        RECT 49.015 136.035 54.525 136.845 ;
        RECT 54.535 136.035 60.045 136.845 ;
        RECT 60.055 136.035 63.725 136.845 ;
        RECT 63.735 136.035 65.105 136.845 ;
        RECT 65.135 135.935 66.485 136.845 ;
        RECT 66.805 136.165 68.640 136.845 ;
        RECT 66.805 135.935 67.735 136.165 ;
        RECT 68.805 135.975 69.235 136.760 ;
        RECT 69.255 136.165 76.565 136.845 ;
        RECT 72.770 135.945 73.680 136.165 ;
        RECT 75.215 135.935 76.565 136.165 ;
        RECT 76.615 135.935 77.965 136.845 ;
        RECT 77.995 136.035 79.365 136.845 ;
        RECT 79.515 136.815 79.685 137.035 ;
        RECT 80.905 136.900 81.065 137.010 ;
        RECT 82.270 136.895 82.390 137.005 ;
        RECT 82.730 136.865 82.905 137.035 ;
        RECT 85.035 136.865 85.205 137.085 ;
        RECT 87.160 137.055 88.105 137.085 ;
        RECT 88.115 137.735 89.045 137.965 ;
        RECT 92.255 137.735 93.185 137.965 ;
        RECT 88.115 137.055 92.015 137.735 ;
        RECT 92.255 137.055 96.155 137.735 ;
        RECT 96.395 137.055 100.065 137.865 ;
        RECT 100.535 137.055 104.405 137.965 ;
        RECT 104.675 137.055 107.425 137.965 ;
        RECT 107.445 137.140 107.875 137.925 ;
        RECT 107.895 137.055 109.725 137.865 ;
        RECT 110.290 137.735 111.210 137.965 ;
        RECT 117.390 137.735 118.300 137.955 ;
        RECT 119.835 137.735 121.185 137.965 ;
        RECT 124.750 137.735 125.660 137.955 ;
        RECT 127.195 137.735 128.545 137.965 ;
        RECT 110.290 137.055 113.755 137.735 ;
        RECT 113.875 137.055 121.185 137.735 ;
        RECT 121.235 137.055 128.545 137.735 ;
        RECT 128.595 137.055 130.425 137.865 ;
        RECT 132.255 137.735 133.185 137.965 ;
        RECT 130.435 137.055 133.185 137.735 ;
        RECT 133.205 137.140 133.635 137.925 ;
        RECT 133.655 137.055 136.865 137.965 ;
        RECT 140.850 137.735 141.760 137.955 ;
        RECT 143.295 137.735 144.645 137.965 ;
        RECT 137.335 137.055 144.645 137.735 ;
        RECT 145.615 137.055 146.985 137.865 ;
        RECT 85.965 136.890 86.125 137.000 ;
        RECT 81.640 136.815 82.585 136.845 ;
        RECT 79.515 136.615 82.585 136.815 ;
        RECT 82.735 136.815 82.905 136.865 ;
        RECT 86.875 136.845 87.045 137.035 ;
        RECT 88.530 136.865 88.700 137.055 ;
        RECT 92.670 136.865 92.840 137.055 ;
        RECT 95.155 136.845 95.325 137.035 ;
        RECT 96.535 136.865 96.705 137.055 ;
        RECT 98.845 136.890 99.005 137.000 ;
        RECT 100.210 136.895 100.330 137.005 ;
        RECT 100.680 136.865 100.850 137.055 ;
        RECT 104.815 136.865 104.985 137.055 ;
        RECT 106.655 136.845 106.825 137.035 ;
        RECT 107.115 136.845 107.285 137.035 ;
        RECT 108.035 136.865 108.205 137.055 ;
        RECT 109.870 136.895 109.990 137.005 ;
        RECT 113.555 136.865 113.725 137.055 ;
        RECT 114.015 136.865 114.185 137.055 ;
        RECT 114.475 136.845 114.645 137.035 ;
        RECT 116.310 136.895 116.430 137.005 ;
        RECT 116.775 136.845 116.945 137.035 ;
        RECT 119.545 136.890 119.705 137.000 ;
        RECT 121.375 136.865 121.545 137.055 ;
        RECT 128.735 137.035 128.905 137.055 ;
        RECT 124.135 136.845 124.305 137.035 ;
        RECT 127.815 136.845 127.985 137.035 ;
        RECT 128.270 136.895 128.390 137.005 ;
        RECT 128.725 136.865 128.905 137.035 ;
        RECT 130.575 136.865 130.745 137.055 ;
        RECT 133.785 136.865 133.955 137.055 ;
        RECT 128.725 136.845 128.895 136.865 ;
        RECT 135.360 136.845 135.530 137.035 ;
        RECT 136.095 136.845 136.265 137.035 ;
        RECT 137.010 136.895 137.130 137.005 ;
        RECT 137.475 136.865 137.645 137.055 ;
        RECT 143.450 136.895 143.570 137.005 ;
        RECT 143.915 136.845 144.085 137.035 ;
        RECT 144.845 136.900 145.005 137.010 ;
        RECT 146.675 136.845 146.845 137.055 ;
        RECT 84.860 136.815 85.805 136.845 ;
        RECT 82.735 136.615 85.805 136.815 ;
        RECT 79.375 136.135 82.585 136.615 ;
        RECT 79.375 135.935 80.305 136.135 ;
        RECT 81.640 135.935 82.585 136.135 ;
        RECT 82.595 136.135 85.805 136.615 ;
        RECT 86.735 136.165 94.465 136.845 ;
        RECT 82.595 135.935 83.525 136.135 ;
        RECT 84.860 135.935 85.805 136.135 ;
        RECT 90.250 135.945 91.160 136.165 ;
        RECT 92.695 135.935 94.465 136.165 ;
        RECT 94.565 135.975 94.995 136.760 ;
        RECT 95.015 136.035 98.685 136.845 ;
        RECT 99.655 136.165 106.965 136.845 ;
        RECT 106.975 136.165 114.285 136.845 ;
        RECT 99.655 135.935 101.005 136.165 ;
        RECT 102.540 135.945 103.450 136.165 ;
        RECT 110.490 135.945 111.400 136.165 ;
        RECT 112.935 135.935 114.285 136.165 ;
        RECT 114.335 136.035 116.165 136.845 ;
        RECT 116.635 135.935 119.385 136.845 ;
        RECT 120.325 135.975 120.755 136.760 ;
        RECT 120.870 136.165 124.335 136.845 ;
        RECT 124.550 136.165 128.015 136.845 ;
        RECT 120.870 135.935 121.790 136.165 ;
        RECT 124.550 135.935 125.470 136.165 ;
        RECT 128.595 135.935 131.805 136.845 ;
        RECT 132.045 136.165 135.945 136.845 ;
        RECT 135.955 136.165 143.265 136.845 ;
        RECT 143.775 136.165 145.605 136.845 ;
        RECT 135.015 135.935 135.945 136.165 ;
        RECT 139.470 135.945 140.380 136.165 ;
        RECT 141.915 135.935 143.265 136.165 ;
        RECT 144.260 135.935 145.605 136.165 ;
        RECT 145.615 136.035 146.985 136.845 ;
      LAYER nwell ;
        RECT 17.080 132.815 147.180 135.645 ;
      LAYER pwell ;
        RECT 17.275 131.615 18.645 132.425 ;
        RECT 22.630 132.295 23.540 132.515 ;
        RECT 25.075 132.295 26.425 132.525 ;
        RECT 19.115 131.615 26.425 132.295 ;
        RECT 27.015 131.615 30.015 132.525 ;
        RECT 30.165 131.700 30.595 132.485 ;
        RECT 30.925 132.295 31.855 132.525 ;
        RECT 30.925 131.615 32.760 132.295 ;
        RECT 32.925 131.615 34.275 132.525 ;
        RECT 34.295 131.615 39.805 132.425 ;
        RECT 39.815 131.615 45.325 132.425 ;
        RECT 45.335 131.615 50.845 132.425 ;
        RECT 50.855 131.615 54.525 132.425 ;
        RECT 54.535 131.615 55.905 132.425 ;
        RECT 55.925 131.700 56.355 132.485 ;
        RECT 56.375 131.615 61.885 132.425 ;
        RECT 65.410 132.295 66.320 132.515 ;
        RECT 67.855 132.295 69.625 132.525 ;
        RECT 61.895 131.615 69.625 132.295 ;
        RECT 69.915 132.435 70.865 132.525 ;
        RECT 69.915 131.615 71.845 132.435 ;
        RECT 75.990 132.295 76.900 132.515 ;
        RECT 78.435 132.295 79.785 132.525 ;
        RECT 72.475 131.615 79.785 132.295 ;
        RECT 79.835 131.615 81.665 132.425 ;
        RECT 81.685 131.700 82.115 132.485 ;
        RECT 82.135 131.615 83.505 132.425 ;
        RECT 86.715 132.295 87.645 132.525 ;
        RECT 91.170 132.295 92.080 132.515 ;
        RECT 93.615 132.295 95.385 132.525 ;
        RECT 83.745 131.615 87.645 132.295 ;
        RECT 87.655 131.615 95.385 132.295 ;
        RECT 95.570 132.295 96.490 132.525 ;
        RECT 102.270 132.295 103.190 132.525 ;
        RECT 106.495 132.295 107.425 132.525 ;
        RECT 95.570 131.615 99.035 132.295 ;
        RECT 99.725 131.615 103.190 132.295 ;
        RECT 103.525 131.615 107.425 132.295 ;
        RECT 107.445 131.700 107.875 132.485 ;
        RECT 111.410 132.295 112.320 132.515 ;
        RECT 113.855 132.295 115.205 132.525 ;
        RECT 107.895 131.615 115.205 132.295 ;
        RECT 115.255 131.615 120.765 132.425 ;
        RECT 120.775 131.615 123.525 132.525 ;
        RECT 123.535 131.615 129.045 132.425 ;
        RECT 129.055 131.615 132.725 132.425 ;
        RECT 133.205 131.700 133.635 132.485 ;
        RECT 135.475 132.295 136.405 132.525 ;
        RECT 133.655 131.615 136.405 132.295 ;
        RECT 136.415 131.615 141.925 132.425 ;
        RECT 142.420 132.295 143.765 132.525 ;
        RECT 144.260 132.295 145.605 132.525 ;
        RECT 141.935 131.615 143.765 132.295 ;
        RECT 143.775 131.615 145.605 132.295 ;
        RECT 145.615 131.615 146.985 132.425 ;
        RECT 17.415 131.405 17.585 131.615 ;
        RECT 18.790 131.455 18.910 131.565 ;
        RECT 19.255 131.425 19.425 131.615 ;
        RECT 20.175 131.405 20.345 131.595 ;
        RECT 20.635 131.405 20.805 131.595 ;
        RECT 22.290 131.405 22.460 131.595 ;
        RECT 26.155 131.405 26.325 131.595 ;
        RECT 26.610 131.455 26.730 131.565 ;
        RECT 27.075 131.425 27.245 131.615 ;
        RECT 32.595 131.595 32.760 131.615 ;
        RECT 31.675 131.405 31.845 131.595 ;
        RECT 32.595 131.425 32.765 131.595 ;
        RECT 33.975 131.425 34.145 131.615 ;
        RECT 34.435 131.425 34.605 131.615 ;
        RECT 37.195 131.405 37.365 131.595 ;
        RECT 39.955 131.425 40.125 131.615 ;
        RECT 42.710 131.455 42.830 131.565 ;
        RECT 43.635 131.405 43.805 131.595 ;
        RECT 45.475 131.425 45.645 131.615 ;
        RECT 49.155 131.405 49.325 131.595 ;
        RECT 50.995 131.425 51.165 131.615 ;
        RECT 54.675 131.405 54.845 131.615 ;
        RECT 56.515 131.425 56.685 131.615 ;
        RECT 60.190 131.455 60.310 131.565 ;
        RECT 60.655 131.405 60.825 131.595 ;
        RECT 62.035 131.425 62.205 131.615 ;
        RECT 71.695 131.595 71.845 131.615 ;
        RECT 63.875 131.405 64.045 131.595 ;
        RECT 69.395 131.405 69.565 131.595 ;
        RECT 71.695 131.425 71.865 131.595 ;
        RECT 72.150 131.455 72.270 131.565 ;
        RECT 72.615 131.425 72.785 131.615 ;
        RECT 79.975 131.425 80.145 131.615 ;
        RECT 82.275 131.425 82.445 131.615 ;
        RECT 84.115 131.405 84.285 131.595 ;
        RECT 84.585 131.450 84.745 131.560 ;
        RECT 85.495 131.405 85.665 131.595 ;
        RECT 87.060 131.425 87.230 131.615 ;
        RECT 87.795 131.425 87.965 131.615 ;
        RECT 93.315 131.405 93.485 131.595 ;
        RECT 95.155 131.405 95.325 131.595 ;
        RECT 97.915 131.405 98.085 131.595 ;
        RECT 98.835 131.425 99.005 131.615 ;
        RECT 99.290 131.455 99.410 131.565 ;
        RECT 99.755 131.425 99.925 131.615 ;
        RECT 101.595 131.405 101.765 131.595 ;
        RECT 105.275 131.405 105.445 131.595 ;
        RECT 106.840 131.425 107.010 131.615 ;
        RECT 108.035 131.425 108.205 131.615 ;
        RECT 109.425 131.405 109.595 131.595 ;
        RECT 109.875 131.405 110.045 131.595 ;
        RECT 111.715 131.405 111.885 131.595 ;
        RECT 115.395 131.425 115.565 131.615 ;
        RECT 119.075 131.405 119.245 131.595 ;
        RECT 120.915 131.425 121.085 131.615 ;
        RECT 123.215 131.405 123.385 131.595 ;
        RECT 123.675 131.405 123.845 131.615 ;
        RECT 129.195 131.565 129.365 131.615 ;
        RECT 129.190 131.455 129.365 131.565 ;
        RECT 129.195 131.425 129.365 131.455 ;
        RECT 129.655 131.405 129.825 131.595 ;
        RECT 132.415 131.405 132.585 131.595 ;
        RECT 132.870 131.455 132.990 131.565 ;
        RECT 133.795 131.425 133.965 131.615 ;
        RECT 135.170 131.455 135.290 131.565 ;
        RECT 135.910 131.405 136.080 131.595 ;
        RECT 136.555 131.425 136.725 131.615 ;
        RECT 139.775 131.405 139.945 131.595 ;
        RECT 142.075 131.425 142.245 131.615 ;
        RECT 143.915 131.425 144.085 131.615 ;
        RECT 145.290 131.455 145.410 131.565 ;
        RECT 146.675 131.405 146.845 131.615 ;
        RECT 17.275 130.595 18.645 131.405 ;
        RECT 18.655 130.725 20.485 131.405 ;
        RECT 18.655 130.495 20.000 130.725 ;
        RECT 20.495 130.595 21.865 131.405 ;
        RECT 21.875 130.725 25.775 131.405 ;
        RECT 21.875 130.495 22.805 130.725 ;
        RECT 26.015 130.595 31.525 131.405 ;
        RECT 31.535 130.595 37.045 131.405 ;
        RECT 37.055 130.595 42.565 131.405 ;
        RECT 43.045 130.535 43.475 131.320 ;
        RECT 43.495 130.595 49.005 131.405 ;
        RECT 49.015 130.595 54.525 131.405 ;
        RECT 54.535 130.595 60.045 131.405 ;
        RECT 60.565 130.495 63.725 131.405 ;
        RECT 63.735 130.725 68.550 131.405 ;
        RECT 68.805 130.535 69.235 131.320 ;
        RECT 69.255 130.725 76.985 131.405 ;
        RECT 72.770 130.505 73.680 130.725 ;
        RECT 75.215 130.495 76.985 130.725 ;
        RECT 77.115 130.725 84.425 131.405 ;
        RECT 85.355 130.725 93.085 131.405 ;
        RECT 77.115 130.495 78.465 130.725 ;
        RECT 80.000 130.505 80.910 130.725 ;
        RECT 88.870 130.505 89.780 130.725 ;
        RECT 91.315 130.495 93.085 130.725 ;
        RECT 93.175 130.595 94.545 131.405 ;
        RECT 94.565 130.535 94.995 131.320 ;
        RECT 95.015 130.595 97.765 131.405 ;
        RECT 97.885 130.725 101.350 131.405 ;
        RECT 100.430 130.495 101.350 130.725 ;
        RECT 101.455 130.595 105.125 131.405 ;
        RECT 105.135 130.595 106.505 131.405 ;
        RECT 106.515 130.495 109.725 131.405 ;
        RECT 109.735 130.595 111.565 131.405 ;
        RECT 111.575 130.725 118.885 131.405 ;
        RECT 115.090 130.505 116.000 130.725 ;
        RECT 117.535 130.495 118.885 130.725 ;
        RECT 118.935 130.595 120.305 131.405 ;
        RECT 120.325 130.535 120.755 131.320 ;
        RECT 120.775 130.725 123.525 131.405 ;
        RECT 120.775 130.495 121.705 130.725 ;
        RECT 123.535 130.595 129.045 131.405 ;
        RECT 129.515 130.725 132.265 131.405 ;
        RECT 131.335 130.495 132.265 130.725 ;
        RECT 132.275 130.595 135.025 131.405 ;
        RECT 135.495 130.725 139.395 131.405 ;
        RECT 135.495 130.495 136.425 130.725 ;
        RECT 139.635 130.595 145.145 131.405 ;
        RECT 145.615 130.595 146.985 131.405 ;
      LAYER nwell ;
        RECT 17.080 127.375 147.180 130.205 ;
      LAYER pwell ;
        RECT 17.275 126.175 18.645 126.985 ;
        RECT 18.655 126.855 20.000 127.085 ;
        RECT 20.495 126.855 21.840 127.085 ;
        RECT 18.655 126.175 20.485 126.855 ;
        RECT 20.495 126.175 22.325 126.855 ;
        RECT 22.335 126.175 26.005 126.985 ;
        RECT 27.065 126.855 27.995 127.085 ;
        RECT 26.160 126.175 27.995 126.855 ;
        RECT 28.315 126.175 30.145 126.985 ;
        RECT 30.165 126.260 30.595 127.045 ;
        RECT 30.615 126.175 36.125 126.985 ;
        RECT 36.135 126.175 41.645 126.985 ;
        RECT 41.655 126.175 47.165 126.985 ;
        RECT 47.175 126.175 52.685 126.985 ;
        RECT 52.695 126.175 55.445 126.985 ;
        RECT 55.925 126.260 56.355 127.045 ;
        RECT 56.375 126.175 61.885 126.985 ;
        RECT 61.895 126.175 64.645 126.985 ;
        RECT 64.655 126.855 65.585 127.085 ;
        RECT 64.655 126.175 68.555 126.855 ;
        RECT 68.795 126.175 71.545 126.985 ;
        RECT 71.555 126.855 72.485 127.085 ;
        RECT 71.555 126.175 75.455 126.855 ;
        RECT 75.695 126.175 81.205 126.985 ;
        RECT 81.685 126.260 82.115 127.045 ;
        RECT 82.135 126.855 83.065 127.085 ;
        RECT 82.135 126.175 86.035 126.855 ;
        RECT 86.275 126.175 89.945 126.985 ;
        RECT 89.955 126.175 91.325 126.985 ;
        RECT 96.395 126.855 97.325 127.085 ;
        RECT 100.535 126.855 101.465 127.085 ;
        RECT 91.570 126.175 96.385 126.855 ;
        RECT 96.395 126.175 100.295 126.855 ;
        RECT 100.535 126.175 104.435 126.855 ;
        RECT 104.675 126.175 107.425 126.985 ;
        RECT 107.445 126.260 107.875 127.045 ;
        RECT 110.635 126.855 111.565 127.085 ;
        RECT 108.815 126.175 111.565 126.855 ;
        RECT 111.575 126.855 112.505 127.085 ;
        RECT 111.575 126.175 115.475 126.855 ;
        RECT 115.715 126.175 117.545 126.985 ;
        RECT 117.555 126.175 120.765 127.085 ;
        RECT 124.290 126.855 125.200 127.075 ;
        RECT 126.735 126.855 128.085 127.085 ;
        RECT 120.775 126.175 128.085 126.855 ;
        RECT 128.135 126.175 129.965 126.985 ;
        RECT 132.255 126.855 133.185 127.085 ;
        RECT 130.435 126.175 133.185 126.855 ;
        RECT 133.205 126.260 133.635 127.045 ;
        RECT 133.655 126.175 136.865 127.085 ;
        RECT 140.850 126.855 141.760 127.075 ;
        RECT 143.295 126.855 144.645 127.085 ;
        RECT 137.335 126.175 144.645 126.855 ;
        RECT 145.615 126.175 146.985 126.985 ;
        RECT 17.415 125.965 17.585 126.175 ;
        RECT 18.805 126.010 18.965 126.120 ;
        RECT 19.715 125.965 19.885 126.155 ;
        RECT 20.175 125.985 20.345 126.175 ;
        RECT 21.555 125.965 21.725 126.155 ;
        RECT 22.015 125.985 22.185 126.175 ;
        RECT 22.475 125.985 22.645 126.175 ;
        RECT 26.160 126.155 26.325 126.175 ;
        RECT 26.155 125.985 26.325 126.155 ;
        RECT 28.455 125.985 28.625 126.175 ;
        RECT 29.835 125.965 30.005 126.155 ;
        RECT 30.295 125.965 30.465 126.155 ;
        RECT 30.755 125.985 30.925 126.175 ;
        RECT 34.435 125.965 34.605 126.155 ;
        RECT 36.275 125.985 36.445 126.175 ;
        RECT 39.955 125.965 40.125 126.155 ;
        RECT 41.795 125.985 41.965 126.175 ;
        RECT 42.710 126.015 42.830 126.125 ;
        RECT 43.635 125.965 43.805 126.155 ;
        RECT 47.315 125.985 47.485 126.175 ;
        RECT 49.155 125.965 49.325 126.155 ;
        RECT 52.835 125.985 53.005 126.175 ;
        RECT 54.675 125.965 54.845 126.155 ;
        RECT 55.590 126.015 55.710 126.125 ;
        RECT 56.515 125.985 56.685 126.175 ;
        RECT 60.195 125.965 60.365 126.155 ;
        RECT 62.035 125.985 62.205 126.175 ;
        RECT 65.070 125.985 65.240 126.175 ;
        RECT 65.715 125.965 65.885 126.155 ;
        RECT 68.470 126.015 68.590 126.125 ;
        RECT 68.935 125.985 69.105 126.175 ;
        RECT 69.395 125.965 69.565 126.155 ;
        RECT 71.970 125.985 72.140 126.175 ;
        RECT 74.915 125.965 75.085 126.155 ;
        RECT 75.835 125.985 76.005 126.175 ;
        RECT 80.435 125.965 80.605 126.155 ;
        RECT 81.350 126.015 81.470 126.125 ;
        RECT 82.550 125.985 82.720 126.175 ;
        RECT 85.965 126.010 86.125 126.120 ;
        RECT 86.415 125.985 86.585 126.175 ;
        RECT 86.875 125.965 87.045 126.155 ;
        RECT 89.635 125.965 89.805 126.155 ;
        RECT 90.095 125.985 90.265 126.175 ;
        RECT 95.155 125.965 95.325 126.155 ;
        RECT 96.075 125.985 96.245 126.175 ;
        RECT 96.810 125.985 96.980 126.175 ;
        RECT 100.950 125.985 101.120 126.175 ;
        RECT 103.890 125.965 104.060 126.155 ;
        RECT 104.355 125.965 104.525 126.155 ;
        RECT 104.815 125.985 104.985 126.175 ;
        RECT 108.045 126.020 108.205 126.130 ;
        RECT 108.955 125.985 109.125 126.175 ;
        RECT 109.875 125.965 110.045 126.155 ;
        RECT 111.990 125.985 112.160 126.175 ;
        RECT 113.550 126.015 113.670 126.125 ;
        RECT 114.290 125.965 114.460 126.155 ;
        RECT 115.855 125.985 116.025 126.175 ;
        RECT 117.685 125.985 117.855 126.175 ;
        RECT 118.155 125.965 118.325 126.155 ;
        RECT 119.990 126.015 120.110 126.125 ;
        RECT 120.915 125.985 121.085 126.175 ;
        RECT 121.835 125.965 122.005 126.155 ;
        RECT 127.170 125.965 127.340 126.155 ;
        RECT 128.275 125.985 128.445 126.175 ;
        RECT 130.110 126.015 130.230 126.125 ;
        RECT 130.575 125.985 130.745 126.175 ;
        RECT 131.035 125.965 131.205 126.155 ;
        RECT 132.415 125.965 132.585 126.155 ;
        RECT 133.785 125.985 133.955 126.175 ;
        RECT 137.010 126.015 137.130 126.125 ;
        RECT 137.475 125.985 137.645 126.175 ;
        RECT 139.775 125.965 139.945 126.155 ;
        RECT 141.610 126.015 141.730 126.125 ;
        RECT 142.075 125.965 142.245 126.155 ;
        RECT 143.915 125.965 144.085 126.155 ;
        RECT 144.845 126.020 145.005 126.130 ;
        RECT 146.675 125.965 146.845 126.175 ;
        RECT 17.275 125.155 18.645 125.965 ;
        RECT 19.575 125.285 21.405 125.965 ;
        RECT 21.415 125.155 22.785 125.965 ;
        RECT 22.835 125.285 30.145 125.965 ;
        RECT 22.835 125.055 24.185 125.285 ;
        RECT 25.720 125.065 26.630 125.285 ;
        RECT 30.155 125.055 34.215 125.965 ;
        RECT 34.295 125.155 39.805 125.965 ;
        RECT 39.815 125.155 42.565 125.965 ;
        RECT 43.045 125.095 43.475 125.880 ;
        RECT 43.495 125.155 49.005 125.965 ;
        RECT 49.015 125.155 54.525 125.965 ;
        RECT 54.535 125.155 60.045 125.965 ;
        RECT 60.055 125.155 65.565 125.965 ;
        RECT 65.575 125.155 68.325 125.965 ;
        RECT 68.805 125.095 69.235 125.880 ;
        RECT 69.255 125.155 74.765 125.965 ;
        RECT 74.775 125.155 80.285 125.965 ;
        RECT 80.295 125.155 85.805 125.965 ;
        RECT 86.735 125.155 88.825 125.965 ;
        RECT 89.495 125.285 94.310 125.965 ;
        RECT 94.565 125.095 94.995 125.880 ;
        RECT 95.015 125.285 102.325 125.965 ;
        RECT 98.530 125.065 99.440 125.285 ;
        RECT 100.975 125.055 102.325 125.285 ;
        RECT 102.435 125.055 104.205 125.965 ;
        RECT 104.215 125.155 109.725 125.965 ;
        RECT 109.735 125.155 113.405 125.965 ;
        RECT 113.875 125.285 117.775 125.965 ;
        RECT 113.875 125.055 114.805 125.285 ;
        RECT 118.015 125.155 119.845 125.965 ;
        RECT 120.325 125.095 120.755 125.880 ;
        RECT 121.695 125.285 126.510 125.965 ;
        RECT 126.755 125.285 130.655 125.965 ;
        RECT 126.755 125.055 127.685 125.285 ;
        RECT 130.895 125.155 132.265 125.965 ;
        RECT 132.275 125.285 139.585 125.965 ;
        RECT 135.790 125.065 136.700 125.285 ;
        RECT 138.235 125.055 139.585 125.285 ;
        RECT 139.635 125.155 141.465 125.965 ;
        RECT 141.935 125.285 143.765 125.965 ;
        RECT 143.775 125.285 145.605 125.965 ;
        RECT 142.420 125.055 143.765 125.285 ;
        RECT 144.260 125.055 145.605 125.285 ;
        RECT 145.615 125.155 146.985 125.965 ;
      LAYER nwell ;
        RECT 17.080 121.935 147.180 124.765 ;
      LAYER pwell ;
        RECT 17.275 120.735 18.645 121.545 ;
        RECT 22.630 121.415 23.540 121.635 ;
        RECT 25.075 121.415 26.425 121.645 ;
        RECT 19.115 120.735 26.425 121.415 ;
        RECT 26.935 121.415 28.300 121.645 ;
        RECT 26.935 120.735 30.145 121.415 ;
        RECT 30.165 120.820 30.595 121.605 ;
        RECT 34.130 121.415 35.040 121.635 ;
        RECT 36.575 121.415 37.925 121.645 ;
        RECT 30.615 120.735 37.925 121.415 ;
        RECT 37.975 120.735 43.485 121.545 ;
        RECT 43.495 120.735 49.005 121.545 ;
        RECT 49.015 120.735 54.525 121.545 ;
        RECT 54.535 120.735 55.905 121.545 ;
        RECT 55.925 120.820 56.355 121.605 ;
        RECT 56.375 120.735 61.885 121.545 ;
        RECT 61.895 120.735 67.405 121.545 ;
        RECT 67.415 120.735 72.925 121.545 ;
        RECT 72.935 120.735 78.445 121.545 ;
        RECT 78.455 120.735 81.205 121.545 ;
        RECT 81.685 120.820 82.115 121.605 ;
        RECT 82.135 120.735 85.805 121.545 ;
        RECT 88.555 121.415 89.485 121.645 ;
        RECT 86.735 120.735 89.485 121.415 ;
        RECT 90.615 120.735 92.705 121.545 ;
        RECT 96.690 121.415 97.600 121.635 ;
        RECT 99.135 121.415 100.485 121.645 ;
        RECT 93.175 120.735 100.485 121.415 ;
        RECT 100.535 120.965 105.125 121.645 ;
        RECT 101.495 120.735 105.125 120.965 ;
        RECT 105.135 120.735 106.965 121.415 ;
        RECT 107.445 120.820 107.875 121.605 ;
        RECT 107.895 120.735 111.105 121.645 ;
        RECT 111.115 120.735 112.945 121.545 ;
        RECT 116.930 121.415 117.840 121.635 ;
        RECT 119.375 121.415 120.725 121.645 ;
        RECT 113.415 120.735 120.725 121.415 ;
        RECT 120.775 120.735 125.590 121.415 ;
        RECT 125.835 120.735 129.505 121.545 ;
        RECT 129.515 120.735 133.170 121.645 ;
        RECT 133.205 120.820 133.635 121.605 ;
        RECT 133.655 121.415 134.585 121.645 ;
        RECT 133.655 120.735 137.555 121.415 ;
        RECT 137.795 120.735 141.465 121.545 ;
        RECT 142.420 121.415 143.765 121.645 ;
        RECT 144.260 121.415 145.605 121.645 ;
        RECT 141.935 120.735 143.765 121.415 ;
        RECT 143.775 120.735 145.605 121.415 ;
        RECT 145.615 120.735 146.985 121.545 ;
        RECT 17.415 120.525 17.585 120.735 ;
        RECT 18.805 120.685 18.975 120.715 ;
        RECT 18.790 120.575 18.975 120.685 ;
        RECT 18.805 120.525 18.975 120.575 ;
        RECT 19.255 120.545 19.425 120.735 ;
        RECT 20.185 120.525 20.355 120.715 ;
        RECT 21.830 120.525 22.000 120.715 ;
        RECT 25.690 120.575 25.810 120.685 ;
        RECT 26.155 120.525 26.325 120.715 ;
        RECT 26.610 120.575 26.730 120.685 ;
        RECT 29.830 120.545 30.000 120.735 ;
        RECT 30.755 120.545 30.925 120.735 ;
        RECT 33.520 120.525 33.690 120.715 ;
        RECT 36.735 120.525 36.905 120.715 ;
        RECT 38.115 120.545 38.285 120.735 ;
        RECT 42.265 120.570 42.425 120.680 ;
        RECT 43.635 120.525 43.805 120.735 ;
        RECT 49.155 120.525 49.325 120.735 ;
        RECT 54.675 120.525 54.845 120.735 ;
        RECT 56.515 120.545 56.685 120.735 ;
        RECT 60.195 120.525 60.365 120.715 ;
        RECT 62.035 120.545 62.205 120.735 ;
        RECT 65.715 120.525 65.885 120.715 ;
        RECT 67.555 120.545 67.725 120.735 ;
        RECT 68.470 120.575 68.590 120.685 ;
        RECT 69.395 120.525 69.565 120.715 ;
        RECT 73.075 120.545 73.245 120.735 ;
        RECT 73.995 120.525 74.165 120.715 ;
        RECT 76.755 120.525 76.925 120.715 ;
        RECT 78.410 120.525 78.580 120.715 ;
        RECT 78.595 120.545 78.765 120.735 ;
        RECT 81.350 120.575 81.470 120.685 ;
        RECT 82.275 120.525 82.445 120.735 ;
        RECT 84.110 120.575 84.230 120.685 ;
        RECT 84.850 120.525 85.020 120.715 ;
        RECT 85.965 120.580 86.125 120.690 ;
        RECT 86.875 120.545 87.045 120.735 ;
        RECT 88.715 120.525 88.885 120.715 ;
        RECT 89.630 120.575 89.750 120.685 ;
        RECT 90.560 120.525 90.730 120.715 ;
        RECT 92.395 120.545 92.565 120.735 ;
        RECT 92.850 120.575 92.970 120.685 ;
        RECT 93.315 120.545 93.485 120.735 ;
        RECT 95.165 120.570 95.325 120.680 ;
        RECT 97.455 120.525 97.625 120.715 ;
        RECT 97.920 120.525 98.090 120.715 ;
        RECT 102.515 120.545 102.685 120.715 ;
        RECT 104.810 120.545 104.980 120.735 ;
        RECT 106.655 120.545 106.825 120.735 ;
        RECT 107.110 120.575 107.230 120.685 ;
        RECT 108.025 120.545 108.195 120.735 ;
        RECT 102.545 120.525 102.685 120.545 ;
        RECT 110.980 120.525 111.150 120.715 ;
        RECT 111.255 120.545 111.425 120.735 ;
        RECT 111.725 120.570 111.885 120.680 ;
        RECT 112.635 120.525 112.805 120.715 ;
        RECT 113.090 120.575 113.210 120.685 ;
        RECT 113.555 120.545 113.725 120.735 ;
        RECT 115.395 120.525 115.565 120.715 ;
        RECT 119.075 120.525 119.245 120.715 ;
        RECT 120.915 120.685 121.085 120.735 ;
        RECT 120.910 120.575 121.085 120.685 ;
        RECT 120.915 120.545 121.085 120.575 ;
        RECT 121.375 120.525 121.545 120.715 ;
        RECT 125.975 120.545 126.145 120.735 ;
        RECT 129.010 120.525 129.180 120.715 ;
        RECT 129.660 120.545 129.830 120.735 ;
        RECT 132.875 120.525 133.045 120.715 ;
        RECT 134.070 120.545 134.240 120.735 ;
        RECT 134.715 120.525 134.885 120.715 ;
        RECT 137.475 120.525 137.645 120.715 ;
        RECT 137.935 120.545 138.105 120.735 ;
        RECT 141.610 120.575 141.730 120.685 ;
        RECT 142.075 120.545 142.245 120.735 ;
        RECT 143.915 120.545 144.085 120.735 ;
        RECT 144.845 120.570 145.005 120.680 ;
        RECT 146.675 120.525 146.845 120.735 ;
        RECT 17.275 119.715 18.645 120.525 ;
        RECT 18.655 119.745 20.025 120.525 ;
        RECT 20.035 119.745 21.405 120.525 ;
        RECT 21.415 119.845 25.315 120.525 ;
        RECT 26.015 119.845 33.325 120.525 ;
        RECT 33.375 119.845 36.585 120.525 ;
        RECT 21.415 119.615 22.345 119.845 ;
        RECT 29.530 119.625 30.440 119.845 ;
        RECT 31.975 119.615 33.325 119.845 ;
        RECT 35.220 119.615 36.585 119.845 ;
        RECT 36.595 119.715 42.105 120.525 ;
        RECT 43.045 119.655 43.475 120.440 ;
        RECT 43.495 119.715 49.005 120.525 ;
        RECT 49.015 119.715 54.525 120.525 ;
        RECT 54.535 119.715 60.045 120.525 ;
        RECT 60.055 119.715 65.565 120.525 ;
        RECT 65.575 119.715 68.325 120.525 ;
        RECT 68.805 119.655 69.235 120.440 ;
        RECT 69.255 119.715 72.925 120.525 ;
        RECT 73.855 119.845 76.605 120.525 ;
        RECT 75.675 119.615 76.605 119.845 ;
        RECT 76.615 119.715 77.985 120.525 ;
        RECT 77.995 119.845 81.895 120.525 ;
        RECT 77.995 119.615 78.925 119.845 ;
        RECT 82.135 119.715 83.965 120.525 ;
        RECT 84.435 119.845 88.335 120.525 ;
        RECT 84.435 119.615 85.365 119.845 ;
        RECT 88.575 119.715 90.405 120.525 ;
        RECT 90.415 119.615 94.285 120.525 ;
        RECT 94.565 119.655 94.995 120.440 ;
        RECT 95.935 119.845 97.765 120.525 ;
        RECT 97.775 120.295 101.405 120.525 ;
        RECT 102.545 120.295 106.315 120.525 ;
        RECT 95.935 119.615 97.280 119.845 ;
        RECT 97.775 119.615 102.365 120.295 ;
        RECT 102.545 119.615 106.895 120.295 ;
        RECT 107.665 119.845 111.565 120.525 ;
        RECT 112.495 119.845 115.245 120.525 ;
        RECT 110.635 119.615 111.565 119.845 ;
        RECT 114.315 119.615 115.245 119.845 ;
        RECT 115.255 119.715 118.925 120.525 ;
        RECT 118.935 119.715 120.305 120.525 ;
        RECT 120.325 119.655 120.755 120.440 ;
        RECT 121.235 119.845 128.545 120.525 ;
        RECT 124.750 119.625 125.660 119.845 ;
        RECT 127.195 119.615 128.545 119.845 ;
        RECT 128.595 119.845 132.495 120.525 ;
        RECT 128.595 119.615 129.525 119.845 ;
        RECT 132.735 119.715 134.565 120.525 ;
        RECT 134.575 119.845 137.325 120.525 ;
        RECT 137.335 119.845 144.645 120.525 ;
        RECT 136.395 119.615 137.325 119.845 ;
        RECT 140.850 119.625 141.760 119.845 ;
        RECT 143.295 119.615 144.645 119.845 ;
        RECT 145.615 119.715 146.985 120.525 ;
      LAYER nwell ;
        RECT 17.080 116.495 147.180 119.325 ;
      LAYER pwell ;
        RECT 17.275 115.295 18.645 116.105 ;
        RECT 18.655 115.295 24.165 116.105 ;
        RECT 24.175 115.295 27.845 116.105 ;
        RECT 28.795 115.295 30.145 116.205 ;
        RECT 30.165 115.380 30.595 116.165 ;
        RECT 30.615 115.295 36.125 116.105 ;
        RECT 36.135 115.295 41.645 116.105 ;
        RECT 41.655 115.295 47.165 116.105 ;
        RECT 47.175 115.295 52.685 116.105 ;
        RECT 52.695 115.295 55.445 116.105 ;
        RECT 55.925 115.380 56.355 116.165 ;
        RECT 56.375 115.295 61.885 116.105 ;
        RECT 61.895 115.295 67.405 116.105 ;
        RECT 67.415 115.295 71.085 116.105 ;
        RECT 72.915 115.975 73.845 116.205 ;
        RECT 77.370 115.975 78.280 116.195 ;
        RECT 79.815 115.975 81.165 116.205 ;
        RECT 71.095 115.295 73.845 115.975 ;
        RECT 73.855 115.295 81.165 115.975 ;
        RECT 81.685 115.380 82.115 116.165 ;
        RECT 85.650 115.975 86.560 116.195 ;
        RECT 88.095 115.975 89.445 116.205 ;
        RECT 82.135 115.295 89.445 115.975 ;
        RECT 90.415 115.975 91.345 116.205 ;
        RECT 90.415 115.295 94.315 115.975 ;
        RECT 94.555 115.295 98.425 116.205 ;
        RECT 98.955 115.295 102.825 116.205 ;
        RECT 103.295 115.975 104.225 116.205 ;
        RECT 103.295 115.295 107.195 115.975 ;
        RECT 107.445 115.380 107.875 116.165 ;
        RECT 107.935 115.975 109.285 116.205 ;
        RECT 110.820 115.975 111.730 116.195 ;
        RECT 107.935 115.295 115.245 115.975 ;
        RECT 115.255 115.295 120.765 116.105 ;
        RECT 123.055 115.975 123.985 116.205 ;
        RECT 121.235 115.295 123.985 115.975 ;
        RECT 123.995 115.975 124.925 116.205 ;
        RECT 123.995 115.295 126.745 115.975 ;
        RECT 126.755 115.295 132.265 116.105 ;
        RECT 133.205 115.380 133.635 116.165 ;
        RECT 133.655 115.295 136.405 116.105 ;
        RECT 136.415 115.975 137.345 116.205 ;
        RECT 136.415 115.295 140.315 115.975 ;
        RECT 140.570 115.295 144.225 116.205 ;
        RECT 144.235 115.295 145.605 116.105 ;
        RECT 145.615 115.295 146.985 116.105 ;
        RECT 17.415 115.085 17.585 115.295 ;
        RECT 18.795 115.105 18.965 115.295 ;
        RECT 20.175 115.085 20.345 115.275 ;
        RECT 20.635 115.085 20.805 115.275 ;
        RECT 24.315 115.105 24.485 115.295 ;
        RECT 25.880 115.085 26.050 115.275 ;
        RECT 26.610 115.135 26.730 115.245 ;
        RECT 27.075 115.085 27.245 115.275 ;
        RECT 28.005 115.140 28.165 115.250 ;
        RECT 29.830 115.105 30.000 115.295 ;
        RECT 30.755 115.105 30.925 115.295 ;
        RECT 34.435 115.085 34.605 115.275 ;
        RECT 36.275 115.105 36.445 115.295 ;
        RECT 39.955 115.085 40.125 115.275 ;
        RECT 41.795 115.105 41.965 115.295 ;
        RECT 42.710 115.135 42.830 115.245 ;
        RECT 43.635 115.085 43.805 115.275 ;
        RECT 47.315 115.105 47.485 115.295 ;
        RECT 49.155 115.085 49.325 115.275 ;
        RECT 52.835 115.105 53.005 115.295 ;
        RECT 54.675 115.085 54.845 115.275 ;
        RECT 55.590 115.135 55.710 115.245 ;
        RECT 56.515 115.105 56.685 115.295 ;
        RECT 60.195 115.085 60.365 115.275 ;
        RECT 62.035 115.105 62.205 115.295 ;
        RECT 65.715 115.085 65.885 115.275 ;
        RECT 67.555 115.105 67.725 115.295 ;
        RECT 68.470 115.135 68.590 115.245 ;
        RECT 69.395 115.085 69.565 115.275 ;
        RECT 71.235 115.085 71.405 115.295 ;
        RECT 73.995 115.105 74.165 115.295 ;
        RECT 78.870 115.085 79.040 115.275 ;
        RECT 81.350 115.135 81.470 115.245 ;
        RECT 82.275 115.105 82.445 115.295 ;
        RECT 82.740 115.085 82.910 115.275 ;
        RECT 86.410 115.135 86.530 115.245 ;
        RECT 86.875 115.085 87.045 115.275 ;
        RECT 89.645 115.140 89.805 115.250 ;
        RECT 90.830 115.105 91.000 115.295 ;
        RECT 94.230 115.135 94.350 115.245 ;
        RECT 94.700 115.105 94.870 115.295 ;
        RECT 102.510 115.275 102.680 115.295 ;
        RECT 98.830 115.085 99.000 115.275 ;
        RECT 99.295 115.085 99.465 115.275 ;
        RECT 102.055 115.085 102.225 115.275 ;
        RECT 102.510 115.105 102.685 115.275 ;
        RECT 102.970 115.135 103.090 115.245 ;
        RECT 103.710 115.105 103.880 115.295 ;
        RECT 102.515 115.085 102.685 115.105 ;
        RECT 109.875 115.085 110.045 115.275 ;
        RECT 113.095 115.085 113.265 115.275 ;
        RECT 114.935 115.105 115.105 115.295 ;
        RECT 115.395 115.105 115.565 115.295 ;
        RECT 118.615 115.085 118.785 115.275 ;
        RECT 120.915 115.245 121.085 115.275 ;
        RECT 120.910 115.135 121.085 115.245 ;
        RECT 120.915 115.085 121.085 115.135 ;
        RECT 121.375 115.105 121.545 115.295 ;
        RECT 122.295 115.085 122.465 115.275 ;
        RECT 126.435 115.105 126.605 115.295 ;
        RECT 126.895 115.105 127.065 115.295 ;
        RECT 129.930 115.085 130.100 115.275 ;
        RECT 132.425 115.140 132.585 115.250 ;
        RECT 133.795 115.085 133.965 115.295 ;
        RECT 135.910 115.085 136.080 115.275 ;
        RECT 136.830 115.105 137.000 115.295 ;
        RECT 143.910 115.275 144.080 115.295 ;
        RECT 140.050 115.085 140.220 115.275 ;
        RECT 143.910 115.105 144.085 115.275 ;
        RECT 144.375 115.105 144.545 115.295 ;
        RECT 143.915 115.085 144.085 115.105 ;
        RECT 146.675 115.085 146.845 115.295 ;
        RECT 17.275 114.275 18.645 115.085 ;
        RECT 18.655 114.405 20.485 115.085 ;
        RECT 18.655 114.175 20.000 114.405 ;
        RECT 20.495 114.275 22.325 115.085 ;
        RECT 22.565 114.405 26.465 115.085 ;
        RECT 26.935 114.405 34.245 115.085 ;
        RECT 25.535 114.175 26.465 114.405 ;
        RECT 30.450 114.185 31.360 114.405 ;
        RECT 32.895 114.175 34.245 114.405 ;
        RECT 34.295 114.275 39.805 115.085 ;
        RECT 39.815 114.275 42.565 115.085 ;
        RECT 43.045 114.215 43.475 115.000 ;
        RECT 43.495 114.275 49.005 115.085 ;
        RECT 49.015 114.275 54.525 115.085 ;
        RECT 54.535 114.275 60.045 115.085 ;
        RECT 60.055 114.275 65.565 115.085 ;
        RECT 65.575 114.275 68.325 115.085 ;
        RECT 68.805 114.215 69.235 115.000 ;
        RECT 69.255 114.275 71.085 115.085 ;
        RECT 71.095 114.405 78.405 115.085 ;
        RECT 74.610 114.185 75.520 114.405 ;
        RECT 77.055 114.175 78.405 114.405 ;
        RECT 78.455 114.405 82.355 115.085 ;
        RECT 78.455 114.175 79.385 114.405 ;
        RECT 82.595 114.175 86.250 115.085 ;
        RECT 86.735 114.405 94.045 115.085 ;
        RECT 90.250 114.185 91.160 114.405 ;
        RECT 92.695 114.175 94.045 114.405 ;
        RECT 94.565 114.215 94.995 115.000 ;
        RECT 95.275 114.175 99.145 115.085 ;
        RECT 99.155 114.275 100.525 115.085 ;
        RECT 100.535 114.405 102.365 115.085 ;
        RECT 102.375 114.405 109.685 115.085 ;
        RECT 105.890 114.185 106.800 114.405 ;
        RECT 108.335 114.175 109.685 114.405 ;
        RECT 109.735 114.175 112.945 115.085 ;
        RECT 112.955 114.275 118.465 115.085 ;
        RECT 118.475 114.275 120.305 115.085 ;
        RECT 120.325 114.215 120.755 115.000 ;
        RECT 120.775 114.275 122.145 115.085 ;
        RECT 122.155 114.405 129.465 115.085 ;
        RECT 125.670 114.185 126.580 114.405 ;
        RECT 128.115 114.175 129.465 114.405 ;
        RECT 129.515 114.405 133.415 115.085 ;
        RECT 129.515 114.175 130.445 114.405 ;
        RECT 133.655 114.275 135.485 115.085 ;
        RECT 135.495 114.405 139.395 115.085 ;
        RECT 139.635 114.405 143.535 115.085 ;
        RECT 143.775 114.405 145.605 115.085 ;
        RECT 135.495 114.175 136.425 114.405 ;
        RECT 139.635 114.175 140.565 114.405 ;
        RECT 144.260 114.175 145.605 114.405 ;
        RECT 145.615 114.275 146.985 115.085 ;
      LAYER nwell ;
        RECT 17.080 111.055 147.180 113.885 ;
      LAYER pwell ;
        RECT 17.275 109.855 18.645 110.665 ;
        RECT 19.155 110.535 20.505 110.765 ;
        RECT 22.040 110.535 22.950 110.755 ;
        RECT 19.155 109.855 26.465 110.535 ;
        RECT 26.475 109.855 30.145 110.665 ;
        RECT 30.165 109.940 30.595 110.725 ;
        RECT 30.615 110.535 31.545 110.765 ;
        RECT 30.615 109.855 34.515 110.535 ;
        RECT 34.755 109.855 40.265 110.665 ;
        RECT 40.275 109.855 45.785 110.665 ;
        RECT 45.795 109.855 51.305 110.665 ;
        RECT 51.315 109.855 54.985 110.665 ;
        RECT 55.925 109.940 56.355 110.725 ;
        RECT 56.375 109.855 61.885 110.665 ;
        RECT 61.895 109.855 63.265 110.665 ;
        RECT 66.790 110.535 67.700 110.755 ;
        RECT 69.235 110.535 70.585 110.765 ;
        RECT 63.275 109.855 70.585 110.535 ;
        RECT 70.635 110.535 71.565 110.765 ;
        RECT 70.635 109.855 74.535 110.535 ;
        RECT 74.775 109.855 80.285 110.665 ;
        RECT 80.295 109.855 81.665 110.665 ;
        RECT 81.685 109.940 82.115 110.725 ;
        RECT 83.955 110.535 84.885 110.765 ;
        RECT 82.135 109.855 84.885 110.535 ;
        RECT 84.895 109.855 88.565 110.665 ;
        RECT 88.575 109.855 91.785 110.765 ;
        RECT 91.795 109.855 97.305 110.665 ;
        RECT 97.315 109.855 102.825 110.665 ;
        RECT 102.835 110.535 103.765 110.765 ;
        RECT 102.835 109.855 105.585 110.535 ;
        RECT 105.595 109.855 107.425 110.665 ;
        RECT 107.445 109.940 107.875 110.725 ;
        RECT 109.715 110.535 110.645 110.765 ;
        RECT 107.895 109.855 110.645 110.535 ;
        RECT 110.655 109.855 112.485 110.665 ;
        RECT 116.155 110.535 117.085 110.765 ;
        RECT 120.610 110.535 121.520 110.755 ;
        RECT 123.055 110.535 124.405 110.765 ;
        RECT 113.185 109.855 117.085 110.535 ;
        RECT 117.095 109.855 124.405 110.535 ;
        RECT 124.455 109.855 129.965 110.665 ;
        RECT 132.255 110.535 133.185 110.765 ;
        RECT 130.435 109.855 133.185 110.535 ;
        RECT 133.205 109.940 133.635 110.725 ;
        RECT 133.655 109.855 135.485 110.665 ;
        RECT 139.470 110.535 140.380 110.755 ;
        RECT 141.915 110.535 143.265 110.765 ;
        RECT 144.260 110.535 145.605 110.765 ;
        RECT 135.955 109.855 143.265 110.535 ;
        RECT 143.775 109.855 145.605 110.535 ;
        RECT 145.615 109.855 146.985 110.665 ;
        RECT 17.415 109.645 17.585 109.855 ;
        RECT 18.790 109.695 18.910 109.805 ;
        RECT 20.175 109.645 20.345 109.835 ;
        RECT 20.630 109.695 20.750 109.805 ;
        RECT 26.155 109.665 26.325 109.855 ;
        RECT 26.615 109.665 26.785 109.855 ;
        RECT 27.995 109.645 28.165 109.835 ;
        RECT 28.730 109.645 28.900 109.835 ;
        RECT 31.030 109.665 31.200 109.855 ;
        RECT 32.595 109.645 32.765 109.835 ;
        RECT 34.895 109.665 35.065 109.855 ;
        RECT 38.115 109.645 38.285 109.835 ;
        RECT 40.415 109.665 40.585 109.855 ;
        RECT 41.795 109.645 41.965 109.835 ;
        RECT 43.635 109.645 43.805 109.835 ;
        RECT 45.935 109.665 46.105 109.855 ;
        RECT 49.155 109.645 49.325 109.835 ;
        RECT 51.455 109.665 51.625 109.855 ;
        RECT 54.675 109.645 54.845 109.835 ;
        RECT 55.145 109.700 55.305 109.810 ;
        RECT 56.515 109.665 56.685 109.855 ;
        RECT 60.195 109.645 60.365 109.835 ;
        RECT 62.035 109.665 62.205 109.855 ;
        RECT 63.415 109.665 63.585 109.855 ;
        RECT 63.870 109.695 63.990 109.805 ;
        RECT 66.635 109.645 66.805 109.835 ;
        RECT 67.095 109.645 67.265 109.835 ;
        RECT 69.395 109.645 69.565 109.835 ;
        RECT 71.050 109.665 71.220 109.855 ;
        RECT 74.915 109.645 75.085 109.855 ;
        RECT 80.435 109.645 80.605 109.855 ;
        RECT 82.275 109.665 82.445 109.855 ;
        RECT 85.035 109.665 85.205 109.855 ;
        RECT 85.955 109.645 86.125 109.835 ;
        RECT 91.475 109.645 91.645 109.855 ;
        RECT 91.935 109.665 92.105 109.855 ;
        RECT 94.230 109.695 94.350 109.805 ;
        RECT 95.155 109.645 95.325 109.835 ;
        RECT 97.455 109.665 97.625 109.855 ;
        RECT 100.675 109.645 100.845 109.835 ;
        RECT 105.275 109.665 105.445 109.855 ;
        RECT 105.735 109.665 105.905 109.855 ;
        RECT 106.205 109.690 106.365 109.800 ;
        RECT 107.115 109.645 107.285 109.835 ;
        RECT 108.035 109.665 108.205 109.855 ;
        RECT 109.875 109.645 110.045 109.835 ;
        RECT 110.795 109.665 110.965 109.855 ;
        RECT 112.630 109.695 112.750 109.805 ;
        RECT 115.405 109.690 115.565 109.800 ;
        RECT 116.315 109.645 116.485 109.835 ;
        RECT 116.500 109.665 116.670 109.855 ;
        RECT 117.235 109.665 117.405 109.855 ;
        RECT 119.075 109.645 119.245 109.835 ;
        RECT 120.915 109.645 121.085 109.835 ;
        RECT 124.595 109.665 124.765 109.855 ;
        RECT 126.435 109.645 126.605 109.835 ;
        RECT 130.110 109.695 130.230 109.805 ;
        RECT 130.575 109.665 130.745 109.855 ;
        RECT 131.955 109.645 132.125 109.835 ;
        RECT 133.795 109.645 133.965 109.855 ;
        RECT 135.630 109.695 135.750 109.805 ;
        RECT 136.095 109.665 136.265 109.855 ;
        RECT 136.555 109.645 136.725 109.835 ;
        RECT 143.450 109.695 143.570 109.805 ;
        RECT 143.915 109.645 144.085 109.855 ;
        RECT 146.675 109.645 146.845 109.855 ;
        RECT 17.275 108.835 18.645 109.645 ;
        RECT 18.655 108.965 20.485 109.645 ;
        RECT 20.995 108.965 28.305 109.645 ;
        RECT 28.315 108.965 32.215 109.645 ;
        RECT 18.655 108.735 20.000 108.965 ;
        RECT 20.995 108.735 22.345 108.965 ;
        RECT 23.880 108.745 24.790 108.965 ;
        RECT 28.315 108.735 29.245 108.965 ;
        RECT 32.455 108.835 37.965 109.645 ;
        RECT 37.975 108.835 41.645 109.645 ;
        RECT 41.655 108.835 43.025 109.645 ;
        RECT 43.045 108.775 43.475 109.560 ;
        RECT 43.495 108.835 49.005 109.645 ;
        RECT 49.015 108.835 54.525 109.645 ;
        RECT 54.535 108.835 60.045 109.645 ;
        RECT 60.055 108.835 63.725 109.645 ;
        RECT 64.195 108.965 66.945 109.645 ;
        RECT 64.195 108.735 65.125 108.965 ;
        RECT 66.955 108.835 68.785 109.645 ;
        RECT 68.805 108.775 69.235 109.560 ;
        RECT 69.255 108.835 74.765 109.645 ;
        RECT 74.775 108.835 80.285 109.645 ;
        RECT 80.295 108.835 85.805 109.645 ;
        RECT 85.815 108.835 91.325 109.645 ;
        RECT 91.335 108.835 94.085 109.645 ;
        RECT 94.565 108.775 94.995 109.560 ;
        RECT 95.015 108.835 100.525 109.645 ;
        RECT 100.535 108.835 106.045 109.645 ;
        RECT 106.975 108.965 109.725 109.645 ;
        RECT 108.795 108.735 109.725 108.965 ;
        RECT 109.735 108.835 115.245 109.645 ;
        RECT 116.175 108.965 118.925 109.645 ;
        RECT 117.995 108.735 118.925 108.965 ;
        RECT 118.935 108.835 120.305 109.645 ;
        RECT 120.325 108.775 120.755 109.560 ;
        RECT 120.775 108.835 126.285 109.645 ;
        RECT 126.295 108.835 131.805 109.645 ;
        RECT 131.815 108.835 133.645 109.645 ;
        RECT 133.655 108.965 136.405 109.645 ;
        RECT 136.415 108.965 143.725 109.645 ;
        RECT 143.775 108.965 145.605 109.645 ;
        RECT 135.475 108.735 136.405 108.965 ;
        RECT 139.930 108.745 140.840 108.965 ;
        RECT 142.375 108.735 143.725 108.965 ;
        RECT 144.260 108.735 145.605 108.965 ;
        RECT 145.615 108.835 146.985 109.645 ;
      LAYER nwell ;
        RECT 17.080 105.615 147.180 108.445 ;
      LAYER pwell ;
        RECT 17.275 104.415 18.645 105.225 ;
        RECT 19.155 105.095 20.505 105.325 ;
        RECT 22.040 105.095 22.950 105.315 ;
        RECT 19.155 104.415 26.465 105.095 ;
        RECT 26.475 104.415 27.845 105.225 ;
        RECT 27.855 105.125 28.810 105.325 ;
        RECT 27.855 104.445 30.135 105.125 ;
        RECT 30.165 104.500 30.595 105.285 ;
        RECT 27.855 104.415 28.810 104.445 ;
        RECT 17.415 104.205 17.585 104.415 ;
        RECT 18.790 104.255 18.910 104.365 ;
        RECT 20.175 104.205 20.345 104.395 ;
        RECT 22.015 104.205 22.185 104.395 ;
        RECT 25.880 104.205 26.050 104.395 ;
        RECT 26.155 104.225 26.325 104.415 ;
        RECT 26.615 104.225 26.785 104.415 ;
        RECT 26.890 104.205 27.060 104.395 ;
        RECT 29.840 104.225 30.010 104.445 ;
        RECT 30.695 104.415 34.145 105.325 ;
        RECT 36.100 105.125 37.045 105.325 ;
        RECT 34.295 104.445 37.045 105.125 ;
        RECT 30.755 104.365 30.925 104.415 ;
        RECT 30.750 104.255 30.925 104.365 ;
        RECT 30.755 104.225 30.925 104.255 ;
        RECT 31.220 104.205 31.390 104.395 ;
        RECT 34.440 104.225 34.610 104.445 ;
        RECT 36.100 104.415 37.045 104.445 ;
        RECT 37.055 104.415 42.565 105.225 ;
        RECT 42.575 104.415 48.085 105.225 ;
        RECT 48.095 104.415 53.605 105.225 ;
        RECT 53.615 104.415 55.445 105.225 ;
        RECT 55.925 104.500 56.355 105.285 ;
        RECT 56.375 104.415 61.885 105.225 ;
        RECT 63.715 105.095 64.645 105.325 ;
        RECT 61.895 104.415 64.645 105.095 ;
        RECT 64.655 104.415 67.405 105.225 ;
        RECT 67.415 105.095 68.345 105.325 ;
        RECT 67.415 104.415 71.315 105.095 ;
        RECT 71.555 104.415 74.765 105.325 ;
        RECT 74.775 104.415 78.445 105.225 ;
        RECT 80.735 105.095 81.665 105.325 ;
        RECT 78.915 104.415 81.665 105.095 ;
        RECT 81.685 104.500 82.115 105.285 ;
        RECT 82.135 104.415 83.965 105.225 ;
        RECT 83.975 105.095 84.905 105.325 ;
        RECT 83.975 104.415 87.875 105.095 ;
        RECT 88.115 104.415 89.945 105.225 ;
        RECT 90.415 104.415 94.070 105.325 ;
        RECT 94.095 104.415 95.465 105.225 ;
        RECT 97.315 105.095 101.245 105.325 ;
        RECT 101.915 105.095 102.845 105.325 ;
        RECT 95.475 104.415 97.305 105.095 ;
        RECT 97.315 104.415 101.730 105.095 ;
        RECT 101.915 104.415 105.815 105.095 ;
        RECT 106.055 104.415 107.425 105.225 ;
        RECT 107.445 104.500 107.875 105.285 ;
        RECT 108.355 105.095 109.285 105.325 ;
        RECT 108.355 104.415 112.255 105.095 ;
        RECT 112.495 104.415 114.325 105.225 ;
        RECT 114.335 104.415 117.990 105.325 ;
        RECT 118.015 104.415 123.525 105.225 ;
        RECT 123.535 104.415 126.285 105.225 ;
        RECT 128.115 105.095 129.045 105.325 ;
        RECT 126.295 104.415 129.045 105.095 ;
        RECT 129.055 104.415 130.885 105.095 ;
        RECT 130.895 104.415 132.725 105.095 ;
        RECT 133.205 104.500 133.635 105.285 ;
        RECT 135.475 105.095 136.405 105.325 ;
        RECT 133.655 104.415 136.405 105.095 ;
        RECT 136.415 104.415 139.625 105.325 ;
        RECT 139.635 104.415 141.465 105.225 ;
        RECT 142.420 105.095 143.765 105.325 ;
        RECT 144.260 105.095 145.605 105.325 ;
        RECT 141.935 104.415 143.765 105.095 ;
        RECT 143.775 104.415 145.605 105.095 ;
        RECT 145.615 104.415 146.985 105.225 ;
        RECT 17.275 103.395 18.645 104.205 ;
        RECT 18.655 103.525 20.485 104.205 ;
        RECT 20.495 103.525 22.325 104.205 ;
        RECT 22.565 103.525 26.465 104.205 ;
        RECT 18.655 103.295 20.000 103.525 ;
        RECT 20.495 103.295 21.840 103.525 ;
        RECT 25.535 103.295 26.465 103.525 ;
        RECT 26.475 103.525 30.375 104.205 ;
        RECT 26.475 103.295 27.405 103.525 ;
        RECT 31.075 103.295 32.425 104.205 ;
        RECT 32.455 104.175 33.405 104.205 ;
        RECT 35.810 104.175 35.980 104.395 ;
        RECT 36.270 104.255 36.390 104.365 ;
        RECT 36.735 104.205 36.905 104.395 ;
        RECT 37.195 104.225 37.365 104.415 ;
        RECT 39.950 104.255 40.070 104.365 ;
        RECT 41.330 104.205 41.500 104.395 ;
        RECT 41.795 104.205 41.965 104.395 ;
        RECT 42.715 104.225 42.885 104.415 ;
        RECT 43.635 104.205 43.805 104.395 ;
        RECT 48.235 104.225 48.405 104.415 ;
        RECT 49.155 104.205 49.325 104.395 ;
        RECT 53.755 104.225 53.925 104.415 ;
        RECT 54.675 104.205 54.845 104.395 ;
        RECT 55.590 104.255 55.710 104.365 ;
        RECT 56.515 104.225 56.685 104.415 ;
        RECT 58.350 104.255 58.470 104.365 ;
        RECT 61.115 104.205 61.285 104.395 ;
        RECT 61.575 104.205 61.745 104.395 ;
        RECT 62.035 104.225 62.205 104.415 ;
        RECT 64.795 104.225 64.965 104.415 ;
        RECT 67.830 104.225 68.000 104.415 ;
        RECT 69.670 104.205 69.840 104.395 ;
        RECT 71.695 104.225 71.865 104.415 ;
        RECT 73.535 104.205 73.705 104.395 ;
        RECT 74.915 104.225 75.085 104.415 ;
        RECT 76.570 104.205 76.740 104.395 ;
        RECT 78.590 104.255 78.710 104.365 ;
        RECT 79.055 104.225 79.225 104.415 ;
        RECT 80.435 104.205 80.605 104.395 ;
        RECT 82.275 104.225 82.445 104.415 ;
        RECT 84.390 104.225 84.560 104.415 ;
        RECT 88.070 104.205 88.240 104.395 ;
        RECT 88.255 104.225 88.425 104.415 ;
        RECT 90.090 104.255 90.210 104.365 ;
        RECT 90.560 104.225 90.730 104.415 ;
        RECT 91.935 104.205 92.105 104.395 ;
        RECT 94.235 104.225 94.405 104.415 ;
        RECT 95.155 104.205 95.325 104.395 ;
        RECT 95.615 104.225 95.785 104.415 ;
        RECT 101.620 104.395 101.730 104.415 ;
        RECT 101.620 104.225 101.790 104.395 ;
        RECT 102.330 104.225 102.500 104.415 ;
        RECT 102.790 104.205 102.960 104.395 ;
        RECT 106.195 104.225 106.365 104.415 ;
        RECT 106.650 104.255 106.770 104.365 ;
        RECT 107.115 104.205 107.285 104.395 ;
        RECT 108.030 104.255 108.150 104.365 ;
        RECT 108.770 104.225 108.940 104.415 ;
        RECT 112.635 104.225 112.805 104.415 ;
        RECT 114.480 104.225 114.650 104.415 ;
        RECT 114.750 104.205 114.920 104.395 ;
        RECT 118.155 104.225 118.325 104.415 ;
        RECT 118.615 104.205 118.785 104.395 ;
        RECT 121.190 104.205 121.360 104.395 ;
        RECT 123.675 104.225 123.845 104.415 ;
        RECT 125.055 104.205 125.225 104.395 ;
        RECT 126.435 104.205 126.605 104.415 ;
        RECT 129.195 104.225 129.365 104.415 ;
        RECT 132.415 104.225 132.585 104.415 ;
        RECT 132.870 104.255 132.990 104.365 ;
        RECT 133.795 104.205 133.965 104.415 ;
        RECT 135.630 104.255 135.750 104.365 ;
        RECT 136.370 104.205 136.540 104.395 ;
        RECT 139.315 104.225 139.485 104.415 ;
        RECT 139.775 104.225 139.945 104.415 ;
        RECT 141.610 104.255 141.730 104.365 ;
        RECT 142.075 104.225 142.245 104.415 ;
        RECT 142.995 104.205 143.165 104.395 ;
        RECT 143.450 104.255 143.570 104.365 ;
        RECT 143.915 104.205 144.085 104.415 ;
        RECT 146.675 104.205 146.845 104.415 ;
        RECT 32.455 103.495 36.125 104.175 ;
        RECT 32.455 103.295 33.405 103.495 ;
        RECT 36.675 103.295 39.675 104.205 ;
        RECT 40.295 103.295 41.645 104.205 ;
        RECT 41.655 103.395 43.025 104.205 ;
        RECT 43.045 103.335 43.475 104.120 ;
        RECT 43.495 103.395 49.005 104.205 ;
        RECT 49.015 103.395 54.525 104.205 ;
        RECT 54.535 103.395 58.205 104.205 ;
        RECT 58.675 103.525 61.425 104.205 ;
        RECT 61.435 103.525 68.745 104.205 ;
        RECT 58.675 103.295 59.605 103.525 ;
        RECT 64.950 103.305 65.860 103.525 ;
        RECT 67.395 103.295 68.745 103.525 ;
        RECT 68.805 103.335 69.235 104.120 ;
        RECT 69.255 103.525 73.155 104.205 ;
        RECT 73.395 103.525 76.145 104.205 ;
        RECT 69.255 103.295 70.185 103.525 ;
        RECT 75.215 103.295 76.145 103.525 ;
        RECT 76.155 103.525 80.055 104.205 ;
        RECT 80.295 103.525 87.605 104.205 ;
        RECT 76.155 103.295 77.085 103.525 ;
        RECT 83.810 103.305 84.720 103.525 ;
        RECT 86.255 103.295 87.605 103.525 ;
        RECT 87.655 103.525 91.555 104.205 ;
        RECT 91.795 103.525 94.545 104.205 ;
        RECT 87.655 103.295 88.585 103.525 ;
        RECT 93.615 103.295 94.545 103.525 ;
        RECT 94.565 103.335 94.995 104.120 ;
        RECT 95.015 103.525 102.325 104.205 ;
        RECT 98.530 103.305 99.440 103.525 ;
        RECT 100.975 103.295 102.325 103.525 ;
        RECT 102.375 103.525 106.275 104.205 ;
        RECT 106.975 103.525 114.285 104.205 ;
        RECT 102.375 103.295 103.305 103.525 ;
        RECT 110.490 103.305 111.400 103.525 ;
        RECT 112.935 103.295 114.285 103.525 ;
        RECT 114.335 103.525 118.235 104.205 ;
        RECT 114.335 103.295 115.265 103.525 ;
        RECT 118.475 103.395 120.305 104.205 ;
        RECT 120.325 103.335 120.755 104.120 ;
        RECT 120.775 103.525 124.675 104.205 ;
        RECT 120.775 103.295 121.705 103.525 ;
        RECT 124.915 103.395 126.285 104.205 ;
        RECT 126.295 103.525 133.605 104.205 ;
        RECT 133.655 103.525 135.485 104.205 ;
        RECT 135.955 103.525 139.855 104.205 ;
        RECT 129.810 103.305 130.720 103.525 ;
        RECT 132.255 103.295 133.605 103.525 ;
        RECT 135.955 103.295 136.885 103.525 ;
        RECT 140.095 103.295 143.305 104.205 ;
        RECT 143.775 103.525 145.605 104.205 ;
        RECT 144.260 103.295 145.605 103.525 ;
        RECT 145.615 103.395 146.985 104.205 ;
      LAYER nwell ;
        RECT 17.080 100.175 147.180 103.005 ;
      LAYER pwell ;
        RECT 17.275 98.975 18.645 99.785 ;
        RECT 18.655 98.975 21.405 99.785 ;
        RECT 24.930 99.655 25.840 99.875 ;
        RECT 27.375 99.655 28.725 99.885 ;
        RECT 21.415 98.975 28.725 99.655 ;
        RECT 28.795 98.975 30.145 99.885 ;
        RECT 30.165 99.060 30.595 99.845 ;
        RECT 31.615 98.975 35.065 99.885 ;
        RECT 35.295 98.975 38.745 99.885 ;
        RECT 38.975 98.975 42.425 99.885 ;
        RECT 42.655 98.975 46.105 99.885 ;
        RECT 48.075 99.655 49.005 99.885 ;
        RECT 46.255 98.975 49.005 99.655 ;
        RECT 49.015 98.975 54.525 99.785 ;
        RECT 54.535 98.975 55.905 99.785 ;
        RECT 55.925 99.060 56.355 99.845 ;
        RECT 56.375 98.975 57.745 99.785 ;
        RECT 61.270 99.655 62.180 99.875 ;
        RECT 63.715 99.655 65.065 99.885 ;
        RECT 68.630 99.655 69.540 99.875 ;
        RECT 71.075 99.655 72.425 99.885 ;
        RECT 72.960 99.655 74.305 99.885 ;
        RECT 77.830 99.655 78.740 99.875 ;
        RECT 80.275 99.655 81.625 99.885 ;
        RECT 57.755 98.975 65.065 99.655 ;
        RECT 65.115 98.975 72.425 99.655 ;
        RECT 72.475 98.975 74.305 99.655 ;
        RECT 74.315 98.975 81.625 99.655 ;
        RECT 81.685 99.060 82.115 99.845 ;
        RECT 82.135 98.975 85.345 99.885 ;
        RECT 85.355 98.975 87.185 99.785 ;
        RECT 90.710 99.655 91.620 99.875 ;
        RECT 93.155 99.655 94.505 99.885 ;
        RECT 87.195 98.975 94.505 99.655 ;
        RECT 94.555 98.975 95.925 99.755 ;
        RECT 99.450 99.655 100.360 99.875 ;
        RECT 101.895 99.655 103.245 99.885 ;
        RECT 95.935 98.975 103.245 99.655 ;
        RECT 103.295 98.975 106.950 99.885 ;
        RECT 107.445 99.060 107.875 99.845 ;
        RECT 111.410 99.655 112.320 99.875 ;
        RECT 113.855 99.655 115.205 99.885 ;
        RECT 118.770 99.655 119.680 99.875 ;
        RECT 121.215 99.655 122.565 99.885 ;
        RECT 126.130 99.655 127.040 99.875 ;
        RECT 128.575 99.655 129.925 99.885 ;
        RECT 107.895 98.975 115.205 99.655 ;
        RECT 115.255 98.975 122.565 99.655 ;
        RECT 122.615 98.975 129.925 99.655 ;
        RECT 129.975 99.655 130.905 99.885 ;
        RECT 129.975 98.975 132.725 99.655 ;
        RECT 133.205 99.060 133.635 99.845 ;
        RECT 137.630 99.655 138.540 99.875 ;
        RECT 140.075 99.655 141.425 99.885 ;
        RECT 134.115 98.975 141.425 99.655 ;
        RECT 141.475 99.655 142.405 99.885 ;
        RECT 141.475 98.975 145.375 99.655 ;
        RECT 145.615 98.975 146.985 99.785 ;
        RECT 17.415 98.765 17.585 98.975 ;
        RECT 18.795 98.925 18.965 98.975 ;
        RECT 18.790 98.815 18.965 98.925 ;
        RECT 18.795 98.785 18.965 98.815 ;
        RECT 21.555 98.785 21.725 98.975 ;
        RECT 26.155 98.765 26.325 98.955 ;
        RECT 26.890 98.765 27.060 98.955 ;
        RECT 29.830 98.785 30.000 98.975 ;
        RECT 31.675 98.955 31.845 98.975 ;
        RECT 30.765 98.810 30.925 98.930 ;
        RECT 31.675 98.785 31.850 98.955 ;
        RECT 31.680 98.765 31.850 98.785 ;
        RECT 34.895 98.765 35.065 98.955 ;
        RECT 35.355 98.785 35.525 98.975 ;
        RECT 39.035 98.785 39.205 98.975 ;
        RECT 17.275 97.955 18.645 98.765 ;
        RECT 19.155 98.085 26.465 98.765 ;
        RECT 26.475 98.085 30.375 98.765 ;
        RECT 19.155 97.855 20.505 98.085 ;
        RECT 22.040 97.865 22.950 98.085 ;
        RECT 26.475 97.855 27.405 98.085 ;
        RECT 31.535 97.855 34.455 98.765 ;
        RECT 34.835 97.855 38.285 98.765 ;
        RECT 38.435 98.735 39.380 98.765 ;
        RECT 40.870 98.735 41.040 98.955 ;
        RECT 41.340 98.765 41.510 98.955 ;
        RECT 42.715 98.925 42.885 98.975 ;
        RECT 42.710 98.815 42.885 98.925 ;
        RECT 42.715 98.785 42.885 98.815 ;
        RECT 43.635 98.765 43.805 98.955 ;
        RECT 46.395 98.765 46.565 98.975 ;
        RECT 49.155 98.785 49.325 98.975 ;
        RECT 51.915 98.765 52.085 98.955 ;
        RECT 54.675 98.785 54.845 98.975 ;
        RECT 56.515 98.785 56.685 98.975 ;
        RECT 57.895 98.785 58.065 98.975 ;
        RECT 58.355 98.765 58.525 98.955 ;
        RECT 58.815 98.765 58.985 98.955 ;
        RECT 60.655 98.765 60.825 98.955 ;
        RECT 65.255 98.785 65.425 98.975 ;
        RECT 68.025 98.810 68.185 98.920 ;
        RECT 69.670 98.765 69.840 98.955 ;
        RECT 72.615 98.785 72.785 98.975 ;
        RECT 73.535 98.765 73.705 98.955 ;
        RECT 74.455 98.785 74.625 98.975 ;
        RECT 76.755 98.765 76.925 98.955 ;
        RECT 82.275 98.765 82.445 98.975 ;
        RECT 83.655 98.765 83.825 98.955 ;
        RECT 85.495 98.785 85.665 98.975 ;
        RECT 87.335 98.785 87.505 98.975 ;
        RECT 91.020 98.765 91.190 98.955 ;
        RECT 95.430 98.765 95.600 98.955 ;
        RECT 95.605 98.785 95.775 98.975 ;
        RECT 96.075 98.785 96.245 98.975 ;
        RECT 99.295 98.765 99.465 98.955 ;
        RECT 102.055 98.765 102.225 98.955 ;
        RECT 103.440 98.785 103.610 98.975 ;
        RECT 104.815 98.765 104.985 98.955 ;
        RECT 107.110 98.815 107.230 98.925 ;
        RECT 107.575 98.765 107.745 98.955 ;
        RECT 108.035 98.785 108.205 98.975 ;
        RECT 111.255 98.765 111.425 98.955 ;
        RECT 112.635 98.765 112.805 98.955 ;
        RECT 115.395 98.925 115.565 98.975 ;
        RECT 115.390 98.815 115.565 98.925 ;
        RECT 115.395 98.785 115.565 98.815 ;
        RECT 116.130 98.765 116.300 98.955 ;
        RECT 119.990 98.815 120.110 98.925 ;
        RECT 120.915 98.765 121.085 98.955 ;
        RECT 122.755 98.785 122.925 98.975 ;
        RECT 123.675 98.765 123.845 98.955 ;
        RECT 131.310 98.765 131.480 98.955 ;
        RECT 132.415 98.785 132.585 98.975 ;
        RECT 132.870 98.815 132.990 98.925 ;
        RECT 133.790 98.815 133.910 98.925 ;
        RECT 134.255 98.785 134.425 98.975 ;
        RECT 136.085 98.765 136.255 98.955 ;
        RECT 136.555 98.765 136.725 98.955 ;
        RECT 141.890 98.785 142.060 98.975 ;
        RECT 143.915 98.765 144.085 98.955 ;
        RECT 146.675 98.765 146.845 98.975 ;
        RECT 38.435 98.055 41.185 98.735 ;
        RECT 38.435 97.855 39.380 98.055 ;
        RECT 41.195 97.855 42.545 98.765 ;
        RECT 43.045 97.895 43.475 98.680 ;
        RECT 43.495 97.855 46.245 98.765 ;
        RECT 46.255 97.955 51.765 98.765 ;
        RECT 51.775 97.955 57.285 98.765 ;
        RECT 57.295 97.985 58.665 98.765 ;
        RECT 58.675 97.955 60.505 98.765 ;
        RECT 60.515 98.085 67.825 98.765 ;
        RECT 64.030 97.865 64.940 98.085 ;
        RECT 66.475 97.855 67.825 98.085 ;
        RECT 68.805 97.895 69.235 98.680 ;
        RECT 69.255 98.085 73.155 98.765 ;
        RECT 69.255 97.855 70.185 98.085 ;
        RECT 73.395 97.855 76.605 98.765 ;
        RECT 76.615 97.955 82.125 98.765 ;
        RECT 82.135 97.955 83.505 98.765 ;
        RECT 83.515 98.085 90.825 98.765 ;
        RECT 87.030 97.865 87.940 98.085 ;
        RECT 89.475 97.855 90.825 98.085 ;
        RECT 90.875 97.855 94.530 98.765 ;
        RECT 94.565 97.895 94.995 98.680 ;
        RECT 95.015 98.085 98.915 98.765 ;
        RECT 99.155 98.085 101.905 98.765 ;
        RECT 95.015 97.855 95.945 98.085 ;
        RECT 100.975 97.855 101.905 98.085 ;
        RECT 101.915 97.955 104.665 98.765 ;
        RECT 104.675 98.085 107.425 98.765 ;
        RECT 106.495 97.855 107.425 98.085 ;
        RECT 107.435 97.955 111.105 98.765 ;
        RECT 111.115 97.955 112.485 98.765 ;
        RECT 112.495 98.085 115.245 98.765 ;
        RECT 114.315 97.855 115.245 98.085 ;
        RECT 115.715 98.085 119.615 98.765 ;
        RECT 115.715 97.855 116.645 98.085 ;
        RECT 120.325 97.895 120.755 98.680 ;
        RECT 120.775 97.955 123.525 98.765 ;
        RECT 123.535 98.085 130.845 98.765 ;
        RECT 127.050 97.865 127.960 98.085 ;
        RECT 129.495 97.855 130.845 98.085 ;
        RECT 130.895 98.085 134.795 98.765 ;
        RECT 130.895 97.855 131.825 98.085 ;
        RECT 135.035 97.985 136.405 98.765 ;
        RECT 136.415 98.085 143.725 98.765 ;
        RECT 143.775 98.085 145.605 98.765 ;
        RECT 139.930 97.865 140.840 98.085 ;
        RECT 142.375 97.855 143.725 98.085 ;
        RECT 144.260 97.855 145.605 98.085 ;
        RECT 145.615 97.955 146.985 98.765 ;
      LAYER nwell ;
        RECT 17.080 94.735 147.180 97.565 ;
      LAYER pwell ;
        RECT 17.275 93.535 18.645 94.345 ;
        RECT 18.655 93.535 20.025 94.315 ;
        RECT 20.035 93.535 21.405 94.315 ;
        RECT 21.875 94.215 23.220 94.445 ;
        RECT 21.875 93.535 23.705 94.215 ;
        RECT 23.715 93.535 25.085 94.315 ;
        RECT 25.095 93.535 26.465 94.315 ;
        RECT 26.475 93.535 28.305 94.345 ;
        RECT 28.800 94.215 30.145 94.445 ;
        RECT 28.315 93.535 30.145 94.215 ;
        RECT 30.165 93.620 30.595 94.405 ;
        RECT 30.615 93.535 31.985 94.315 ;
        RECT 32.075 93.535 35.075 94.445 ;
        RECT 35.215 93.535 36.585 94.315 ;
        RECT 36.595 93.535 37.965 94.345 ;
        RECT 37.975 93.535 39.345 94.315 ;
        RECT 39.355 93.535 41.185 94.345 ;
        RECT 41.195 93.535 42.565 94.315 ;
        RECT 43.045 93.620 43.475 94.405 ;
        RECT 44.415 93.535 45.785 94.315 ;
        RECT 45.795 93.535 47.625 94.345 ;
        RECT 47.635 93.535 49.005 94.315 ;
        RECT 49.015 93.535 50.845 94.345 ;
        RECT 50.855 93.535 52.225 94.315 ;
        RECT 52.235 93.535 54.065 94.345 ;
        RECT 54.075 93.535 55.445 94.315 ;
        RECT 55.925 93.620 56.355 94.405 ;
        RECT 56.375 94.215 57.720 94.445 ;
        RECT 58.215 94.215 59.560 94.445 ;
        RECT 60.055 94.215 61.400 94.445 ;
        RECT 61.895 94.215 62.825 94.445 ;
        RECT 67.395 94.215 68.325 94.445 ;
        RECT 56.375 93.535 58.205 94.215 ;
        RECT 58.215 93.535 60.045 94.215 ;
        RECT 60.055 93.535 61.885 94.215 ;
        RECT 61.895 93.535 64.645 94.215 ;
        RECT 65.575 93.535 68.325 94.215 ;
        RECT 68.805 93.620 69.235 94.405 ;
        RECT 69.255 94.215 70.185 94.445 ;
        RECT 73.880 94.215 75.225 94.445 ;
        RECT 69.255 93.535 73.155 94.215 ;
        RECT 73.395 93.535 75.225 94.215 ;
        RECT 76.155 94.215 77.500 94.445 ;
        RECT 78.480 94.215 79.825 94.445 ;
        RECT 80.320 94.215 81.665 94.445 ;
        RECT 76.155 93.535 77.985 94.215 ;
        RECT 77.995 93.535 79.825 94.215 ;
        RECT 79.835 93.535 81.665 94.215 ;
        RECT 81.685 93.620 82.115 94.405 ;
        RECT 82.135 93.535 83.505 94.345 ;
        RECT 85.335 94.215 86.265 94.445 ;
        RECT 89.015 94.215 89.945 94.445 ;
        RECT 83.515 93.535 86.265 94.215 ;
        RECT 87.195 93.535 89.945 94.215 ;
        RECT 89.955 94.215 91.300 94.445 ;
        RECT 92.280 94.215 93.625 94.445 ;
        RECT 89.955 93.535 91.785 94.215 ;
        RECT 91.795 93.535 93.625 94.215 ;
        RECT 94.565 93.620 94.995 94.405 ;
        RECT 95.500 94.215 96.845 94.445 ;
        RECT 97.340 94.215 98.685 94.445 ;
        RECT 95.015 93.535 96.845 94.215 ;
        RECT 96.855 93.535 98.685 94.215 ;
        RECT 99.155 94.215 100.500 94.445 ;
        RECT 99.155 93.535 100.985 94.215 ;
        RECT 100.995 93.535 102.365 94.345 ;
        RECT 102.375 94.215 103.720 94.445 ;
        RECT 102.375 93.535 104.205 94.215 ;
        RECT 104.215 93.535 105.585 94.345 ;
        RECT 105.595 94.215 106.940 94.445 ;
        RECT 105.595 93.535 107.425 94.215 ;
        RECT 107.445 93.620 107.875 94.405 ;
        RECT 108.815 94.215 110.160 94.445 ;
        RECT 108.815 93.535 110.645 94.215 ;
        RECT 110.655 93.535 112.025 94.345 ;
        RECT 112.035 94.215 113.380 94.445 ;
        RECT 115.695 94.215 116.625 94.445 ;
        RECT 112.035 93.535 113.865 94.215 ;
        RECT 113.875 93.535 116.625 94.215 ;
        RECT 117.095 93.535 120.305 94.445 ;
        RECT 120.325 93.620 120.755 94.405 ;
        RECT 121.260 94.215 122.605 94.445 ;
        RECT 123.100 94.215 124.445 94.445 ;
        RECT 120.775 93.535 122.605 94.215 ;
        RECT 122.615 93.535 124.445 94.215 ;
        RECT 124.455 94.215 125.800 94.445 ;
        RECT 129.495 94.215 130.425 94.445 ;
        RECT 130.920 94.215 132.265 94.445 ;
        RECT 124.455 93.535 126.285 94.215 ;
        RECT 126.525 93.535 130.425 94.215 ;
        RECT 130.435 93.535 132.265 94.215 ;
        RECT 133.205 93.620 133.635 94.405 ;
        RECT 133.670 93.535 137.325 94.445 ;
        RECT 139.155 94.215 140.085 94.445 ;
        RECT 140.580 94.215 141.925 94.445 ;
        RECT 142.420 94.215 143.765 94.445 ;
        RECT 144.260 94.215 145.605 94.445 ;
        RECT 137.335 93.535 140.085 94.215 ;
        RECT 140.095 93.535 141.925 94.215 ;
        RECT 141.935 93.535 143.765 94.215 ;
        RECT 143.775 93.535 145.605 94.215 ;
        RECT 145.615 93.535 146.985 94.345 ;
        RECT 17.415 93.345 17.585 93.535 ;
        RECT 18.805 93.345 18.975 93.535 ;
        RECT 20.175 93.345 20.345 93.535 ;
        RECT 21.550 93.375 21.670 93.485 ;
        RECT 23.395 93.345 23.565 93.535 ;
        RECT 23.865 93.345 24.035 93.535 ;
        RECT 25.245 93.345 25.415 93.535 ;
        RECT 26.615 93.345 26.785 93.535 ;
        RECT 28.455 93.345 28.625 93.535 ;
        RECT 30.765 93.345 30.935 93.535 ;
        RECT 32.135 93.345 32.305 93.535 ;
        RECT 35.355 93.345 35.525 93.535 ;
        RECT 36.735 93.345 36.905 93.535 ;
        RECT 38.115 93.345 38.285 93.535 ;
        RECT 39.495 93.345 39.665 93.535 ;
        RECT 42.245 93.345 42.415 93.535 ;
        RECT 42.710 93.375 42.830 93.485 ;
        RECT 43.645 93.380 43.805 93.490 ;
        RECT 45.465 93.345 45.635 93.535 ;
        RECT 45.935 93.345 46.105 93.535 ;
        RECT 48.685 93.345 48.855 93.535 ;
        RECT 49.155 93.345 49.325 93.535 ;
        RECT 51.915 93.345 52.085 93.535 ;
        RECT 52.375 93.345 52.545 93.535 ;
        RECT 55.135 93.345 55.305 93.535 ;
        RECT 55.590 93.375 55.710 93.485 ;
        RECT 57.895 93.345 58.065 93.535 ;
        RECT 59.735 93.345 59.905 93.535 ;
        RECT 61.575 93.345 61.745 93.535 ;
        RECT 64.335 93.345 64.505 93.535 ;
        RECT 64.805 93.380 64.965 93.490 ;
        RECT 65.715 93.345 65.885 93.535 ;
        RECT 68.470 93.375 68.590 93.485 ;
        RECT 69.670 93.345 69.840 93.535 ;
        RECT 73.535 93.345 73.705 93.535 ;
        RECT 75.385 93.380 75.545 93.490 ;
        RECT 77.675 93.345 77.845 93.535 ;
        RECT 78.135 93.345 78.305 93.535 ;
        RECT 79.975 93.345 80.145 93.535 ;
        RECT 82.275 93.345 82.445 93.535 ;
        RECT 83.655 93.345 83.825 93.535 ;
        RECT 86.425 93.380 86.585 93.490 ;
        RECT 87.335 93.345 87.505 93.535 ;
        RECT 91.475 93.345 91.645 93.535 ;
        RECT 91.935 93.345 92.105 93.535 ;
        RECT 93.785 93.380 93.945 93.490 ;
        RECT 95.155 93.345 95.325 93.535 ;
        RECT 96.995 93.345 97.165 93.535 ;
        RECT 98.830 93.375 98.950 93.485 ;
        RECT 100.675 93.345 100.845 93.535 ;
        RECT 101.135 93.345 101.305 93.535 ;
        RECT 103.895 93.345 104.065 93.535 ;
        RECT 104.355 93.345 104.525 93.535 ;
        RECT 107.115 93.345 107.285 93.535 ;
        RECT 108.045 93.380 108.205 93.490 ;
        RECT 110.335 93.345 110.505 93.535 ;
        RECT 110.795 93.345 110.965 93.535 ;
        RECT 113.555 93.345 113.725 93.535 ;
        RECT 114.015 93.345 114.185 93.535 ;
        RECT 116.770 93.375 116.890 93.485 ;
        RECT 119.995 93.345 120.165 93.535 ;
        RECT 120.915 93.345 121.085 93.535 ;
        RECT 122.755 93.345 122.925 93.535 ;
        RECT 125.975 93.345 126.145 93.535 ;
        RECT 129.840 93.345 130.010 93.535 ;
        RECT 130.575 93.345 130.745 93.535 ;
        RECT 132.425 93.380 132.585 93.490 ;
        RECT 137.010 93.345 137.180 93.535 ;
        RECT 137.475 93.345 137.645 93.535 ;
        RECT 140.235 93.345 140.405 93.535 ;
        RECT 142.075 93.345 142.245 93.535 ;
        RECT 143.915 93.345 144.085 93.535 ;
        RECT 146.675 93.345 146.845 93.535 ;
      LAYER nwell ;
        RECT 54.490 67.690 67.660 75.530 ;
      LAYER pwell ;
        RECT 54.500 63.190 67.670 66.980 ;
        RECT 54.500 55.700 68.350 62.920 ;
        RECT 72.890 58.540 74.900 76.510 ;
      LAYER nwell ;
        RECT 74.900 65.670 87.150 75.860 ;
        RECT 89.880 65.650 102.130 75.840 ;
        RECT 104.890 65.650 117.140 75.840 ;
        RECT 119.900 65.650 132.150 75.840 ;
        RECT 134.890 65.650 147.140 75.840 ;
      LAYER pwell ;
        RECT 84.700 64.440 86.810 64.450 ;
        RECT 54.500 49.710 65.390 55.700 ;
      LAYER nwell ;
        RECT 54.540 37.650 66.790 47.840 ;
      LAYER pwell ;
        RECT 64.340 36.420 66.450 36.430 ;
        RECT 54.550 33.640 66.450 36.420 ;
        RECT 54.550 31.680 64.370 33.640 ;
        RECT 54.550 30.520 64.770 31.680 ;
      LAYER nwell ;
        RECT 66.450 31.530 68.560 36.370 ;
      LAYER pwell ;
        RECT 54.550 30.320 64.370 30.520 ;
      LAYER nwell ;
        RECT 61.320 22.420 66.970 28.610 ;
      LAYER pwell ;
        RECT 71.410 28.590 74.900 58.540 ;
        RECT 74.910 61.660 86.810 64.440 ;
        RECT 99.680 64.420 101.790 64.430 ;
        RECT 114.690 64.420 116.800 64.430 ;
        RECT 129.700 64.420 131.810 64.430 ;
        RECT 144.690 64.420 146.800 64.430 ;
        RECT 74.910 59.700 84.730 61.660 ;
        RECT 74.910 58.540 85.130 59.700 ;
      LAYER nwell ;
        RECT 86.810 59.550 88.920 64.390 ;
      LAYER pwell ;
        RECT 89.890 61.640 101.790 64.420 ;
        RECT 89.890 59.680 99.710 61.640 ;
        RECT 74.910 58.340 84.730 58.540 ;
        RECT 89.890 58.520 100.110 59.680 ;
      LAYER nwell ;
        RECT 101.790 59.530 103.900 64.370 ;
      LAYER pwell ;
        RECT 104.900 61.640 116.800 64.420 ;
        RECT 104.900 59.680 114.720 61.640 ;
        RECT 104.900 58.520 115.120 59.680 ;
      LAYER nwell ;
        RECT 116.800 59.530 118.910 64.370 ;
      LAYER pwell ;
        RECT 119.910 61.640 131.810 64.420 ;
        RECT 119.910 59.680 129.730 61.640 ;
        RECT 119.910 58.520 130.130 59.680 ;
      LAYER nwell ;
        RECT 131.810 59.530 133.920 64.370 ;
      LAYER pwell ;
        RECT 134.900 61.640 146.800 64.420 ;
        RECT 134.900 59.680 144.720 61.640 ;
        RECT 134.900 58.520 145.120 59.680 ;
      LAYER nwell ;
        RECT 146.800 59.530 148.910 64.370 ;
      LAYER pwell ;
        RECT 89.890 58.320 99.710 58.520 ;
        RECT 104.900 58.320 114.720 58.520 ;
        RECT 119.910 58.320 129.730 58.520 ;
        RECT 134.900 58.320 144.720 58.520 ;
      LAYER nwell ;
        RECT 74.900 46.660 87.150 56.850 ;
        RECT 89.880 46.650 102.130 56.840 ;
        RECT 104.920 46.650 117.170 56.840 ;
        RECT 119.900 46.650 132.150 56.840 ;
        RECT 134.910 46.680 147.160 56.870 ;
      LAYER pwell ;
        RECT 144.710 45.450 146.820 45.460 ;
        RECT 84.700 45.430 86.810 45.440 ;
        RECT 74.910 42.650 86.810 45.430 ;
        RECT 99.680 45.420 101.790 45.430 ;
        RECT 114.720 45.420 116.830 45.430 ;
        RECT 129.700 45.420 131.810 45.430 ;
        RECT 74.910 40.690 84.730 42.650 ;
        RECT 74.910 39.530 85.130 40.690 ;
      LAYER nwell ;
        RECT 86.810 40.540 88.920 45.380 ;
      LAYER pwell ;
        RECT 89.890 42.640 101.790 45.420 ;
        RECT 89.890 40.680 99.710 42.640 ;
        RECT 74.910 39.330 84.730 39.530 ;
        RECT 89.890 39.520 100.110 40.680 ;
      LAYER nwell ;
        RECT 101.790 40.530 103.900 45.370 ;
      LAYER pwell ;
        RECT 104.930 42.640 116.830 45.420 ;
        RECT 104.930 40.680 114.750 42.640 ;
        RECT 104.930 39.520 115.150 40.680 ;
      LAYER nwell ;
        RECT 116.830 40.530 118.940 45.370 ;
      LAYER pwell ;
        RECT 119.910 42.640 131.810 45.420 ;
        RECT 119.910 40.680 129.730 42.640 ;
        RECT 119.910 39.520 130.130 40.680 ;
      LAYER nwell ;
        RECT 131.810 40.530 133.920 45.370 ;
      LAYER pwell ;
        RECT 134.920 42.670 146.820 45.450 ;
        RECT 134.920 40.710 144.740 42.670 ;
        RECT 134.920 39.550 145.140 40.710 ;
      LAYER nwell ;
        RECT 146.820 40.560 148.930 45.400 ;
      LAYER pwell ;
        RECT 89.890 39.320 99.710 39.520 ;
        RECT 104.930 39.320 114.750 39.520 ;
        RECT 119.910 39.320 129.730 39.520 ;
        RECT 134.920 39.350 144.740 39.550 ;
        RECT 69.930 22.070 74.900 28.590 ;
      LAYER nwell ;
        RECT 74.940 27.650 87.190 37.840 ;
        RECT 89.880 27.650 102.130 37.840 ;
        RECT 104.890 27.650 117.140 37.840 ;
        RECT 119.930 27.650 132.180 37.840 ;
        RECT 134.890 27.650 147.140 37.840 ;
      LAYER pwell ;
        RECT 84.740 26.420 86.850 26.430 ;
        RECT 99.680 26.420 101.790 26.430 ;
        RECT 114.690 26.420 116.800 26.430 ;
        RECT 129.730 26.420 131.840 26.430 ;
        RECT 144.690 26.420 146.800 26.430 ;
        RECT 74.950 23.640 86.850 26.420 ;
        RECT 61.310 18.960 66.960 22.060 ;
        RECT 74.950 21.680 84.770 23.640 ;
        RECT 74.950 20.520 85.170 21.680 ;
      LAYER nwell ;
        RECT 86.850 21.530 88.960 26.370 ;
      LAYER pwell ;
        RECT 89.890 23.640 101.790 26.420 ;
        RECT 89.890 21.680 99.710 23.640 ;
        RECT 89.890 20.520 100.110 21.680 ;
      LAYER nwell ;
        RECT 101.790 21.530 103.900 26.370 ;
      LAYER pwell ;
        RECT 104.900 23.640 116.800 26.420 ;
        RECT 104.900 21.680 114.720 23.640 ;
        RECT 104.900 20.520 115.120 21.680 ;
      LAYER nwell ;
        RECT 116.800 21.530 118.910 26.370 ;
      LAYER pwell ;
        RECT 119.940 23.640 131.840 26.420 ;
        RECT 119.940 21.680 129.760 23.640 ;
        RECT 119.940 20.520 130.160 21.680 ;
      LAYER nwell ;
        RECT 131.840 21.530 133.950 26.370 ;
      LAYER pwell ;
        RECT 134.900 23.640 146.800 26.420 ;
        RECT 134.900 21.680 144.720 23.640 ;
        RECT 134.900 20.520 145.120 21.680 ;
      LAYER nwell ;
        RECT 146.800 21.530 148.910 26.370 ;
      LAYER pwell ;
        RECT 74.950 20.320 84.770 20.520 ;
        RECT 89.890 20.320 99.710 20.520 ;
        RECT 104.900 20.320 114.720 20.520 ;
        RECT 119.940 20.320 129.760 20.520 ;
        RECT 134.900 20.320 144.720 20.520 ;
      LAYER li1 ;
        RECT 33.300 224.810 33.870 225.380 ;
        RECT 33.430 221.355 33.730 224.810 ;
        RECT 17.270 221.185 146.990 221.355 ;
        RECT 17.355 220.095 18.565 221.185 ;
        RECT 18.735 220.750 24.080 221.185 ;
        RECT 24.255 220.750 29.600 221.185 ;
        RECT 17.355 219.385 17.875 219.925 ;
        RECT 18.045 219.555 18.565 220.095 ;
        RECT 17.355 218.635 18.565 219.385 ;
        RECT 20.320 219.180 20.660 220.010 ;
        RECT 22.140 219.500 22.490 220.750 ;
        RECT 25.840 219.180 26.180 220.010 ;
        RECT 27.660 219.500 28.010 220.750 ;
        RECT 30.235 220.020 30.525 221.185 ;
        RECT 30.695 220.750 36.040 221.185 ;
        RECT 36.215 220.750 41.560 221.185 ;
        RECT 18.735 218.635 24.080 219.180 ;
        RECT 24.255 218.635 29.600 219.180 ;
        RECT 30.235 218.635 30.525 219.360 ;
        RECT 32.280 219.180 32.620 220.010 ;
        RECT 34.100 219.500 34.450 220.750 ;
        RECT 37.800 219.180 38.140 220.010 ;
        RECT 39.620 219.500 39.970 220.750 ;
        RECT 41.735 220.095 42.945 221.185 ;
        RECT 41.735 219.385 42.255 219.925 ;
        RECT 42.425 219.555 42.945 220.095 ;
        RECT 43.115 220.020 43.405 221.185 ;
        RECT 43.575 220.750 48.920 221.185 ;
        RECT 49.095 220.750 54.440 221.185 ;
        RECT 30.695 218.635 36.040 219.180 ;
        RECT 36.215 218.635 41.560 219.180 ;
        RECT 41.735 218.635 42.945 219.385 ;
        RECT 43.115 218.635 43.405 219.360 ;
        RECT 45.160 219.180 45.500 220.010 ;
        RECT 46.980 219.500 47.330 220.750 ;
        RECT 50.680 219.180 51.020 220.010 ;
        RECT 52.500 219.500 52.850 220.750 ;
        RECT 54.615 220.095 55.825 221.185 ;
        RECT 54.615 219.385 55.135 219.925 ;
        RECT 55.305 219.555 55.825 220.095 ;
        RECT 55.995 220.020 56.285 221.185 ;
        RECT 56.455 220.095 59.965 221.185 ;
        RECT 56.455 219.405 58.105 219.925 ;
        RECT 58.275 219.575 59.965 220.095 ;
        RECT 60.605 220.205 60.935 221.015 ;
        RECT 61.105 220.385 61.345 221.185 ;
        RECT 60.605 220.035 61.320 220.205 ;
        RECT 60.600 219.625 60.980 219.865 ;
        RECT 61.150 219.795 61.320 220.035 ;
        RECT 61.525 220.165 61.695 221.015 ;
        RECT 61.865 220.385 62.195 221.185 ;
        RECT 62.365 220.165 62.535 221.015 ;
        RECT 61.525 219.995 62.535 220.165 ;
        RECT 62.705 220.035 63.035 221.185 ;
        RECT 63.355 220.750 68.700 221.185 ;
        RECT 61.150 219.625 61.650 219.795 ;
        RECT 61.150 219.455 61.320 219.625 ;
        RECT 62.040 219.485 62.535 219.995 ;
        RECT 62.035 219.455 62.535 219.485 ;
        RECT 43.575 218.635 48.920 219.180 ;
        RECT 49.095 218.635 54.440 219.180 ;
        RECT 54.615 218.635 55.825 219.385 ;
        RECT 55.995 218.635 56.285 219.360 ;
        RECT 56.455 218.635 59.965 219.405 ;
        RECT 60.685 219.285 61.320 219.455 ;
        RECT 61.525 219.285 62.535 219.455 ;
        RECT 60.685 218.805 60.855 219.285 ;
        RECT 61.035 218.635 61.275 219.115 ;
        RECT 61.525 218.805 61.695 219.285 ;
        RECT 61.865 218.635 62.195 219.115 ;
        RECT 62.365 218.805 62.535 219.285 ;
        RECT 62.705 218.635 63.035 219.435 ;
        RECT 64.940 219.180 65.280 220.010 ;
        RECT 66.760 219.500 67.110 220.750 ;
        RECT 68.875 220.020 69.165 221.185 ;
        RECT 69.335 220.750 74.680 221.185 ;
        RECT 63.355 218.635 68.700 219.180 ;
        RECT 68.875 218.635 69.165 219.360 ;
        RECT 70.920 219.180 71.260 220.010 ;
        RECT 72.740 219.500 73.090 220.750 ;
        RECT 74.855 220.095 78.365 221.185 ;
        RECT 78.535 220.095 79.745 221.185 ;
        RECT 74.855 219.405 76.505 219.925 ;
        RECT 76.675 219.575 78.365 220.095 ;
        RECT 69.335 218.635 74.680 219.180 ;
        RECT 74.855 218.635 78.365 219.405 ;
        RECT 78.535 219.385 79.055 219.925 ;
        RECT 79.225 219.555 79.745 220.095 ;
        RECT 79.920 220.035 80.180 221.185 ;
        RECT 80.355 220.110 80.610 221.015 ;
        RECT 80.780 220.425 81.110 221.185 ;
        RECT 81.325 220.255 81.495 221.015 ;
        RECT 78.535 218.635 79.745 219.385 ;
        RECT 79.920 218.635 80.180 219.475 ;
        RECT 80.355 219.380 80.525 220.110 ;
        RECT 80.780 220.085 81.495 220.255 ;
        RECT 80.780 219.875 80.950 220.085 ;
        RECT 81.755 220.020 82.045 221.185 ;
        RECT 83.215 220.255 83.395 221.015 ;
        RECT 83.575 220.425 83.905 221.185 ;
        RECT 83.215 220.085 83.890 220.255 ;
        RECT 84.075 220.110 84.345 221.015 ;
        RECT 83.720 219.940 83.890 220.085 ;
        RECT 80.695 219.545 80.950 219.875 ;
        RECT 80.355 218.805 80.610 219.380 ;
        RECT 80.780 219.355 80.950 219.545 ;
        RECT 81.230 219.535 81.585 219.905 ;
        RECT 83.155 219.535 83.495 219.905 ;
        RECT 83.720 219.610 83.995 219.940 ;
        RECT 80.780 219.185 81.495 219.355 ;
        RECT 80.780 218.635 81.110 219.015 ;
        RECT 81.325 218.805 81.495 219.185 ;
        RECT 81.755 218.635 82.045 219.360 ;
        RECT 83.720 219.355 83.890 219.610 ;
        RECT 83.225 219.185 83.890 219.355 ;
        RECT 84.165 219.310 84.345 220.110 ;
        RECT 83.225 218.805 83.395 219.185 ;
        RECT 83.575 218.635 83.905 219.015 ;
        RECT 84.085 218.805 84.345 219.310 ;
        RECT 85.435 220.465 85.895 221.015 ;
        RECT 86.085 220.465 86.415 221.185 ;
        RECT 85.435 219.095 85.685 220.465 ;
        RECT 86.615 220.295 86.915 220.845 ;
        RECT 87.085 220.515 87.365 221.185 ;
        RECT 85.975 220.125 86.915 220.295 ;
        RECT 87.815 220.255 87.995 221.015 ;
        RECT 88.175 220.425 88.505 221.185 ;
        RECT 85.975 219.875 86.145 220.125 ;
        RECT 87.285 219.875 87.550 220.235 ;
        RECT 87.815 220.085 88.490 220.255 ;
        RECT 88.675 220.110 88.945 221.015 ;
        RECT 88.320 219.940 88.490 220.085 ;
        RECT 85.855 219.545 86.145 219.875 ;
        RECT 86.315 219.625 86.655 219.875 ;
        RECT 86.875 219.625 87.550 219.875 ;
        RECT 85.975 219.455 86.145 219.545 ;
        RECT 87.755 219.535 88.095 219.905 ;
        RECT 88.320 219.610 88.595 219.940 ;
        RECT 85.975 219.265 87.365 219.455 ;
        RECT 88.320 219.355 88.490 219.610 ;
        RECT 85.435 218.805 85.995 219.095 ;
        RECT 86.165 218.635 86.415 219.095 ;
        RECT 87.035 218.905 87.365 219.265 ;
        RECT 87.825 219.185 88.490 219.355 ;
        RECT 88.765 219.310 88.945 220.110 ;
        RECT 89.115 220.095 90.325 221.185 ;
        RECT 87.825 218.805 87.995 219.185 ;
        RECT 88.175 218.635 88.505 219.015 ;
        RECT 88.685 218.805 88.945 219.310 ;
        RECT 89.115 219.385 89.635 219.925 ;
        RECT 89.805 219.555 90.325 220.095 ;
        RECT 90.535 220.045 90.765 221.185 ;
        RECT 90.935 220.035 91.265 221.015 ;
        RECT 91.435 220.045 91.645 221.185 ;
        RECT 91.875 220.095 94.465 221.185 ;
        RECT 90.515 219.625 90.845 219.875 ;
        RECT 89.115 218.635 90.325 219.385 ;
        RECT 90.535 218.635 90.765 219.455 ;
        RECT 91.015 219.435 91.265 220.035 ;
        RECT 90.935 218.805 91.265 219.435 ;
        RECT 91.435 218.635 91.645 219.455 ;
        RECT 91.875 219.405 93.085 219.925 ;
        RECT 93.255 219.575 94.465 220.095 ;
        RECT 94.635 220.020 94.925 221.185 ;
        RECT 96.020 220.035 96.280 221.185 ;
        RECT 96.455 220.110 96.710 221.015 ;
        RECT 96.880 220.425 97.210 221.185 ;
        RECT 97.425 220.255 97.595 221.015 ;
        RECT 97.855 220.750 103.200 221.185 ;
        RECT 91.875 218.635 94.465 219.405 ;
        RECT 94.635 218.635 94.925 219.360 ;
        RECT 96.020 218.635 96.280 219.475 ;
        RECT 96.455 219.380 96.625 220.110 ;
        RECT 96.880 220.085 97.595 220.255 ;
        RECT 96.880 219.875 97.050 220.085 ;
        RECT 96.795 219.545 97.050 219.875 ;
        RECT 96.455 218.805 96.710 219.380 ;
        RECT 96.880 219.355 97.050 219.545 ;
        RECT 97.330 219.535 97.685 219.905 ;
        RECT 96.880 219.185 97.595 219.355 ;
        RECT 96.880 218.635 97.210 219.015 ;
        RECT 97.425 218.805 97.595 219.185 ;
        RECT 99.440 219.180 99.780 220.010 ;
        RECT 101.260 219.500 101.610 220.750 ;
        RECT 103.375 220.095 106.885 221.185 ;
        RECT 103.375 219.405 105.025 219.925 ;
        RECT 105.195 219.575 106.885 220.095 ;
        RECT 107.515 220.020 107.805 221.185 ;
        RECT 107.975 220.750 113.320 221.185 ;
        RECT 113.495 220.750 118.840 221.185 ;
        RECT 97.855 218.635 103.200 219.180 ;
        RECT 103.375 218.635 106.885 219.405 ;
        RECT 107.515 218.635 107.805 219.360 ;
        RECT 109.560 219.180 109.900 220.010 ;
        RECT 111.380 219.500 111.730 220.750 ;
        RECT 115.080 219.180 115.420 220.010 ;
        RECT 116.900 219.500 117.250 220.750 ;
        RECT 119.015 220.095 120.225 221.185 ;
        RECT 119.015 219.385 119.535 219.925 ;
        RECT 119.705 219.555 120.225 220.095 ;
        RECT 120.395 220.020 120.685 221.185 ;
        RECT 120.855 220.750 126.200 221.185 ;
        RECT 126.375 220.750 131.720 221.185 ;
        RECT 107.975 218.635 113.320 219.180 ;
        RECT 113.495 218.635 118.840 219.180 ;
        RECT 119.015 218.635 120.225 219.385 ;
        RECT 120.395 218.635 120.685 219.360 ;
        RECT 122.440 219.180 122.780 220.010 ;
        RECT 124.260 219.500 124.610 220.750 ;
        RECT 127.960 219.180 128.300 220.010 ;
        RECT 129.780 219.500 130.130 220.750 ;
        RECT 131.895 220.095 133.105 221.185 ;
        RECT 131.895 219.385 132.415 219.925 ;
        RECT 132.585 219.555 133.105 220.095 ;
        RECT 133.275 220.020 133.565 221.185 ;
        RECT 133.735 220.750 139.080 221.185 ;
        RECT 139.255 220.750 144.600 221.185 ;
        RECT 120.855 218.635 126.200 219.180 ;
        RECT 126.375 218.635 131.720 219.180 ;
        RECT 131.895 218.635 133.105 219.385 ;
        RECT 133.275 218.635 133.565 219.360 ;
        RECT 135.320 219.180 135.660 220.010 ;
        RECT 137.140 219.500 137.490 220.750 ;
        RECT 140.840 219.180 141.180 220.010 ;
        RECT 142.660 219.500 143.010 220.750 ;
        RECT 145.695 220.095 146.905 221.185 ;
        RECT 145.695 219.555 146.215 220.095 ;
        RECT 146.385 219.385 146.905 219.925 ;
        RECT 133.735 218.635 139.080 219.180 ;
        RECT 139.255 218.635 144.600 219.180 ;
        RECT 145.695 218.635 146.905 219.385 ;
        RECT 17.270 218.465 146.990 218.635 ;
        RECT 17.355 217.715 18.565 218.465 ;
        RECT 18.735 217.920 24.080 218.465 ;
        RECT 24.255 217.920 29.600 218.465 ;
        RECT 29.775 217.920 35.120 218.465 ;
        RECT 35.295 217.920 40.640 218.465 ;
        RECT 17.355 217.175 17.875 217.715 ;
        RECT 18.045 217.005 18.565 217.545 ;
        RECT 20.320 217.090 20.660 217.920 ;
        RECT 17.355 215.915 18.565 217.005 ;
        RECT 22.140 216.350 22.490 217.600 ;
        RECT 25.840 217.090 26.180 217.920 ;
        RECT 27.660 216.350 28.010 217.600 ;
        RECT 31.360 217.090 31.700 217.920 ;
        RECT 33.180 216.350 33.530 217.600 ;
        RECT 36.880 217.090 37.220 217.920 ;
        RECT 40.815 217.695 42.485 218.465 ;
        RECT 43.115 217.740 43.405 218.465 ;
        RECT 43.575 217.920 48.920 218.465 ;
        RECT 38.700 216.350 39.050 217.600 ;
        RECT 40.815 217.175 41.565 217.695 ;
        RECT 41.735 217.005 42.485 217.525 ;
        RECT 45.160 217.090 45.500 217.920 ;
        RECT 49.095 217.695 51.685 218.465 ;
        RECT 52.385 218.065 52.715 218.465 ;
        RECT 52.885 217.895 53.055 218.165 ;
        RECT 53.225 218.065 53.555 218.465 ;
        RECT 53.725 217.895 53.980 218.165 ;
        RECT 54.225 218.065 54.555 218.465 ;
        RECT 54.725 217.895 54.895 218.165 ;
        RECT 55.065 218.065 55.395 218.465 ;
        RECT 55.565 217.895 55.820 218.165 ;
        RECT 18.735 215.915 24.080 216.350 ;
        RECT 24.255 215.915 29.600 216.350 ;
        RECT 29.775 215.915 35.120 216.350 ;
        RECT 35.295 215.915 40.640 216.350 ;
        RECT 40.815 215.915 42.485 217.005 ;
        RECT 43.115 215.915 43.405 217.080 ;
        RECT 46.980 216.350 47.330 217.600 ;
        RECT 49.095 217.175 50.305 217.695 ;
        RECT 50.475 217.005 51.685 217.525 ;
        RECT 43.575 215.915 48.920 216.350 ;
        RECT 49.095 215.915 51.685 217.005 ;
        RECT 52.315 216.885 52.585 217.895 ;
        RECT 52.755 217.725 53.980 217.895 ;
        RECT 52.755 217.055 52.925 217.725 ;
        RECT 53.095 217.225 53.475 217.555 ;
        RECT 53.645 217.225 53.980 217.555 ;
        RECT 52.755 216.885 53.070 217.055 ;
        RECT 52.320 215.915 52.635 216.715 ;
        RECT 52.900 216.270 53.070 216.885 ;
        RECT 53.240 216.545 53.475 217.225 ;
        RECT 53.645 216.270 53.980 217.055 ;
        RECT 54.155 216.885 54.425 217.895 ;
        RECT 54.595 217.725 55.820 217.895 ;
        RECT 57.030 217.835 57.315 218.295 ;
        RECT 57.485 218.005 57.755 218.465 ;
        RECT 54.595 217.055 54.765 217.725 ;
        RECT 57.030 217.665 57.985 217.835 ;
        RECT 54.935 217.225 55.315 217.555 ;
        RECT 55.485 217.225 55.820 217.555 ;
        RECT 54.595 216.885 54.910 217.055 ;
        RECT 52.900 216.100 53.980 216.270 ;
        RECT 54.160 215.915 54.475 216.715 ;
        RECT 54.740 216.270 54.910 216.885 ;
        RECT 55.080 216.545 55.315 217.225 ;
        RECT 55.485 216.270 55.820 217.055 ;
        RECT 56.915 216.935 57.605 217.495 ;
        RECT 57.775 216.765 57.985 217.665 ;
        RECT 54.740 216.100 55.820 216.270 ;
        RECT 57.030 216.545 57.985 216.765 ;
        RECT 58.155 217.495 58.555 218.295 ;
        RECT 58.745 217.835 59.025 218.295 ;
        RECT 59.545 218.005 59.870 218.465 ;
        RECT 58.745 217.665 59.870 217.835 ;
        RECT 60.040 217.725 60.425 218.295 ;
        RECT 59.420 217.555 59.870 217.665 ;
        RECT 58.155 216.935 59.250 217.495 ;
        RECT 59.420 217.225 59.975 217.555 ;
        RECT 57.030 216.085 57.315 216.545 ;
        RECT 57.485 215.915 57.755 216.375 ;
        RECT 58.155 216.085 58.555 216.935 ;
        RECT 59.420 216.765 59.870 217.225 ;
        RECT 60.145 217.055 60.425 217.725 ;
        RECT 60.615 217.655 60.855 218.465 ;
        RECT 61.025 217.655 61.355 218.295 ;
        RECT 61.525 217.655 61.795 218.465 ;
        RECT 61.975 217.695 65.485 218.465 ;
        RECT 65.655 217.715 66.865 218.465 ;
        RECT 67.045 217.735 67.345 218.465 ;
        RECT 60.595 217.225 60.945 217.475 ;
        RECT 61.115 217.055 61.285 217.655 ;
        RECT 61.455 217.225 61.805 217.475 ;
        RECT 61.975 217.175 63.625 217.695 ;
        RECT 58.745 216.545 59.870 216.765 ;
        RECT 58.745 216.085 59.025 216.545 ;
        RECT 59.545 215.915 59.870 216.375 ;
        RECT 60.040 216.085 60.425 217.055 ;
        RECT 60.605 216.885 61.285 217.055 ;
        RECT 60.605 216.100 60.935 216.885 ;
        RECT 61.465 215.915 61.795 217.055 ;
        RECT 63.795 217.005 65.485 217.525 ;
        RECT 65.655 217.175 66.175 217.715 ;
        RECT 67.525 217.555 67.755 218.175 ;
        RECT 67.955 217.905 68.180 218.285 ;
        RECT 68.350 218.075 68.680 218.465 ;
        RECT 67.955 217.725 68.285 217.905 ;
        RECT 66.345 217.005 66.865 217.545 ;
        RECT 67.050 217.225 67.345 217.555 ;
        RECT 67.525 217.225 67.940 217.555 ;
        RECT 68.110 217.055 68.285 217.725 ;
        RECT 68.455 217.225 68.695 217.875 ;
        RECT 68.875 217.740 69.165 218.465 ;
        RECT 69.355 217.655 69.595 218.465 ;
        RECT 69.765 217.655 70.095 218.295 ;
        RECT 70.265 217.655 70.535 218.465 ;
        RECT 70.715 217.920 76.060 218.465 ;
        RECT 69.335 217.225 69.685 217.475 ;
        RECT 61.975 215.915 65.485 217.005 ;
        RECT 65.655 215.915 66.865 217.005 ;
        RECT 67.045 216.695 67.940 217.025 ;
        RECT 68.110 216.865 68.695 217.055 ;
        RECT 67.045 216.525 68.250 216.695 ;
        RECT 67.045 216.095 67.375 216.525 ;
        RECT 67.555 215.915 67.750 216.355 ;
        RECT 67.920 216.095 68.250 216.525 ;
        RECT 68.420 216.095 68.695 216.865 ;
        RECT 68.875 215.915 69.165 217.080 ;
        RECT 69.855 217.055 70.025 217.655 ;
        RECT 70.195 217.225 70.545 217.475 ;
        RECT 72.300 217.090 72.640 217.920 ;
        RECT 76.235 217.695 79.745 218.465 ;
        RECT 80.950 217.835 81.235 218.295 ;
        RECT 81.405 218.005 81.675 218.465 ;
        RECT 69.345 216.885 70.025 217.055 ;
        RECT 69.345 216.100 69.675 216.885 ;
        RECT 70.205 215.915 70.535 217.055 ;
        RECT 74.120 216.350 74.470 217.600 ;
        RECT 76.235 217.175 77.885 217.695 ;
        RECT 80.950 217.665 81.905 217.835 ;
        RECT 78.055 217.005 79.745 217.525 ;
        RECT 70.715 215.915 76.060 216.350 ;
        RECT 76.235 215.915 79.745 217.005 ;
        RECT 80.835 216.935 81.525 217.495 ;
        RECT 81.695 216.765 81.905 217.665 ;
        RECT 80.950 216.545 81.905 216.765 ;
        RECT 82.075 217.495 82.475 218.295 ;
        RECT 82.665 217.835 82.945 218.295 ;
        RECT 83.465 218.005 83.790 218.465 ;
        RECT 82.665 217.665 83.790 217.835 ;
        RECT 83.960 217.725 84.345 218.295 ;
        RECT 83.340 217.555 83.790 217.665 ;
        RECT 82.075 216.935 83.170 217.495 ;
        RECT 83.340 217.225 83.895 217.555 ;
        RECT 80.950 216.085 81.235 216.545 ;
        RECT 81.405 215.915 81.675 216.375 ;
        RECT 82.075 216.085 82.475 216.935 ;
        RECT 83.340 216.765 83.790 217.225 ;
        RECT 84.065 217.055 84.345 217.725 ;
        RECT 84.515 217.715 85.725 218.465 ;
        RECT 86.010 217.835 86.295 218.295 ;
        RECT 86.465 218.005 86.735 218.465 ;
        RECT 84.515 217.175 85.035 217.715 ;
        RECT 86.010 217.665 86.965 217.835 ;
        RECT 82.665 216.545 83.790 216.765 ;
        RECT 82.665 216.085 82.945 216.545 ;
        RECT 83.465 215.915 83.790 216.375 ;
        RECT 83.960 216.085 84.345 217.055 ;
        RECT 85.205 217.005 85.725 217.545 ;
        RECT 84.515 215.915 85.725 217.005 ;
        RECT 85.895 216.935 86.585 217.495 ;
        RECT 86.755 216.765 86.965 217.665 ;
        RECT 86.010 216.545 86.965 216.765 ;
        RECT 87.135 217.495 87.535 218.295 ;
        RECT 87.725 217.835 88.005 218.295 ;
        RECT 88.525 218.005 88.850 218.465 ;
        RECT 87.725 217.665 88.850 217.835 ;
        RECT 89.020 217.725 89.405 218.295 ;
        RECT 88.400 217.555 88.850 217.665 ;
        RECT 87.135 216.935 88.230 217.495 ;
        RECT 88.400 217.225 88.955 217.555 ;
        RECT 86.010 216.085 86.295 216.545 ;
        RECT 86.465 215.915 86.735 216.375 ;
        RECT 87.135 216.085 87.535 216.935 ;
        RECT 88.400 216.765 88.850 217.225 ;
        RECT 89.125 217.055 89.405 217.725 ;
        RECT 87.725 216.545 88.850 216.765 ;
        RECT 87.725 216.085 88.005 216.545 ;
        RECT 88.525 215.915 88.850 216.375 ;
        RECT 89.020 216.085 89.405 217.055 ;
        RECT 89.585 217.740 89.915 218.250 ;
        RECT 90.085 218.065 90.415 218.465 ;
        RECT 91.465 217.895 91.795 218.235 ;
        RECT 91.965 218.065 92.295 218.465 ;
        RECT 89.585 216.975 89.775 217.740 ;
        RECT 90.085 217.725 92.450 217.895 ;
        RECT 90.085 217.555 90.255 217.725 ;
        RECT 89.945 217.225 90.255 217.555 ;
        RECT 90.425 217.225 90.730 217.555 ;
        RECT 89.585 216.125 89.915 216.975 ;
        RECT 90.085 215.915 90.335 217.055 ;
        RECT 90.515 216.895 90.730 217.225 ;
        RECT 90.905 216.895 91.190 217.555 ;
        RECT 91.385 216.895 91.650 217.555 ;
        RECT 91.865 216.895 92.110 217.555 ;
        RECT 92.280 216.725 92.450 217.725 ;
        RECT 93.255 217.665 93.565 218.465 ;
        RECT 93.770 217.665 94.465 218.295 ;
        RECT 94.635 217.740 94.925 218.465 ;
        RECT 93.265 217.225 93.600 217.495 ;
        RECT 93.770 217.105 93.940 217.665 ;
        RECT 95.095 217.645 95.355 218.465 ;
        RECT 95.525 217.645 95.855 218.065 ;
        RECT 96.035 217.980 96.825 218.245 ;
        RECT 95.605 217.555 95.855 217.645 ;
        RECT 94.110 217.225 94.445 217.475 ;
        RECT 93.770 217.065 93.945 217.105 ;
        RECT 90.525 216.555 91.815 216.725 ;
        RECT 90.525 216.135 90.775 216.555 ;
        RECT 91.005 215.915 91.335 216.385 ;
        RECT 91.565 216.135 91.815 216.555 ;
        RECT 91.995 216.555 92.450 216.725 ;
        RECT 91.995 216.125 92.325 216.555 ;
        RECT 93.255 215.915 93.535 217.055 ;
        RECT 93.705 216.085 94.035 217.065 ;
        RECT 94.205 215.915 94.465 217.055 ;
        RECT 94.635 215.915 94.925 217.080 ;
        RECT 95.095 216.595 95.435 217.475 ;
        RECT 95.605 217.305 96.400 217.555 ;
        RECT 95.095 215.915 95.355 216.425 ;
        RECT 95.605 216.085 95.775 217.305 ;
        RECT 96.570 217.125 96.825 217.980 ;
        RECT 96.995 217.825 97.195 218.245 ;
        RECT 97.385 218.005 97.715 218.465 ;
        RECT 96.995 217.305 97.405 217.825 ;
        RECT 97.885 217.815 98.145 218.295 ;
        RECT 97.575 217.125 97.805 217.555 ;
        RECT 96.015 216.955 97.805 217.125 ;
        RECT 96.015 216.590 96.265 216.955 ;
        RECT 96.435 216.595 96.765 216.785 ;
        RECT 96.985 216.660 97.700 216.955 ;
        RECT 97.975 216.785 98.145 217.815 ;
        RECT 96.435 216.420 96.630 216.595 ;
        RECT 96.015 215.915 96.630 216.420 ;
        RECT 96.800 216.085 97.275 216.425 ;
        RECT 97.445 215.915 97.660 216.460 ;
        RECT 97.870 216.085 98.145 216.785 ;
        RECT 99.235 217.725 99.700 218.270 ;
        RECT 99.235 216.765 99.405 217.725 ;
        RECT 100.205 217.645 100.375 218.465 ;
        RECT 100.545 217.815 100.875 218.295 ;
        RECT 101.045 218.075 101.395 218.465 ;
        RECT 101.565 217.895 101.795 218.295 ;
        RECT 101.285 217.815 101.795 217.895 ;
        RECT 100.545 217.725 101.795 217.815 ;
        RECT 101.965 217.725 102.285 218.205 ;
        RECT 102.620 217.955 102.860 218.465 ;
        RECT 103.040 217.955 103.320 218.285 ;
        RECT 103.550 217.955 103.765 218.465 ;
        RECT 100.545 217.645 101.455 217.725 ;
        RECT 99.575 217.105 99.820 217.555 ;
        RECT 100.080 217.275 100.775 217.475 ;
        RECT 100.945 217.305 101.545 217.475 ;
        RECT 100.945 217.105 101.115 217.305 ;
        RECT 101.775 217.135 101.945 217.555 ;
        RECT 99.575 216.935 101.115 217.105 ;
        RECT 101.285 216.965 101.945 217.135 ;
        RECT 101.285 216.765 101.455 216.965 ;
        RECT 102.115 216.795 102.285 217.725 ;
        RECT 102.515 217.225 102.870 217.785 ;
        RECT 103.040 217.055 103.210 217.955 ;
        RECT 103.380 217.225 103.645 217.785 ;
        RECT 103.935 217.725 104.550 218.295 ;
        RECT 104.755 217.920 110.100 218.465 ;
        RECT 110.275 217.920 115.620 218.465 ;
        RECT 103.895 217.055 104.065 217.555 ;
        RECT 99.235 216.595 101.455 216.765 ;
        RECT 101.625 216.595 102.285 216.795 ;
        RECT 102.640 216.885 104.065 217.055 ;
        RECT 102.640 216.710 103.030 216.885 ;
        RECT 99.235 215.915 99.535 216.425 ;
        RECT 99.705 216.085 100.035 216.595 ;
        RECT 101.625 216.425 101.795 216.595 ;
        RECT 100.205 215.915 100.835 216.425 ;
        RECT 101.415 216.255 101.795 216.425 ;
        RECT 101.965 215.915 102.265 216.425 ;
        RECT 103.515 215.915 103.845 216.715 ;
        RECT 104.235 216.705 104.550 217.725 ;
        RECT 106.340 217.090 106.680 217.920 ;
        RECT 104.015 216.085 104.550 216.705 ;
        RECT 108.160 216.350 108.510 217.600 ;
        RECT 111.860 217.090 112.200 217.920 ;
        RECT 115.795 217.695 119.305 218.465 ;
        RECT 120.395 217.740 120.685 218.465 ;
        RECT 120.855 217.920 126.200 218.465 ;
        RECT 126.375 217.920 131.720 218.465 ;
        RECT 131.895 217.920 137.240 218.465 ;
        RECT 137.415 217.920 142.760 218.465 ;
        RECT 113.680 216.350 114.030 217.600 ;
        RECT 115.795 217.175 117.445 217.695 ;
        RECT 117.615 217.005 119.305 217.525 ;
        RECT 122.440 217.090 122.780 217.920 ;
        RECT 104.755 215.915 110.100 216.350 ;
        RECT 110.275 215.915 115.620 216.350 ;
        RECT 115.795 215.915 119.305 217.005 ;
        RECT 120.395 215.915 120.685 217.080 ;
        RECT 124.260 216.350 124.610 217.600 ;
        RECT 127.960 217.090 128.300 217.920 ;
        RECT 129.780 216.350 130.130 217.600 ;
        RECT 133.480 217.090 133.820 217.920 ;
        RECT 135.300 216.350 135.650 217.600 ;
        RECT 139.000 217.090 139.340 217.920 ;
        RECT 142.935 217.695 145.525 218.465 ;
        RECT 145.695 217.715 146.905 218.465 ;
        RECT 140.820 216.350 141.170 217.600 ;
        RECT 142.935 217.175 144.145 217.695 ;
        RECT 144.315 217.005 145.525 217.525 ;
        RECT 120.855 215.915 126.200 216.350 ;
        RECT 126.375 215.915 131.720 216.350 ;
        RECT 131.895 215.915 137.240 216.350 ;
        RECT 137.415 215.915 142.760 216.350 ;
        RECT 142.935 215.915 145.525 217.005 ;
        RECT 145.695 217.005 146.215 217.545 ;
        RECT 146.385 217.175 146.905 217.715 ;
        RECT 145.695 215.915 146.905 217.005 ;
        RECT 17.270 215.745 146.990 215.915 ;
        RECT 17.355 214.655 18.565 215.745 ;
        RECT 18.735 215.310 24.080 215.745 ;
        RECT 24.255 215.310 29.600 215.745 ;
        RECT 17.355 213.945 17.875 214.485 ;
        RECT 18.045 214.115 18.565 214.655 ;
        RECT 17.355 213.195 18.565 213.945 ;
        RECT 20.320 213.740 20.660 214.570 ;
        RECT 22.140 214.060 22.490 215.310 ;
        RECT 25.840 213.740 26.180 214.570 ;
        RECT 27.660 214.060 28.010 215.310 ;
        RECT 30.235 214.580 30.525 215.745 ;
        RECT 30.695 215.310 36.040 215.745 ;
        RECT 36.215 215.310 41.560 215.745 ;
        RECT 41.735 215.310 47.080 215.745 ;
        RECT 18.735 213.195 24.080 213.740 ;
        RECT 24.255 213.195 29.600 213.740 ;
        RECT 30.235 213.195 30.525 213.920 ;
        RECT 32.280 213.740 32.620 214.570 ;
        RECT 34.100 214.060 34.450 215.310 ;
        RECT 37.800 213.740 38.140 214.570 ;
        RECT 39.620 214.060 39.970 215.310 ;
        RECT 43.320 213.740 43.660 214.570 ;
        RECT 45.140 214.060 45.490 215.310 ;
        RECT 47.255 214.655 48.925 215.745 ;
        RECT 47.255 213.965 48.005 214.485 ;
        RECT 48.175 214.135 48.925 214.655 ;
        RECT 49.095 214.605 49.480 215.575 ;
        RECT 49.650 215.285 49.975 215.745 ;
        RECT 50.495 215.115 50.775 215.575 ;
        RECT 49.650 214.895 50.775 215.115 ;
        RECT 30.695 213.195 36.040 213.740 ;
        RECT 36.215 213.195 41.560 213.740 ;
        RECT 41.735 213.195 47.080 213.740 ;
        RECT 47.255 213.195 48.925 213.965 ;
        RECT 49.095 213.935 49.375 214.605 ;
        RECT 49.650 214.435 50.100 214.895 ;
        RECT 50.965 214.725 51.365 215.575 ;
        RECT 51.765 215.285 52.035 215.745 ;
        RECT 52.205 215.115 52.490 215.575 ;
        RECT 52.795 215.235 53.095 215.745 ;
        RECT 53.265 215.235 53.645 215.405 ;
        RECT 54.225 215.235 54.855 215.745 ;
        RECT 49.545 214.105 50.100 214.435 ;
        RECT 50.270 214.165 51.365 214.725 ;
        RECT 49.650 213.995 50.100 214.105 ;
        RECT 49.095 213.365 49.480 213.935 ;
        RECT 49.650 213.825 50.775 213.995 ;
        RECT 49.650 213.195 49.975 213.655 ;
        RECT 50.495 213.365 50.775 213.825 ;
        RECT 50.965 213.365 51.365 214.165 ;
        RECT 51.535 214.895 52.490 215.115 ;
        RECT 53.265 215.065 53.435 215.235 ;
        RECT 55.025 215.065 55.355 215.575 ;
        RECT 55.525 215.235 55.825 215.745 ;
        RECT 51.535 213.995 51.745 214.895 ;
        RECT 52.775 214.865 53.435 215.065 ;
        RECT 53.605 214.895 55.825 215.065 ;
        RECT 51.915 214.165 52.605 214.725 ;
        RECT 51.535 213.825 52.490 213.995 ;
        RECT 51.765 213.195 52.035 213.655 ;
        RECT 52.205 213.365 52.490 213.825 ;
        RECT 52.775 213.935 52.945 214.865 ;
        RECT 53.605 214.695 53.775 214.895 ;
        RECT 53.115 214.525 53.775 214.695 ;
        RECT 53.945 214.555 55.485 214.725 ;
        RECT 53.115 214.105 53.285 214.525 ;
        RECT 53.945 214.355 54.115 214.555 ;
        RECT 53.515 214.185 54.115 214.355 ;
        RECT 54.285 214.185 54.980 214.385 ;
        RECT 55.240 214.105 55.485 214.555 ;
        RECT 53.605 213.935 54.515 214.015 ;
        RECT 52.775 213.455 53.095 213.935 ;
        RECT 53.265 213.845 54.515 213.935 ;
        RECT 53.265 213.765 53.775 213.845 ;
        RECT 53.265 213.365 53.495 213.765 ;
        RECT 53.665 213.195 54.015 213.585 ;
        RECT 54.185 213.365 54.515 213.845 ;
        RECT 54.685 213.195 54.855 214.015 ;
        RECT 55.655 213.935 55.825 214.895 ;
        RECT 55.995 214.580 56.285 215.745 ;
        RECT 56.515 214.685 56.845 215.530 ;
        RECT 57.015 214.735 57.185 215.745 ;
        RECT 57.355 215.015 57.695 215.575 ;
        RECT 57.925 215.245 58.240 215.745 ;
        RECT 58.420 215.275 59.305 215.445 ;
        RECT 56.455 214.605 56.845 214.685 ;
        RECT 57.355 214.640 58.250 215.015 ;
        RECT 55.360 213.390 55.825 213.935 ;
        RECT 56.455 214.555 56.670 214.605 ;
        RECT 56.455 213.975 56.625 214.555 ;
        RECT 57.355 214.435 57.545 214.640 ;
        RECT 58.420 214.435 58.590 215.275 ;
        RECT 59.530 215.245 59.780 215.575 ;
        RECT 56.795 214.105 57.545 214.435 ;
        RECT 57.715 214.105 58.590 214.435 ;
        RECT 56.455 213.935 56.680 213.975 ;
        RECT 57.345 213.935 57.545 214.105 ;
        RECT 55.995 213.195 56.285 213.920 ;
        RECT 56.455 213.850 56.835 213.935 ;
        RECT 56.505 213.415 56.835 213.850 ;
        RECT 57.005 213.195 57.175 213.805 ;
        RECT 57.345 213.410 57.675 213.935 ;
        RECT 57.935 213.195 58.145 213.725 ;
        RECT 58.420 213.645 58.590 214.105 ;
        RECT 58.760 214.145 59.080 215.105 ;
        RECT 59.250 214.355 59.440 215.075 ;
        RECT 59.610 214.175 59.780 215.245 ;
        RECT 59.950 214.945 60.120 215.745 ;
        RECT 60.290 215.300 61.395 215.470 ;
        RECT 60.290 214.685 60.460 215.300 ;
        RECT 61.605 215.150 61.855 215.575 ;
        RECT 62.025 215.285 62.290 215.745 ;
        RECT 60.630 214.765 61.160 215.130 ;
        RECT 61.605 215.020 61.910 215.150 ;
        RECT 59.950 214.595 60.460 214.685 ;
        RECT 59.950 214.425 60.820 214.595 ;
        RECT 59.950 214.355 60.120 214.425 ;
        RECT 60.240 214.175 60.440 214.205 ;
        RECT 58.760 213.815 59.225 214.145 ;
        RECT 59.610 213.875 60.440 214.175 ;
        RECT 59.610 213.645 59.780 213.875 ;
        RECT 58.420 213.475 59.205 213.645 ;
        RECT 59.375 213.475 59.780 213.645 ;
        RECT 59.960 213.195 60.330 213.695 ;
        RECT 60.650 213.645 60.820 214.425 ;
        RECT 60.990 214.065 61.160 214.765 ;
        RECT 61.330 214.235 61.570 214.830 ;
        RECT 60.990 213.845 61.515 214.065 ;
        RECT 61.740 213.915 61.910 215.020 ;
        RECT 61.685 213.785 61.910 213.915 ;
        RECT 62.080 213.825 62.360 214.775 ;
        RECT 61.685 213.645 61.855 213.785 ;
        RECT 60.650 213.475 61.325 213.645 ;
        RECT 61.520 213.475 61.855 213.645 ;
        RECT 62.025 213.195 62.275 213.655 ;
        RECT 62.530 213.455 62.715 215.575 ;
        RECT 62.885 215.245 63.215 215.745 ;
        RECT 63.385 215.075 63.555 215.575 ;
        RECT 62.890 214.905 63.555 215.075 ;
        RECT 62.890 213.915 63.120 214.905 ;
        RECT 63.290 214.085 63.640 214.735 ;
        RECT 64.335 214.685 64.665 215.530 ;
        RECT 64.835 214.735 65.005 215.745 ;
        RECT 65.175 215.015 65.515 215.575 ;
        RECT 65.745 215.245 66.060 215.745 ;
        RECT 66.240 215.275 67.125 215.445 ;
        RECT 64.275 214.605 64.665 214.685 ;
        RECT 65.175 214.640 66.070 215.015 ;
        RECT 64.275 214.555 64.490 214.605 ;
        RECT 64.275 213.975 64.445 214.555 ;
        RECT 65.175 214.435 65.365 214.640 ;
        RECT 66.240 214.435 66.410 215.275 ;
        RECT 67.350 215.245 67.600 215.575 ;
        RECT 64.615 214.105 65.365 214.435 ;
        RECT 65.535 214.105 66.410 214.435 ;
        RECT 64.275 213.935 64.500 213.975 ;
        RECT 65.165 213.935 65.365 214.105 ;
        RECT 62.890 213.745 63.555 213.915 ;
        RECT 64.275 213.850 64.655 213.935 ;
        RECT 62.885 213.195 63.215 213.575 ;
        RECT 63.385 213.455 63.555 213.745 ;
        RECT 64.325 213.415 64.655 213.850 ;
        RECT 64.825 213.195 64.995 213.805 ;
        RECT 65.165 213.410 65.495 213.935 ;
        RECT 65.755 213.195 65.965 213.725 ;
        RECT 66.240 213.645 66.410 214.105 ;
        RECT 66.580 214.145 66.900 215.105 ;
        RECT 67.070 214.355 67.260 215.075 ;
        RECT 67.430 214.175 67.600 215.245 ;
        RECT 67.770 214.945 67.940 215.745 ;
        RECT 68.110 215.300 69.215 215.470 ;
        RECT 68.110 214.685 68.280 215.300 ;
        RECT 69.425 215.150 69.675 215.575 ;
        RECT 69.845 215.285 70.110 215.745 ;
        RECT 68.450 214.765 68.980 215.130 ;
        RECT 69.425 215.020 69.730 215.150 ;
        RECT 67.770 214.595 68.280 214.685 ;
        RECT 67.770 214.425 68.640 214.595 ;
        RECT 67.770 214.355 67.940 214.425 ;
        RECT 68.060 214.175 68.260 214.205 ;
        RECT 66.580 213.815 67.045 214.145 ;
        RECT 67.430 213.875 68.260 214.175 ;
        RECT 67.430 213.645 67.600 213.875 ;
        RECT 66.240 213.475 67.025 213.645 ;
        RECT 67.195 213.475 67.600 213.645 ;
        RECT 67.780 213.195 68.150 213.695 ;
        RECT 68.470 213.645 68.640 214.425 ;
        RECT 68.810 214.065 68.980 214.765 ;
        RECT 69.150 214.235 69.390 214.830 ;
        RECT 68.810 213.845 69.335 214.065 ;
        RECT 69.560 213.915 69.730 215.020 ;
        RECT 69.505 213.785 69.730 213.915 ;
        RECT 69.900 213.825 70.180 214.775 ;
        RECT 69.505 213.645 69.675 213.785 ;
        RECT 68.470 213.475 69.145 213.645 ;
        RECT 69.340 213.475 69.675 213.645 ;
        RECT 69.845 213.195 70.095 213.655 ;
        RECT 70.350 213.455 70.535 215.575 ;
        RECT 70.705 215.245 71.035 215.745 ;
        RECT 71.205 215.075 71.375 215.575 ;
        RECT 71.635 215.310 76.980 215.745 ;
        RECT 70.710 214.905 71.375 215.075 ;
        RECT 70.710 213.915 70.940 214.905 ;
        RECT 71.110 214.085 71.460 214.735 ;
        RECT 70.710 213.745 71.375 213.915 ;
        RECT 70.705 213.195 71.035 213.575 ;
        RECT 71.205 213.455 71.375 213.745 ;
        RECT 73.220 213.740 73.560 214.570 ;
        RECT 75.040 214.060 75.390 215.310 ;
        RECT 77.155 214.655 80.665 215.745 ;
        RECT 77.155 213.965 78.805 214.485 ;
        RECT 78.975 214.135 80.665 214.655 ;
        RECT 81.755 214.580 82.045 215.745 ;
        RECT 82.735 214.685 83.065 215.530 ;
        RECT 83.235 214.735 83.405 215.745 ;
        RECT 83.575 215.015 83.915 215.575 ;
        RECT 84.145 215.245 84.460 215.745 ;
        RECT 84.640 215.275 85.525 215.445 ;
        RECT 82.675 214.605 83.065 214.685 ;
        RECT 83.575 214.640 84.470 215.015 ;
        RECT 82.675 214.555 82.890 214.605 ;
        RECT 82.675 213.975 82.845 214.555 ;
        RECT 83.575 214.435 83.765 214.640 ;
        RECT 84.640 214.435 84.810 215.275 ;
        RECT 85.750 215.245 86.000 215.575 ;
        RECT 83.015 214.105 83.765 214.435 ;
        RECT 83.935 214.105 84.810 214.435 ;
        RECT 71.635 213.195 76.980 213.740 ;
        RECT 77.155 213.195 80.665 213.965 ;
        RECT 82.675 213.935 82.900 213.975 ;
        RECT 83.565 213.935 83.765 214.105 ;
        RECT 81.755 213.195 82.045 213.920 ;
        RECT 82.675 213.850 83.055 213.935 ;
        RECT 82.725 213.415 83.055 213.850 ;
        RECT 83.225 213.195 83.395 213.805 ;
        RECT 83.565 213.410 83.895 213.935 ;
        RECT 84.155 213.195 84.365 213.725 ;
        RECT 84.640 213.645 84.810 214.105 ;
        RECT 84.980 214.145 85.300 215.105 ;
        RECT 85.470 214.355 85.660 215.075 ;
        RECT 85.830 214.175 86.000 215.245 ;
        RECT 86.170 214.945 86.340 215.745 ;
        RECT 86.510 215.300 87.615 215.470 ;
        RECT 86.510 214.685 86.680 215.300 ;
        RECT 87.825 215.150 88.075 215.575 ;
        RECT 88.245 215.285 88.510 215.745 ;
        RECT 86.850 214.765 87.380 215.130 ;
        RECT 87.825 215.020 88.130 215.150 ;
        RECT 86.170 214.595 86.680 214.685 ;
        RECT 86.170 214.425 87.040 214.595 ;
        RECT 86.170 214.355 86.340 214.425 ;
        RECT 86.460 214.175 86.660 214.205 ;
        RECT 84.980 213.815 85.445 214.145 ;
        RECT 85.830 213.875 86.660 214.175 ;
        RECT 85.830 213.645 86.000 213.875 ;
        RECT 84.640 213.475 85.425 213.645 ;
        RECT 85.595 213.475 86.000 213.645 ;
        RECT 86.180 213.195 86.550 213.695 ;
        RECT 86.870 213.645 87.040 214.425 ;
        RECT 87.210 214.065 87.380 214.765 ;
        RECT 87.550 214.235 87.790 214.830 ;
        RECT 87.210 213.845 87.735 214.065 ;
        RECT 87.960 213.915 88.130 215.020 ;
        RECT 87.905 213.785 88.130 213.915 ;
        RECT 88.300 213.825 88.580 214.775 ;
        RECT 87.905 213.645 88.075 213.785 ;
        RECT 86.870 213.475 87.545 213.645 ;
        RECT 87.740 213.475 88.075 213.645 ;
        RECT 88.245 213.195 88.495 213.655 ;
        RECT 88.750 213.455 88.935 215.575 ;
        RECT 89.105 215.245 89.435 215.745 ;
        RECT 89.605 215.075 89.775 215.575 ;
        RECT 89.110 214.905 89.775 215.075 ;
        RECT 90.125 215.075 90.295 215.575 ;
        RECT 90.465 215.245 90.795 215.745 ;
        RECT 90.125 214.905 90.790 215.075 ;
        RECT 89.110 213.915 89.340 214.905 ;
        RECT 89.510 214.085 89.860 214.735 ;
        RECT 90.040 214.085 90.390 214.735 ;
        RECT 90.560 213.915 90.790 214.905 ;
        RECT 89.110 213.745 89.775 213.915 ;
        RECT 89.105 213.195 89.435 213.575 ;
        RECT 89.605 213.455 89.775 213.745 ;
        RECT 90.125 213.745 90.790 213.915 ;
        RECT 90.125 213.455 90.295 213.745 ;
        RECT 90.465 213.195 90.795 213.575 ;
        RECT 90.965 213.455 91.150 215.575 ;
        RECT 91.390 215.285 91.655 215.745 ;
        RECT 91.825 215.150 92.075 215.575 ;
        RECT 92.285 215.300 93.390 215.470 ;
        RECT 91.770 215.020 92.075 215.150 ;
        RECT 91.320 213.825 91.600 214.775 ;
        RECT 91.770 213.915 91.940 215.020 ;
        RECT 92.110 214.235 92.350 214.830 ;
        RECT 92.520 214.765 93.050 215.130 ;
        RECT 92.520 214.065 92.690 214.765 ;
        RECT 93.220 214.685 93.390 215.300 ;
        RECT 93.560 214.945 93.730 215.745 ;
        RECT 93.900 215.245 94.150 215.575 ;
        RECT 94.375 215.275 95.260 215.445 ;
        RECT 93.220 214.595 93.730 214.685 ;
        RECT 91.770 213.785 91.995 213.915 ;
        RECT 92.165 213.845 92.690 214.065 ;
        RECT 92.860 214.425 93.730 214.595 ;
        RECT 91.405 213.195 91.655 213.655 ;
        RECT 91.825 213.645 91.995 213.785 ;
        RECT 92.860 213.645 93.030 214.425 ;
        RECT 93.560 214.355 93.730 214.425 ;
        RECT 93.240 214.175 93.440 214.205 ;
        RECT 93.900 214.175 94.070 215.245 ;
        RECT 94.240 214.355 94.430 215.075 ;
        RECT 93.240 213.875 94.070 214.175 ;
        RECT 94.600 214.145 94.920 215.105 ;
        RECT 91.825 213.475 92.160 213.645 ;
        RECT 92.355 213.475 93.030 213.645 ;
        RECT 93.350 213.195 93.720 213.695 ;
        RECT 93.900 213.645 94.070 213.875 ;
        RECT 94.455 213.815 94.920 214.145 ;
        RECT 95.090 214.435 95.260 215.275 ;
        RECT 95.440 215.245 95.755 215.745 ;
        RECT 95.985 215.015 96.325 215.575 ;
        RECT 95.430 214.640 96.325 215.015 ;
        RECT 96.495 214.735 96.665 215.745 ;
        RECT 96.135 214.435 96.325 214.640 ;
        RECT 96.835 214.685 97.165 215.530 ;
        RECT 97.485 215.075 97.655 215.575 ;
        RECT 97.825 215.245 98.155 215.745 ;
        RECT 97.485 214.905 98.150 215.075 ;
        RECT 96.835 214.605 97.225 214.685 ;
        RECT 97.010 214.555 97.225 214.605 ;
        RECT 95.090 214.105 95.965 214.435 ;
        RECT 96.135 214.105 96.885 214.435 ;
        RECT 95.090 213.645 95.260 214.105 ;
        RECT 96.135 213.935 96.335 214.105 ;
        RECT 97.055 213.975 97.225 214.555 ;
        RECT 97.400 214.085 97.750 214.735 ;
        RECT 97.000 213.935 97.225 213.975 ;
        RECT 93.900 213.475 94.305 213.645 ;
        RECT 94.475 213.475 95.260 213.645 ;
        RECT 95.535 213.195 95.745 213.725 ;
        RECT 96.005 213.410 96.335 213.935 ;
        RECT 96.845 213.850 97.225 213.935 ;
        RECT 97.920 213.915 98.150 214.905 ;
        RECT 96.505 213.195 96.675 213.805 ;
        RECT 96.845 213.415 97.175 213.850 ;
        RECT 97.485 213.745 98.150 213.915 ;
        RECT 97.485 213.455 97.655 213.745 ;
        RECT 97.825 213.195 98.155 213.575 ;
        RECT 98.325 213.455 98.510 215.575 ;
        RECT 98.750 215.285 99.015 215.745 ;
        RECT 99.185 215.150 99.435 215.575 ;
        RECT 99.645 215.300 100.750 215.470 ;
        RECT 99.130 215.020 99.435 215.150 ;
        RECT 98.680 213.825 98.960 214.775 ;
        RECT 99.130 213.915 99.300 215.020 ;
        RECT 99.470 214.235 99.710 214.830 ;
        RECT 99.880 214.765 100.410 215.130 ;
        RECT 99.880 214.065 100.050 214.765 ;
        RECT 100.580 214.685 100.750 215.300 ;
        RECT 100.920 214.945 101.090 215.745 ;
        RECT 101.260 215.245 101.510 215.575 ;
        RECT 101.735 215.275 102.620 215.445 ;
        RECT 100.580 214.595 101.090 214.685 ;
        RECT 99.130 213.785 99.355 213.915 ;
        RECT 99.525 213.845 100.050 214.065 ;
        RECT 100.220 214.425 101.090 214.595 ;
        RECT 98.765 213.195 99.015 213.655 ;
        RECT 99.185 213.645 99.355 213.785 ;
        RECT 100.220 213.645 100.390 214.425 ;
        RECT 100.920 214.355 101.090 214.425 ;
        RECT 100.600 214.175 100.800 214.205 ;
        RECT 101.260 214.175 101.430 215.245 ;
        RECT 101.600 214.355 101.790 215.075 ;
        RECT 100.600 213.875 101.430 214.175 ;
        RECT 101.960 214.145 102.280 215.105 ;
        RECT 99.185 213.475 99.520 213.645 ;
        RECT 99.715 213.475 100.390 213.645 ;
        RECT 100.710 213.195 101.080 213.695 ;
        RECT 101.260 213.645 101.430 213.875 ;
        RECT 101.815 213.815 102.280 214.145 ;
        RECT 102.450 214.435 102.620 215.275 ;
        RECT 102.800 215.245 103.115 215.745 ;
        RECT 103.345 215.015 103.685 215.575 ;
        RECT 102.790 214.640 103.685 215.015 ;
        RECT 103.855 214.735 104.025 215.745 ;
        RECT 103.495 214.435 103.685 214.640 ;
        RECT 104.195 214.685 104.525 215.530 ;
        RECT 104.810 214.875 105.095 215.745 ;
        RECT 105.265 215.115 105.525 215.575 ;
        RECT 105.700 215.285 105.955 215.745 ;
        RECT 106.125 215.115 106.385 215.575 ;
        RECT 105.265 214.945 106.385 215.115 ;
        RECT 106.555 214.945 106.865 215.745 ;
        RECT 105.265 214.695 105.525 214.945 ;
        RECT 107.035 214.775 107.345 215.575 ;
        RECT 104.195 214.605 104.585 214.685 ;
        RECT 104.370 214.555 104.585 214.605 ;
        RECT 102.450 214.105 103.325 214.435 ;
        RECT 103.495 214.105 104.245 214.435 ;
        RECT 102.450 213.645 102.620 214.105 ;
        RECT 103.495 213.935 103.695 214.105 ;
        RECT 104.415 213.975 104.585 214.555 ;
        RECT 104.360 213.935 104.585 213.975 ;
        RECT 101.260 213.475 101.665 213.645 ;
        RECT 101.835 213.475 102.620 213.645 ;
        RECT 102.895 213.195 103.105 213.725 ;
        RECT 103.365 213.410 103.695 213.935 ;
        RECT 104.205 213.850 104.585 213.935 ;
        RECT 104.770 214.525 105.525 214.695 ;
        RECT 106.315 214.605 107.345 214.775 ;
        RECT 104.770 214.015 105.175 214.525 ;
        RECT 106.315 214.355 106.485 214.605 ;
        RECT 105.345 214.185 106.485 214.355 ;
        RECT 103.865 213.195 104.035 213.805 ;
        RECT 104.205 213.415 104.535 213.850 ;
        RECT 104.770 213.845 106.420 214.015 ;
        RECT 106.655 213.865 107.005 214.435 ;
        RECT 104.815 213.195 105.095 213.675 ;
        RECT 105.265 213.455 105.525 213.845 ;
        RECT 105.700 213.195 105.955 213.675 ;
        RECT 106.125 213.455 106.420 213.845 ;
        RECT 107.175 213.695 107.345 214.605 ;
        RECT 107.515 214.580 107.805 215.745 ;
        RECT 107.975 215.310 113.320 215.745 ;
        RECT 113.495 215.310 118.840 215.745 ;
        RECT 119.015 215.310 124.360 215.745 ;
        RECT 124.535 215.310 129.880 215.745 ;
        RECT 106.600 213.195 106.875 213.675 ;
        RECT 107.045 213.365 107.345 213.695 ;
        RECT 107.515 213.195 107.805 213.920 ;
        RECT 109.560 213.740 109.900 214.570 ;
        RECT 111.380 214.060 111.730 215.310 ;
        RECT 115.080 213.740 115.420 214.570 ;
        RECT 116.900 214.060 117.250 215.310 ;
        RECT 120.600 213.740 120.940 214.570 ;
        RECT 122.420 214.060 122.770 215.310 ;
        RECT 126.120 213.740 126.460 214.570 ;
        RECT 127.940 214.060 128.290 215.310 ;
        RECT 130.055 214.655 132.645 215.745 ;
        RECT 130.055 213.965 131.265 214.485 ;
        RECT 131.435 214.135 132.645 214.655 ;
        RECT 133.275 214.580 133.565 215.745 ;
        RECT 133.735 215.310 139.080 215.745 ;
        RECT 139.255 215.310 144.600 215.745 ;
        RECT 107.975 213.195 113.320 213.740 ;
        RECT 113.495 213.195 118.840 213.740 ;
        RECT 119.015 213.195 124.360 213.740 ;
        RECT 124.535 213.195 129.880 213.740 ;
        RECT 130.055 213.195 132.645 213.965 ;
        RECT 133.275 213.195 133.565 213.920 ;
        RECT 135.320 213.740 135.660 214.570 ;
        RECT 137.140 214.060 137.490 215.310 ;
        RECT 140.840 213.740 141.180 214.570 ;
        RECT 142.660 214.060 143.010 215.310 ;
        RECT 145.695 214.655 146.905 215.745 ;
        RECT 145.695 214.115 146.215 214.655 ;
        RECT 146.385 213.945 146.905 214.485 ;
        RECT 133.735 213.195 139.080 213.740 ;
        RECT 139.255 213.195 144.600 213.740 ;
        RECT 145.695 213.195 146.905 213.945 ;
        RECT 17.270 213.025 146.990 213.195 ;
        RECT 17.355 212.275 18.565 213.025 ;
        RECT 18.735 212.480 24.080 213.025 ;
        RECT 24.255 212.480 29.600 213.025 ;
        RECT 29.775 212.480 35.120 213.025 ;
        RECT 35.295 212.480 40.640 213.025 ;
        RECT 17.355 211.735 17.875 212.275 ;
        RECT 18.045 211.565 18.565 212.105 ;
        RECT 20.320 211.650 20.660 212.480 ;
        RECT 17.355 210.475 18.565 211.565 ;
        RECT 22.140 210.910 22.490 212.160 ;
        RECT 25.840 211.650 26.180 212.480 ;
        RECT 27.660 210.910 28.010 212.160 ;
        RECT 31.360 211.650 31.700 212.480 ;
        RECT 33.180 210.910 33.530 212.160 ;
        RECT 36.880 211.650 37.220 212.480 ;
        RECT 40.815 212.255 42.485 213.025 ;
        RECT 43.115 212.300 43.405 213.025 ;
        RECT 43.575 212.275 44.785 213.025 ;
        RECT 38.700 210.910 39.050 212.160 ;
        RECT 40.815 211.735 41.565 212.255 ;
        RECT 41.735 211.565 42.485 212.085 ;
        RECT 43.575 211.735 44.095 212.275 ;
        RECT 44.965 212.215 45.235 213.025 ;
        RECT 45.405 212.215 45.735 212.855 ;
        RECT 45.905 212.215 46.145 213.025 ;
        RECT 46.425 212.475 46.595 212.765 ;
        RECT 46.765 212.645 47.095 213.025 ;
        RECT 46.425 212.305 47.090 212.475 ;
        RECT 18.735 210.475 24.080 210.910 ;
        RECT 24.255 210.475 29.600 210.910 ;
        RECT 29.775 210.475 35.120 210.910 ;
        RECT 35.295 210.475 40.640 210.910 ;
        RECT 40.815 210.475 42.485 211.565 ;
        RECT 43.115 210.475 43.405 211.640 ;
        RECT 44.265 211.565 44.785 212.105 ;
        RECT 44.955 211.785 45.305 212.035 ;
        RECT 45.475 211.615 45.645 212.215 ;
        RECT 45.815 211.785 46.165 212.035 ;
        RECT 43.575 210.475 44.785 211.565 ;
        RECT 44.965 210.475 45.295 211.615 ;
        RECT 45.475 211.445 46.155 211.615 ;
        RECT 46.340 211.485 46.690 212.135 ;
        RECT 45.825 210.660 46.155 211.445 ;
        RECT 46.860 211.315 47.090 212.305 ;
        RECT 46.425 211.145 47.090 211.315 ;
        RECT 46.425 210.645 46.595 211.145 ;
        RECT 46.765 210.475 47.095 210.975 ;
        RECT 47.265 210.645 47.450 212.765 ;
        RECT 47.705 212.565 47.955 213.025 ;
        RECT 48.125 212.575 48.460 212.745 ;
        RECT 48.655 212.575 49.330 212.745 ;
        RECT 48.125 212.435 48.295 212.575 ;
        RECT 47.620 211.445 47.900 212.395 ;
        RECT 48.070 212.305 48.295 212.435 ;
        RECT 48.070 211.200 48.240 212.305 ;
        RECT 48.465 212.155 48.990 212.375 ;
        RECT 48.410 211.390 48.650 211.985 ;
        RECT 48.820 211.455 48.990 212.155 ;
        RECT 49.160 211.795 49.330 212.575 ;
        RECT 49.650 212.525 50.020 213.025 ;
        RECT 50.200 212.575 50.605 212.745 ;
        RECT 50.775 212.575 51.560 212.745 ;
        RECT 50.200 212.345 50.370 212.575 ;
        RECT 49.540 212.045 50.370 212.345 ;
        RECT 50.755 212.075 51.220 212.405 ;
        RECT 49.540 212.015 49.740 212.045 ;
        RECT 49.860 211.795 50.030 211.865 ;
        RECT 49.160 211.625 50.030 211.795 ;
        RECT 49.520 211.535 50.030 211.625 ;
        RECT 48.070 211.070 48.375 211.200 ;
        RECT 48.820 211.090 49.350 211.455 ;
        RECT 47.690 210.475 47.955 210.935 ;
        RECT 48.125 210.645 48.375 211.070 ;
        RECT 49.520 210.920 49.690 211.535 ;
        RECT 48.585 210.750 49.690 210.920 ;
        RECT 49.860 210.475 50.030 211.275 ;
        RECT 50.200 210.975 50.370 212.045 ;
        RECT 50.540 211.145 50.730 211.865 ;
        RECT 50.900 211.115 51.220 212.075 ;
        RECT 51.390 212.115 51.560 212.575 ;
        RECT 51.835 212.495 52.045 213.025 ;
        RECT 52.305 212.285 52.635 212.810 ;
        RECT 52.805 212.415 52.975 213.025 ;
        RECT 53.145 212.370 53.475 212.805 ;
        RECT 53.785 212.475 53.955 212.765 ;
        RECT 54.125 212.645 54.455 213.025 ;
        RECT 53.145 212.285 53.525 212.370 ;
        RECT 53.785 212.305 54.450 212.475 ;
        RECT 52.435 212.115 52.635 212.285 ;
        RECT 53.300 212.245 53.525 212.285 ;
        RECT 51.390 211.785 52.265 212.115 ;
        RECT 52.435 211.785 53.185 212.115 ;
        RECT 50.200 210.645 50.450 210.975 ;
        RECT 51.390 210.945 51.560 211.785 ;
        RECT 52.435 211.580 52.625 211.785 ;
        RECT 53.355 211.665 53.525 212.245 ;
        RECT 53.310 211.615 53.525 211.665 ;
        RECT 51.730 211.205 52.625 211.580 ;
        RECT 53.135 211.535 53.525 211.615 ;
        RECT 50.675 210.775 51.560 210.945 ;
        RECT 51.740 210.475 52.055 210.975 ;
        RECT 52.285 210.645 52.625 211.205 ;
        RECT 52.795 210.475 52.965 211.485 ;
        RECT 53.135 210.690 53.465 211.535 ;
        RECT 53.700 211.485 54.050 212.135 ;
        RECT 54.220 211.315 54.450 212.305 ;
        RECT 53.785 211.145 54.450 211.315 ;
        RECT 53.785 210.645 53.955 211.145 ;
        RECT 54.125 210.475 54.455 210.975 ;
        RECT 54.625 210.645 54.810 212.765 ;
        RECT 55.065 212.565 55.315 213.025 ;
        RECT 55.485 212.575 55.820 212.745 ;
        RECT 56.015 212.575 56.690 212.745 ;
        RECT 55.485 212.435 55.655 212.575 ;
        RECT 54.980 211.445 55.260 212.395 ;
        RECT 55.430 212.305 55.655 212.435 ;
        RECT 55.430 211.200 55.600 212.305 ;
        RECT 55.825 212.155 56.350 212.375 ;
        RECT 55.770 211.390 56.010 211.985 ;
        RECT 56.180 211.455 56.350 212.155 ;
        RECT 56.520 211.795 56.690 212.575 ;
        RECT 57.010 212.525 57.380 213.025 ;
        RECT 57.560 212.575 57.965 212.745 ;
        RECT 58.135 212.575 58.920 212.745 ;
        RECT 57.560 212.345 57.730 212.575 ;
        RECT 56.900 212.045 57.730 212.345 ;
        RECT 58.115 212.075 58.580 212.405 ;
        RECT 56.900 212.015 57.100 212.045 ;
        RECT 57.220 211.795 57.390 211.865 ;
        RECT 56.520 211.625 57.390 211.795 ;
        RECT 56.880 211.535 57.390 211.625 ;
        RECT 55.430 211.070 55.735 211.200 ;
        RECT 56.180 211.090 56.710 211.455 ;
        RECT 55.050 210.475 55.315 210.935 ;
        RECT 55.485 210.645 55.735 211.070 ;
        RECT 56.880 210.920 57.050 211.535 ;
        RECT 55.945 210.750 57.050 210.920 ;
        RECT 57.220 210.475 57.390 211.275 ;
        RECT 57.560 210.975 57.730 212.045 ;
        RECT 57.900 211.145 58.090 211.865 ;
        RECT 58.260 211.115 58.580 212.075 ;
        RECT 58.750 212.115 58.920 212.575 ;
        RECT 59.195 212.495 59.405 213.025 ;
        RECT 59.665 212.285 59.995 212.810 ;
        RECT 60.165 212.415 60.335 213.025 ;
        RECT 60.505 212.370 60.835 212.805 ;
        RECT 60.505 212.285 60.885 212.370 ;
        RECT 59.795 212.115 59.995 212.285 ;
        RECT 60.660 212.245 60.885 212.285 ;
        RECT 58.750 211.785 59.625 212.115 ;
        RECT 59.795 211.785 60.545 212.115 ;
        RECT 57.560 210.645 57.810 210.975 ;
        RECT 58.750 210.945 58.920 211.785 ;
        RECT 59.795 211.580 59.985 211.785 ;
        RECT 60.715 211.665 60.885 212.245 ;
        RECT 60.670 211.615 60.885 211.665 ;
        RECT 59.090 211.205 59.985 211.580 ;
        RECT 60.495 211.535 60.885 211.615 ;
        RECT 61.055 212.285 61.440 212.855 ;
        RECT 61.610 212.565 61.935 213.025 ;
        RECT 62.455 212.395 62.735 212.855 ;
        RECT 61.055 211.615 61.335 212.285 ;
        RECT 61.610 212.225 62.735 212.395 ;
        RECT 61.610 212.115 62.060 212.225 ;
        RECT 61.505 211.785 62.060 212.115 ;
        RECT 62.925 212.055 63.325 212.855 ;
        RECT 63.725 212.565 63.995 213.025 ;
        RECT 64.165 212.395 64.450 212.855 ;
        RECT 58.035 210.775 58.920 210.945 ;
        RECT 59.100 210.475 59.415 210.975 ;
        RECT 59.645 210.645 59.985 211.205 ;
        RECT 60.155 210.475 60.325 211.485 ;
        RECT 60.495 210.690 60.825 211.535 ;
        RECT 61.055 210.645 61.440 211.615 ;
        RECT 61.610 211.325 62.060 211.785 ;
        RECT 62.230 211.495 63.325 212.055 ;
        RECT 61.610 211.105 62.735 211.325 ;
        RECT 61.610 210.475 61.935 210.935 ;
        RECT 62.455 210.645 62.735 211.105 ;
        RECT 62.925 210.645 63.325 211.495 ;
        RECT 63.495 212.225 64.450 212.395 ;
        RECT 65.310 212.395 65.595 212.855 ;
        RECT 65.765 212.565 66.035 213.025 ;
        RECT 65.310 212.225 66.265 212.395 ;
        RECT 63.495 211.325 63.705 212.225 ;
        RECT 63.875 211.495 64.565 212.055 ;
        RECT 65.195 211.495 65.885 212.055 ;
        RECT 66.055 211.325 66.265 212.225 ;
        RECT 63.495 211.105 64.450 211.325 ;
        RECT 63.725 210.475 63.995 210.935 ;
        RECT 64.165 210.645 64.450 211.105 ;
        RECT 65.310 211.105 66.265 211.325 ;
        RECT 66.435 212.055 66.835 212.855 ;
        RECT 67.025 212.395 67.305 212.855 ;
        RECT 67.825 212.565 68.150 213.025 ;
        RECT 67.025 212.225 68.150 212.395 ;
        RECT 68.320 212.285 68.705 212.855 ;
        RECT 68.875 212.300 69.165 213.025 ;
        RECT 69.490 212.375 69.820 212.840 ;
        RECT 69.990 212.555 70.160 213.025 ;
        RECT 70.330 212.375 70.660 212.855 ;
        RECT 67.700 212.115 68.150 212.225 ;
        RECT 66.435 211.495 67.530 212.055 ;
        RECT 67.700 211.785 68.255 212.115 ;
        RECT 65.310 210.645 65.595 211.105 ;
        RECT 65.765 210.475 66.035 210.935 ;
        RECT 66.435 210.645 66.835 211.495 ;
        RECT 67.700 211.325 68.150 211.785 ;
        RECT 68.425 211.615 68.705 212.285 ;
        RECT 69.490 212.205 70.660 212.375 ;
        RECT 69.335 211.825 69.980 212.035 ;
        RECT 70.150 211.825 70.720 212.035 ;
        RECT 70.890 211.655 71.060 212.855 ;
        RECT 71.600 212.455 71.770 212.660 ;
        RECT 67.025 211.105 68.150 211.325 ;
        RECT 67.025 210.645 67.305 211.105 ;
        RECT 67.825 210.475 68.150 210.935 ;
        RECT 68.320 210.645 68.705 211.615 ;
        RECT 68.875 210.475 69.165 211.640 ;
        RECT 69.550 210.475 69.880 211.575 ;
        RECT 70.355 211.245 71.060 211.655 ;
        RECT 71.230 212.285 71.770 212.455 ;
        RECT 72.050 212.285 72.220 213.025 ;
        RECT 72.485 212.285 72.845 212.660 ;
        RECT 73.105 212.475 73.275 212.765 ;
        RECT 73.445 212.645 73.775 213.025 ;
        RECT 73.105 212.305 73.770 212.475 ;
        RECT 71.230 211.585 71.400 212.285 ;
        RECT 71.570 211.785 71.900 212.115 ;
        RECT 72.070 211.785 72.420 212.115 ;
        RECT 71.230 211.415 71.855 211.585 ;
        RECT 72.070 211.245 72.335 211.785 ;
        RECT 72.590 211.630 72.845 212.285 ;
        RECT 70.355 211.075 72.335 211.245 ;
        RECT 70.355 210.645 70.680 211.075 ;
        RECT 70.850 210.475 71.180 210.895 ;
        RECT 71.925 210.475 72.335 210.905 ;
        RECT 72.505 210.645 72.845 211.630 ;
        RECT 73.020 211.485 73.370 212.135 ;
        RECT 73.540 211.315 73.770 212.305 ;
        RECT 73.105 211.145 73.770 211.315 ;
        RECT 73.105 210.645 73.275 211.145 ;
        RECT 73.445 210.475 73.775 210.975 ;
        RECT 73.945 210.645 74.130 212.765 ;
        RECT 74.385 212.565 74.635 213.025 ;
        RECT 74.805 212.575 75.140 212.745 ;
        RECT 75.335 212.575 76.010 212.745 ;
        RECT 74.805 212.435 74.975 212.575 ;
        RECT 74.300 211.445 74.580 212.395 ;
        RECT 74.750 212.305 74.975 212.435 ;
        RECT 74.750 211.200 74.920 212.305 ;
        RECT 75.145 212.155 75.670 212.375 ;
        RECT 75.090 211.390 75.330 211.985 ;
        RECT 75.500 211.455 75.670 212.155 ;
        RECT 75.840 211.795 76.010 212.575 ;
        RECT 76.330 212.525 76.700 213.025 ;
        RECT 76.880 212.575 77.285 212.745 ;
        RECT 77.455 212.575 78.240 212.745 ;
        RECT 76.880 212.345 77.050 212.575 ;
        RECT 76.220 212.045 77.050 212.345 ;
        RECT 77.435 212.075 77.900 212.405 ;
        RECT 76.220 212.015 76.420 212.045 ;
        RECT 76.540 211.795 76.710 211.865 ;
        RECT 75.840 211.625 76.710 211.795 ;
        RECT 76.200 211.535 76.710 211.625 ;
        RECT 74.750 211.070 75.055 211.200 ;
        RECT 75.500 211.090 76.030 211.455 ;
        RECT 74.370 210.475 74.635 210.935 ;
        RECT 74.805 210.645 75.055 211.070 ;
        RECT 76.200 210.920 76.370 211.535 ;
        RECT 75.265 210.750 76.370 210.920 ;
        RECT 76.540 210.475 76.710 211.275 ;
        RECT 76.880 210.975 77.050 212.045 ;
        RECT 77.220 211.145 77.410 211.865 ;
        RECT 77.580 211.115 77.900 212.075 ;
        RECT 78.070 212.115 78.240 212.575 ;
        RECT 78.515 212.495 78.725 213.025 ;
        RECT 78.985 212.285 79.315 212.810 ;
        RECT 79.485 212.415 79.655 213.025 ;
        RECT 79.825 212.370 80.155 212.805 ;
        RECT 80.465 212.475 80.635 212.765 ;
        RECT 80.805 212.645 81.135 213.025 ;
        RECT 79.825 212.285 80.205 212.370 ;
        RECT 80.465 212.305 81.130 212.475 ;
        RECT 79.115 212.115 79.315 212.285 ;
        RECT 79.980 212.245 80.205 212.285 ;
        RECT 78.070 211.785 78.945 212.115 ;
        RECT 79.115 211.785 79.865 212.115 ;
        RECT 76.880 210.645 77.130 210.975 ;
        RECT 78.070 210.945 78.240 211.785 ;
        RECT 79.115 211.580 79.305 211.785 ;
        RECT 80.035 211.665 80.205 212.245 ;
        RECT 79.990 211.615 80.205 211.665 ;
        RECT 78.410 211.205 79.305 211.580 ;
        RECT 79.815 211.535 80.205 211.615 ;
        RECT 77.355 210.775 78.240 210.945 ;
        RECT 78.420 210.475 78.735 210.975 ;
        RECT 78.965 210.645 79.305 211.205 ;
        RECT 79.475 210.475 79.645 211.485 ;
        RECT 79.815 210.690 80.145 211.535 ;
        RECT 80.380 211.485 80.730 212.135 ;
        RECT 80.900 211.315 81.130 212.305 ;
        RECT 80.465 211.145 81.130 211.315 ;
        RECT 80.465 210.645 80.635 211.145 ;
        RECT 80.805 210.475 81.135 210.975 ;
        RECT 81.305 210.645 81.490 212.765 ;
        RECT 81.745 212.565 81.995 213.025 ;
        RECT 82.165 212.575 82.500 212.745 ;
        RECT 82.695 212.575 83.370 212.745 ;
        RECT 82.165 212.435 82.335 212.575 ;
        RECT 81.660 211.445 81.940 212.395 ;
        RECT 82.110 212.305 82.335 212.435 ;
        RECT 82.110 211.200 82.280 212.305 ;
        RECT 82.505 212.155 83.030 212.375 ;
        RECT 82.450 211.390 82.690 211.985 ;
        RECT 82.860 211.455 83.030 212.155 ;
        RECT 83.200 211.795 83.370 212.575 ;
        RECT 83.690 212.525 84.060 213.025 ;
        RECT 84.240 212.575 84.645 212.745 ;
        RECT 84.815 212.575 85.600 212.745 ;
        RECT 84.240 212.345 84.410 212.575 ;
        RECT 83.580 212.045 84.410 212.345 ;
        RECT 84.795 212.075 85.260 212.405 ;
        RECT 83.580 212.015 83.780 212.045 ;
        RECT 83.900 211.795 84.070 211.865 ;
        RECT 83.200 211.625 84.070 211.795 ;
        RECT 83.560 211.535 84.070 211.625 ;
        RECT 82.110 211.070 82.415 211.200 ;
        RECT 82.860 211.090 83.390 211.455 ;
        RECT 81.730 210.475 81.995 210.935 ;
        RECT 82.165 210.645 82.415 211.070 ;
        RECT 83.560 210.920 83.730 211.535 ;
        RECT 82.625 210.750 83.730 210.920 ;
        RECT 83.900 210.475 84.070 211.275 ;
        RECT 84.240 210.975 84.410 212.045 ;
        RECT 84.580 211.145 84.770 211.865 ;
        RECT 84.940 211.115 85.260 212.075 ;
        RECT 85.430 212.115 85.600 212.575 ;
        RECT 85.875 212.495 86.085 213.025 ;
        RECT 86.345 212.285 86.675 212.810 ;
        RECT 86.845 212.415 87.015 213.025 ;
        RECT 87.185 212.370 87.515 212.805 ;
        RECT 88.745 212.375 88.915 212.855 ;
        RECT 89.085 212.545 89.415 213.025 ;
        RECT 89.640 212.605 91.175 212.855 ;
        RECT 89.640 212.375 89.810 212.605 ;
        RECT 87.185 212.285 87.565 212.370 ;
        RECT 86.475 212.115 86.675 212.285 ;
        RECT 87.340 212.245 87.565 212.285 ;
        RECT 85.430 211.785 86.305 212.115 ;
        RECT 86.475 211.785 87.225 212.115 ;
        RECT 84.240 210.645 84.490 210.975 ;
        RECT 85.430 210.945 85.600 211.785 ;
        RECT 86.475 211.580 86.665 211.785 ;
        RECT 87.395 211.665 87.565 212.245 ;
        RECT 88.745 212.205 89.810 212.375 ;
        RECT 89.990 212.035 90.270 212.435 ;
        RECT 88.660 211.825 89.010 212.035 ;
        RECT 89.180 211.835 89.625 212.035 ;
        RECT 89.795 211.835 90.270 212.035 ;
        RECT 90.540 212.035 90.825 212.435 ;
        RECT 91.005 212.375 91.175 212.605 ;
        RECT 91.345 212.545 91.675 213.025 ;
        RECT 91.890 212.525 92.145 212.855 ;
        RECT 91.935 212.515 92.145 212.525 ;
        RECT 91.960 212.445 92.145 212.515 ;
        RECT 91.005 212.205 91.805 212.375 ;
        RECT 90.540 211.835 90.870 212.035 ;
        RECT 91.040 211.835 91.405 212.035 ;
        RECT 87.350 211.615 87.565 211.665 ;
        RECT 91.635 211.655 91.805 212.205 ;
        RECT 85.770 211.205 86.665 211.580 ;
        RECT 87.175 211.535 87.565 211.615 ;
        RECT 84.715 210.775 85.600 210.945 ;
        RECT 85.780 210.475 86.095 210.975 ;
        RECT 86.325 210.645 86.665 211.205 ;
        RECT 86.835 210.475 87.005 211.485 ;
        RECT 87.175 210.690 87.505 211.535 ;
        RECT 88.745 211.485 91.805 211.655 ;
        RECT 88.745 210.645 88.915 211.485 ;
        RECT 91.975 211.315 92.145 212.445 ;
        RECT 92.395 212.205 92.605 213.025 ;
        RECT 92.775 212.225 93.105 212.855 ;
        RECT 92.775 211.625 93.025 212.225 ;
        RECT 93.275 212.205 93.505 213.025 ;
        RECT 94.635 212.300 94.925 213.025 ;
        RECT 95.110 212.455 95.365 212.805 ;
        RECT 95.535 212.625 95.865 213.025 ;
        RECT 96.035 212.455 96.205 212.805 ;
        RECT 96.375 212.625 96.755 213.025 ;
        RECT 95.110 212.285 96.775 212.455 ;
        RECT 96.945 212.350 97.220 212.695 ;
        RECT 96.605 212.115 96.775 212.285 ;
        RECT 93.195 211.785 93.525 212.035 ;
        RECT 95.095 211.785 95.440 212.115 ;
        RECT 95.610 211.785 96.435 212.115 ;
        RECT 96.605 211.785 96.880 212.115 ;
        RECT 89.085 210.815 89.415 211.315 ;
        RECT 89.585 211.075 91.220 211.315 ;
        RECT 89.585 210.985 89.815 211.075 ;
        RECT 89.925 210.815 90.255 210.855 ;
        RECT 89.085 210.645 90.255 210.815 ;
        RECT 90.445 210.475 90.800 210.895 ;
        RECT 90.970 210.645 91.220 211.075 ;
        RECT 91.390 210.475 91.720 211.235 ;
        RECT 91.890 210.645 92.145 211.315 ;
        RECT 92.395 210.475 92.605 211.615 ;
        RECT 92.775 210.645 93.105 211.625 ;
        RECT 93.275 210.475 93.505 211.615 ;
        RECT 94.635 210.475 94.925 211.640 ;
        RECT 95.115 211.325 95.440 211.615 ;
        RECT 95.610 211.495 95.805 211.785 ;
        RECT 96.605 211.615 96.775 211.785 ;
        RECT 97.050 211.615 97.220 212.350 ;
        RECT 96.115 211.445 96.775 211.615 ;
        RECT 96.115 211.325 96.285 211.445 ;
        RECT 95.115 211.155 96.285 211.325 ;
        RECT 95.095 210.695 96.285 210.985 ;
        RECT 96.455 210.475 96.735 211.275 ;
        RECT 96.945 210.645 97.220 211.615 ;
        RECT 97.395 212.300 97.655 212.855 ;
        RECT 97.825 212.580 98.255 213.025 ;
        RECT 98.490 212.455 98.660 212.855 ;
        RECT 98.830 212.625 99.550 213.025 ;
        RECT 97.395 211.585 97.570 212.300 ;
        RECT 98.490 212.285 99.370 212.455 ;
        RECT 99.720 212.410 99.890 212.855 ;
        RECT 100.465 212.515 100.865 213.025 ;
        RECT 97.740 211.785 97.995 212.115 ;
        RECT 97.395 210.645 97.655 211.585 ;
        RECT 97.825 211.305 97.995 211.785 ;
        RECT 98.220 211.495 98.550 212.115 ;
        RECT 98.720 211.735 99.010 212.115 ;
        RECT 99.200 211.565 99.370 212.285 ;
        RECT 98.850 211.395 99.370 211.565 ;
        RECT 99.540 212.240 99.890 212.410 ;
        RECT 101.125 212.370 101.455 212.805 ;
        RECT 101.625 212.415 101.795 213.025 ;
        RECT 97.825 211.135 98.585 211.305 ;
        RECT 98.850 211.205 99.020 211.395 ;
        RECT 99.540 211.215 99.710 212.240 ;
        RECT 100.130 211.755 100.390 212.345 ;
        RECT 99.910 211.455 100.390 211.755 ;
        RECT 100.590 211.455 100.850 212.345 ;
        RECT 101.075 212.285 101.455 212.370 ;
        RECT 101.965 212.285 102.295 212.810 ;
        RECT 102.555 212.495 102.765 213.025 ;
        RECT 103.040 212.575 103.825 212.745 ;
        RECT 103.995 212.575 104.400 212.745 ;
        RECT 101.075 212.245 101.300 212.285 ;
        RECT 101.075 211.665 101.245 212.245 ;
        RECT 101.965 212.115 102.165 212.285 ;
        RECT 103.040 212.115 103.210 212.575 ;
        RECT 101.415 211.785 102.165 212.115 ;
        RECT 102.335 211.785 103.210 212.115 ;
        RECT 101.075 211.615 101.290 211.665 ;
        RECT 101.075 211.535 101.465 211.615 ;
        RECT 98.415 210.910 98.585 211.135 ;
        RECT 99.300 211.045 99.710 211.215 ;
        RECT 99.885 211.105 100.825 211.275 ;
        RECT 99.300 210.910 99.555 211.045 ;
        RECT 97.825 210.475 98.155 210.875 ;
        RECT 98.415 210.740 99.555 210.910 ;
        RECT 99.885 210.855 100.055 211.105 ;
        RECT 99.300 210.645 99.555 210.740 ;
        RECT 99.725 210.685 100.055 210.855 ;
        RECT 100.225 210.475 100.475 210.935 ;
        RECT 100.645 210.645 100.825 211.105 ;
        RECT 101.135 210.690 101.465 211.535 ;
        RECT 101.975 211.580 102.165 211.785 ;
        RECT 101.635 210.475 101.805 211.485 ;
        RECT 101.975 211.205 102.870 211.580 ;
        RECT 101.975 210.645 102.315 211.205 ;
        RECT 102.545 210.475 102.860 210.975 ;
        RECT 103.040 210.945 103.210 211.785 ;
        RECT 103.380 212.075 103.845 212.405 ;
        RECT 104.230 212.345 104.400 212.575 ;
        RECT 104.580 212.525 104.950 213.025 ;
        RECT 105.270 212.575 105.945 212.745 ;
        RECT 106.140 212.575 106.475 212.745 ;
        RECT 103.380 211.115 103.700 212.075 ;
        RECT 104.230 212.045 105.060 212.345 ;
        RECT 103.870 211.145 104.060 211.865 ;
        RECT 104.230 210.975 104.400 212.045 ;
        RECT 104.860 212.015 105.060 212.045 ;
        RECT 104.570 211.795 104.740 211.865 ;
        RECT 105.270 211.795 105.440 212.575 ;
        RECT 106.305 212.435 106.475 212.575 ;
        RECT 106.645 212.565 106.895 213.025 ;
        RECT 104.570 211.625 105.440 211.795 ;
        RECT 105.610 212.155 106.135 212.375 ;
        RECT 106.305 212.305 106.530 212.435 ;
        RECT 104.570 211.535 105.080 211.625 ;
        RECT 103.040 210.775 103.925 210.945 ;
        RECT 104.150 210.645 104.400 210.975 ;
        RECT 104.570 210.475 104.740 211.275 ;
        RECT 104.910 210.920 105.080 211.535 ;
        RECT 105.610 211.455 105.780 212.155 ;
        RECT 105.250 211.090 105.780 211.455 ;
        RECT 105.950 211.390 106.190 211.985 ;
        RECT 106.360 211.200 106.530 212.305 ;
        RECT 106.700 211.445 106.980 212.395 ;
        RECT 106.225 211.070 106.530 211.200 ;
        RECT 104.910 210.750 106.015 210.920 ;
        RECT 106.225 210.645 106.475 211.070 ;
        RECT 106.645 210.475 106.910 210.935 ;
        RECT 107.150 210.645 107.335 212.765 ;
        RECT 107.505 212.645 107.835 213.025 ;
        RECT 108.005 212.475 108.175 212.765 ;
        RECT 108.435 212.480 113.780 213.025 ;
        RECT 113.955 212.480 119.300 213.025 ;
        RECT 107.510 212.305 108.175 212.475 ;
        RECT 107.510 211.315 107.740 212.305 ;
        RECT 107.910 211.485 108.260 212.135 ;
        RECT 110.020 211.650 110.360 212.480 ;
        RECT 107.510 211.145 108.175 211.315 ;
        RECT 107.505 210.475 107.835 210.975 ;
        RECT 108.005 210.645 108.175 211.145 ;
        RECT 111.840 210.910 112.190 212.160 ;
        RECT 115.540 211.650 115.880 212.480 ;
        RECT 120.395 212.300 120.685 213.025 ;
        RECT 120.855 212.480 126.200 213.025 ;
        RECT 126.375 212.480 131.720 213.025 ;
        RECT 131.895 212.480 137.240 213.025 ;
        RECT 137.415 212.480 142.760 213.025 ;
        RECT 117.360 210.910 117.710 212.160 ;
        RECT 122.440 211.650 122.780 212.480 ;
        RECT 108.435 210.475 113.780 210.910 ;
        RECT 113.955 210.475 119.300 210.910 ;
        RECT 120.395 210.475 120.685 211.640 ;
        RECT 124.260 210.910 124.610 212.160 ;
        RECT 127.960 211.650 128.300 212.480 ;
        RECT 129.780 210.910 130.130 212.160 ;
        RECT 133.480 211.650 133.820 212.480 ;
        RECT 135.300 210.910 135.650 212.160 ;
        RECT 139.000 211.650 139.340 212.480 ;
        RECT 142.935 212.255 145.525 213.025 ;
        RECT 145.695 212.275 146.905 213.025 ;
        RECT 140.820 210.910 141.170 212.160 ;
        RECT 142.935 211.735 144.145 212.255 ;
        RECT 144.315 211.565 145.525 212.085 ;
        RECT 120.855 210.475 126.200 210.910 ;
        RECT 126.375 210.475 131.720 210.910 ;
        RECT 131.895 210.475 137.240 210.910 ;
        RECT 137.415 210.475 142.760 210.910 ;
        RECT 142.935 210.475 145.525 211.565 ;
        RECT 145.695 211.565 146.215 212.105 ;
        RECT 146.385 211.735 146.905 212.275 ;
        RECT 145.695 210.475 146.905 211.565 ;
        RECT 17.270 210.305 146.990 210.475 ;
        RECT 17.355 209.215 18.565 210.305 ;
        RECT 18.735 209.870 24.080 210.305 ;
        RECT 24.255 209.870 29.600 210.305 ;
        RECT 17.355 208.505 17.875 209.045 ;
        RECT 18.045 208.675 18.565 209.215 ;
        RECT 17.355 207.755 18.565 208.505 ;
        RECT 20.320 208.300 20.660 209.130 ;
        RECT 22.140 208.620 22.490 209.870 ;
        RECT 25.840 208.300 26.180 209.130 ;
        RECT 27.660 208.620 28.010 209.870 ;
        RECT 30.235 209.140 30.525 210.305 ;
        RECT 30.695 209.870 36.040 210.305 ;
        RECT 36.215 209.870 41.560 210.305 ;
        RECT 18.735 207.755 24.080 208.300 ;
        RECT 24.255 207.755 29.600 208.300 ;
        RECT 30.235 207.755 30.525 208.480 ;
        RECT 32.280 208.300 32.620 209.130 ;
        RECT 34.100 208.620 34.450 209.870 ;
        RECT 37.800 208.300 38.140 209.130 ;
        RECT 39.620 208.620 39.970 209.870 ;
        RECT 41.735 209.215 45.245 210.305 ;
        RECT 45.965 209.635 46.135 210.135 ;
        RECT 46.305 209.805 46.635 210.305 ;
        RECT 45.965 209.465 46.630 209.635 ;
        RECT 41.735 208.525 43.385 209.045 ;
        RECT 43.555 208.695 45.245 209.215 ;
        RECT 45.880 208.645 46.230 209.295 ;
        RECT 30.695 207.755 36.040 208.300 ;
        RECT 36.215 207.755 41.560 208.300 ;
        RECT 41.735 207.755 45.245 208.525 ;
        RECT 46.400 208.475 46.630 209.465 ;
        RECT 45.965 208.305 46.630 208.475 ;
        RECT 45.965 208.015 46.135 208.305 ;
        RECT 46.305 207.755 46.635 208.135 ;
        RECT 46.805 208.015 46.990 210.135 ;
        RECT 47.230 209.845 47.495 210.305 ;
        RECT 47.665 209.710 47.915 210.135 ;
        RECT 48.125 209.860 49.230 210.030 ;
        RECT 47.610 209.580 47.915 209.710 ;
        RECT 47.160 208.385 47.440 209.335 ;
        RECT 47.610 208.475 47.780 209.580 ;
        RECT 47.950 208.795 48.190 209.390 ;
        RECT 48.360 209.325 48.890 209.690 ;
        RECT 48.360 208.625 48.530 209.325 ;
        RECT 49.060 209.245 49.230 209.860 ;
        RECT 49.400 209.505 49.570 210.305 ;
        RECT 49.740 209.805 49.990 210.135 ;
        RECT 50.215 209.835 51.100 210.005 ;
        RECT 49.060 209.155 49.570 209.245 ;
        RECT 47.610 208.345 47.835 208.475 ;
        RECT 48.005 208.405 48.530 208.625 ;
        RECT 48.700 208.985 49.570 209.155 ;
        RECT 47.245 207.755 47.495 208.215 ;
        RECT 47.665 208.205 47.835 208.345 ;
        RECT 48.700 208.205 48.870 208.985 ;
        RECT 49.400 208.915 49.570 208.985 ;
        RECT 49.080 208.735 49.280 208.765 ;
        RECT 49.740 208.735 49.910 209.805 ;
        RECT 50.080 208.915 50.270 209.635 ;
        RECT 49.080 208.435 49.910 208.735 ;
        RECT 50.440 208.705 50.760 209.665 ;
        RECT 47.665 208.035 48.000 208.205 ;
        RECT 48.195 208.035 48.870 208.205 ;
        RECT 49.190 207.755 49.560 208.255 ;
        RECT 49.740 208.205 49.910 208.435 ;
        RECT 50.295 208.375 50.760 208.705 ;
        RECT 50.930 208.995 51.100 209.835 ;
        RECT 51.280 209.805 51.595 210.305 ;
        RECT 51.825 209.575 52.165 210.135 ;
        RECT 51.270 209.200 52.165 209.575 ;
        RECT 52.335 209.295 52.505 210.305 ;
        RECT 51.975 208.995 52.165 209.200 ;
        RECT 52.675 209.245 53.005 210.090 ;
        RECT 54.165 209.695 54.495 210.125 ;
        RECT 54.675 209.865 54.870 210.305 ;
        RECT 55.040 209.695 55.370 210.125 ;
        RECT 54.165 209.525 55.370 209.695 ;
        RECT 52.675 209.165 53.065 209.245 ;
        RECT 54.165 209.195 55.060 209.525 ;
        RECT 55.540 209.355 55.815 210.125 ;
        RECT 52.850 209.115 53.065 209.165 ;
        RECT 50.930 208.665 51.805 208.995 ;
        RECT 51.975 208.665 52.725 208.995 ;
        RECT 50.930 208.205 51.100 208.665 ;
        RECT 51.975 208.495 52.175 208.665 ;
        RECT 52.895 208.535 53.065 209.115 ;
        RECT 55.230 209.165 55.815 209.355 ;
        RECT 54.170 208.665 54.465 208.995 ;
        RECT 54.645 208.665 55.060 208.995 ;
        RECT 52.840 208.495 53.065 208.535 ;
        RECT 49.740 208.035 50.145 208.205 ;
        RECT 50.315 208.035 51.100 208.205 ;
        RECT 51.375 207.755 51.585 208.285 ;
        RECT 51.845 207.970 52.175 208.495 ;
        RECT 52.685 208.410 53.065 208.495 ;
        RECT 52.345 207.755 52.515 208.365 ;
        RECT 52.685 207.975 53.015 208.410 ;
        RECT 54.165 207.755 54.465 208.485 ;
        RECT 54.645 208.045 54.875 208.665 ;
        RECT 55.230 208.495 55.405 209.165 ;
        RECT 55.995 209.140 56.285 210.305 ;
        RECT 56.460 209.925 56.795 210.305 ;
        RECT 55.075 208.315 55.405 208.495 ;
        RECT 55.575 208.345 55.815 208.995 ;
        RECT 55.075 207.935 55.300 208.315 ;
        RECT 55.470 207.755 55.800 208.145 ;
        RECT 55.995 207.755 56.285 208.480 ;
        RECT 56.455 208.435 56.695 209.745 ;
        RECT 56.965 209.335 57.215 210.135 ;
        RECT 57.435 209.585 57.765 210.305 ;
        RECT 57.950 209.335 58.200 210.135 ;
        RECT 58.665 209.505 58.995 210.305 ;
        RECT 59.165 209.875 59.505 210.135 ;
        RECT 56.865 209.165 59.055 209.335 ;
        RECT 56.865 208.255 57.035 209.165 ;
        RECT 58.740 208.995 59.055 209.165 ;
        RECT 56.540 207.925 57.035 208.255 ;
        RECT 57.255 208.030 57.605 208.995 ;
        RECT 57.785 208.025 58.085 208.995 ;
        RECT 58.265 208.025 58.545 208.995 ;
        RECT 58.740 208.745 59.070 208.995 ;
        RECT 58.725 207.755 58.995 208.555 ;
        RECT 59.245 208.475 59.505 209.875 ;
        RECT 59.165 207.965 59.505 208.475 ;
        RECT 60.135 209.435 60.410 210.135 ;
        RECT 60.580 209.760 60.835 210.305 ;
        RECT 61.005 209.795 61.485 210.135 ;
        RECT 61.660 209.750 62.265 210.305 ;
        RECT 62.435 209.795 62.735 210.305 ;
        RECT 61.650 209.650 62.265 209.750 ;
        RECT 61.650 209.625 61.835 209.650 ;
        RECT 62.905 209.625 63.235 210.135 ;
        RECT 63.405 209.795 64.035 210.305 ;
        RECT 64.615 209.795 64.995 209.965 ;
        RECT 65.165 209.795 65.465 210.305 ;
        RECT 64.825 209.625 64.995 209.795 ;
        RECT 65.745 209.635 65.915 210.135 ;
        RECT 66.085 209.805 66.415 210.305 ;
        RECT 60.135 208.405 60.305 209.435 ;
        RECT 60.580 209.305 61.335 209.555 ;
        RECT 61.505 209.380 61.835 209.625 ;
        RECT 60.580 209.270 61.350 209.305 ;
        RECT 60.580 209.260 61.365 209.270 ;
        RECT 60.475 209.245 61.370 209.260 ;
        RECT 60.475 209.230 61.390 209.245 ;
        RECT 60.475 209.220 61.410 209.230 ;
        RECT 60.475 209.210 61.435 209.220 ;
        RECT 60.475 209.180 61.505 209.210 ;
        RECT 60.475 209.150 61.525 209.180 ;
        RECT 60.475 209.120 61.545 209.150 ;
        RECT 60.475 209.095 61.575 209.120 ;
        RECT 60.475 209.060 61.610 209.095 ;
        RECT 60.475 209.055 61.640 209.060 ;
        RECT 60.475 208.660 60.705 209.055 ;
        RECT 61.250 209.050 61.640 209.055 ;
        RECT 61.275 209.040 61.640 209.050 ;
        RECT 61.290 209.035 61.640 209.040 ;
        RECT 61.305 209.030 61.640 209.035 ;
        RECT 62.005 209.030 62.265 209.480 ;
        RECT 61.305 209.025 62.265 209.030 ;
        RECT 61.315 209.015 62.265 209.025 ;
        RECT 61.325 209.010 62.265 209.015 ;
        RECT 61.335 209.000 62.265 209.010 ;
        RECT 61.340 208.990 62.265 209.000 ;
        RECT 61.345 208.985 62.265 208.990 ;
        RECT 61.355 208.970 62.265 208.985 ;
        RECT 61.360 208.955 62.265 208.970 ;
        RECT 61.370 208.930 62.265 208.955 ;
        RECT 60.875 208.460 61.205 208.885 ;
        RECT 60.135 207.925 60.395 208.405 ;
        RECT 60.565 207.755 60.815 208.295 ;
        RECT 60.985 207.975 61.205 208.460 ;
        RECT 61.375 208.860 62.265 208.930 ;
        RECT 62.435 209.455 64.655 209.625 ;
        RECT 61.375 208.135 61.545 208.860 ;
        RECT 61.715 208.305 62.265 208.690 ;
        RECT 62.435 208.495 62.605 209.455 ;
        RECT 62.775 209.115 64.315 209.285 ;
        RECT 62.775 208.665 63.020 209.115 ;
        RECT 63.280 208.745 63.975 208.945 ;
        RECT 64.145 208.915 64.315 209.115 ;
        RECT 64.485 209.255 64.655 209.455 ;
        RECT 64.825 209.425 65.485 209.625 ;
        RECT 65.745 209.465 66.410 209.635 ;
        RECT 64.485 209.085 65.145 209.255 ;
        RECT 64.145 208.745 64.745 208.915 ;
        RECT 64.975 208.665 65.145 209.085 ;
        RECT 61.375 207.965 62.265 208.135 ;
        RECT 62.435 207.950 62.900 208.495 ;
        RECT 63.405 207.755 63.575 208.575 ;
        RECT 63.745 208.495 64.655 208.575 ;
        RECT 65.315 208.495 65.485 209.425 ;
        RECT 65.660 208.645 66.010 209.295 ;
        RECT 63.745 208.405 64.995 208.495 ;
        RECT 63.745 207.925 64.075 208.405 ;
        RECT 64.485 208.325 64.995 208.405 ;
        RECT 64.245 207.755 64.595 208.145 ;
        RECT 64.765 207.925 64.995 208.325 ;
        RECT 65.165 208.015 65.485 208.495 ;
        RECT 66.180 208.475 66.410 209.465 ;
        RECT 65.745 208.305 66.410 208.475 ;
        RECT 65.745 208.015 65.915 208.305 ;
        RECT 66.085 207.755 66.415 208.135 ;
        RECT 66.585 208.015 66.770 210.135 ;
        RECT 67.010 209.845 67.275 210.305 ;
        RECT 67.445 209.710 67.695 210.135 ;
        RECT 67.905 209.860 69.010 210.030 ;
        RECT 67.390 209.580 67.695 209.710 ;
        RECT 66.940 208.385 67.220 209.335 ;
        RECT 67.390 208.475 67.560 209.580 ;
        RECT 67.730 208.795 67.970 209.390 ;
        RECT 68.140 209.325 68.670 209.690 ;
        RECT 68.140 208.625 68.310 209.325 ;
        RECT 68.840 209.245 69.010 209.860 ;
        RECT 69.180 209.505 69.350 210.305 ;
        RECT 69.520 209.805 69.770 210.135 ;
        RECT 69.995 209.835 70.880 210.005 ;
        RECT 68.840 209.155 69.350 209.245 ;
        RECT 67.390 208.345 67.615 208.475 ;
        RECT 67.785 208.405 68.310 208.625 ;
        RECT 68.480 208.985 69.350 209.155 ;
        RECT 67.025 207.755 67.275 208.215 ;
        RECT 67.445 208.205 67.615 208.345 ;
        RECT 68.480 208.205 68.650 208.985 ;
        RECT 69.180 208.915 69.350 208.985 ;
        RECT 68.860 208.735 69.060 208.765 ;
        RECT 69.520 208.735 69.690 209.805 ;
        RECT 69.860 208.915 70.050 209.635 ;
        RECT 68.860 208.435 69.690 208.735 ;
        RECT 70.220 208.705 70.540 209.665 ;
        RECT 67.445 208.035 67.780 208.205 ;
        RECT 67.975 208.035 68.650 208.205 ;
        RECT 68.970 207.755 69.340 208.255 ;
        RECT 69.520 208.205 69.690 208.435 ;
        RECT 70.075 208.375 70.540 208.705 ;
        RECT 70.710 208.995 70.880 209.835 ;
        RECT 71.060 209.805 71.375 210.305 ;
        RECT 71.605 209.575 71.945 210.135 ;
        RECT 71.050 209.200 71.945 209.575 ;
        RECT 72.115 209.295 72.285 210.305 ;
        RECT 71.755 208.995 71.945 209.200 ;
        RECT 72.455 209.245 72.785 210.090 ;
        RECT 73.015 209.795 74.205 210.085 ;
        RECT 73.035 209.455 74.205 209.625 ;
        RECT 74.375 209.505 74.655 210.305 ;
        RECT 72.455 209.165 72.845 209.245 ;
        RECT 73.035 209.165 73.360 209.455 ;
        RECT 74.035 209.335 74.205 209.455 ;
        RECT 72.630 209.115 72.845 209.165 ;
        RECT 70.710 208.665 71.585 208.995 ;
        RECT 71.755 208.665 72.505 208.995 ;
        RECT 70.710 208.205 70.880 208.665 ;
        RECT 71.755 208.495 71.955 208.665 ;
        RECT 72.675 208.535 72.845 209.115 ;
        RECT 73.530 208.995 73.725 209.285 ;
        RECT 74.035 209.165 74.695 209.335 ;
        RECT 74.865 209.165 75.140 210.135 ;
        RECT 75.315 209.870 80.660 210.305 ;
        RECT 74.525 208.995 74.695 209.165 ;
        RECT 73.015 208.665 73.360 208.995 ;
        RECT 73.530 208.665 74.355 208.995 ;
        RECT 74.525 208.665 74.800 208.995 ;
        RECT 72.620 208.495 72.845 208.535 ;
        RECT 74.525 208.495 74.695 208.665 ;
        RECT 69.520 208.035 69.925 208.205 ;
        RECT 70.095 208.035 70.880 208.205 ;
        RECT 71.155 207.755 71.365 208.285 ;
        RECT 71.625 207.970 71.955 208.495 ;
        RECT 72.465 208.410 72.845 208.495 ;
        RECT 72.125 207.755 72.295 208.365 ;
        RECT 72.465 207.975 72.795 208.410 ;
        RECT 73.030 208.325 74.695 208.495 ;
        RECT 74.970 208.430 75.140 209.165 ;
        RECT 73.030 207.975 73.285 208.325 ;
        RECT 73.455 207.755 73.785 208.155 ;
        RECT 73.955 207.975 74.125 208.325 ;
        RECT 74.295 207.755 74.675 208.155 ;
        RECT 74.865 208.085 75.140 208.430 ;
        RECT 76.900 208.300 77.240 209.130 ;
        RECT 78.720 208.620 79.070 209.870 ;
        RECT 81.755 209.140 82.045 210.305 ;
        RECT 75.315 207.755 80.660 208.300 ;
        RECT 81.755 207.755 82.045 208.480 ;
        RECT 82.690 207.935 82.970 210.125 ;
        RECT 83.160 209.165 83.445 210.305 ;
        RECT 83.710 209.655 83.880 210.125 ;
        RECT 84.055 209.825 84.385 210.305 ;
        RECT 84.555 209.655 84.735 210.125 ;
        RECT 83.710 209.455 84.735 209.655 ;
        RECT 83.170 208.485 83.430 208.995 ;
        RECT 83.640 208.665 83.900 209.285 ;
        RECT 84.095 208.665 84.520 209.285 ;
        RECT 84.905 209.015 85.235 210.125 ;
        RECT 85.405 209.895 85.755 210.305 ;
        RECT 85.925 209.715 86.165 210.105 ;
        RECT 84.690 208.715 85.235 209.015 ;
        RECT 85.415 209.515 86.165 209.715 ;
        RECT 85.415 208.835 85.755 209.515 ;
        RECT 84.690 208.485 84.910 208.715 ;
        RECT 83.170 208.295 84.910 208.485 ;
        RECT 83.170 207.755 83.900 208.125 ;
        RECT 84.480 207.935 84.910 208.295 ;
        RECT 85.080 207.755 85.325 208.535 ;
        RECT 85.525 207.935 85.755 208.835 ;
        RECT 85.935 207.995 86.165 209.335 ;
        RECT 86.355 209.165 86.740 210.135 ;
        RECT 86.910 209.845 87.235 210.305 ;
        RECT 87.755 209.675 88.035 210.135 ;
        RECT 86.910 209.455 88.035 209.675 ;
        RECT 86.355 208.495 86.635 209.165 ;
        RECT 86.910 208.995 87.360 209.455 ;
        RECT 88.225 209.285 88.625 210.135 ;
        RECT 89.025 209.845 89.295 210.305 ;
        RECT 89.465 209.675 89.750 210.135 ;
        RECT 86.805 208.665 87.360 208.995 ;
        RECT 87.530 208.725 88.625 209.285 ;
        RECT 86.910 208.555 87.360 208.665 ;
        RECT 86.355 207.925 86.740 208.495 ;
        RECT 86.910 208.385 88.035 208.555 ;
        RECT 86.910 207.755 87.235 208.215 ;
        RECT 87.755 207.925 88.035 208.385 ;
        RECT 88.225 207.925 88.625 208.725 ;
        RECT 88.795 209.455 89.750 209.675 ;
        RECT 88.795 208.555 89.005 209.455 ;
        RECT 89.175 208.725 89.865 209.285 ;
        RECT 90.035 209.165 90.310 210.135 ;
        RECT 90.520 209.505 90.800 210.305 ;
        RECT 90.970 209.795 92.585 210.125 ;
        RECT 90.970 209.455 92.145 209.625 ;
        RECT 90.970 209.335 91.140 209.455 ;
        RECT 90.480 209.165 91.140 209.335 ;
        RECT 88.795 208.385 89.750 208.555 ;
        RECT 89.025 207.755 89.295 208.215 ;
        RECT 89.465 207.925 89.750 208.385 ;
        RECT 90.035 208.430 90.205 209.165 ;
        RECT 90.480 208.995 90.650 209.165 ;
        RECT 91.400 208.995 91.645 209.285 ;
        RECT 91.815 209.165 92.145 209.455 ;
        RECT 92.405 208.995 92.575 209.555 ;
        RECT 92.825 209.165 93.085 210.305 ;
        RECT 93.440 209.335 93.830 209.510 ;
        RECT 94.315 209.505 94.645 210.305 ;
        RECT 94.815 209.515 95.350 210.135 ;
        RECT 93.440 209.165 94.865 209.335 ;
        RECT 90.375 208.665 90.650 208.995 ;
        RECT 90.820 208.665 91.645 208.995 ;
        RECT 91.860 208.665 92.575 208.995 ;
        RECT 92.745 208.745 93.080 208.995 ;
        RECT 90.480 208.495 90.650 208.665 ;
        RECT 92.325 208.575 92.575 208.665 ;
        RECT 90.035 208.085 90.310 208.430 ;
        RECT 90.480 208.325 92.145 208.495 ;
        RECT 90.500 207.755 90.875 208.155 ;
        RECT 91.045 207.975 91.215 208.325 ;
        RECT 91.385 207.755 91.715 208.155 ;
        RECT 91.885 207.925 92.145 208.325 ;
        RECT 92.325 208.155 92.655 208.575 ;
        RECT 92.825 207.755 93.085 208.575 ;
        RECT 93.315 208.435 93.670 208.995 ;
        RECT 93.840 208.265 94.010 209.165 ;
        RECT 94.180 208.435 94.445 208.995 ;
        RECT 94.695 208.665 94.865 209.165 ;
        RECT 95.035 208.495 95.350 209.515 ;
        RECT 95.555 209.215 97.225 210.305 ;
        RECT 93.420 207.755 93.660 208.265 ;
        RECT 93.840 207.935 94.120 208.265 ;
        RECT 94.350 207.755 94.565 208.265 ;
        RECT 94.735 207.925 95.350 208.495 ;
        RECT 95.555 208.525 96.305 209.045 ;
        RECT 96.475 208.695 97.225 209.215 ;
        RECT 97.395 209.335 97.685 210.135 ;
        RECT 97.855 209.505 98.090 210.305 ;
        RECT 98.275 209.965 99.810 210.135 ;
        RECT 98.275 209.335 98.605 209.965 ;
        RECT 97.395 209.165 98.605 209.335 ;
        RECT 97.395 208.665 97.640 208.995 ;
        RECT 95.555 207.755 97.225 208.525 ;
        RECT 97.810 208.495 97.980 209.165 ;
        RECT 98.775 208.995 99.010 209.740 ;
        RECT 98.150 208.665 98.550 208.995 ;
        RECT 98.720 208.665 99.010 208.995 ;
        RECT 99.200 208.995 99.470 209.740 ;
        RECT 99.640 209.335 99.810 209.965 ;
        RECT 99.980 209.505 100.385 210.305 ;
        RECT 99.640 209.165 100.385 209.335 ;
        RECT 99.200 208.665 99.540 208.995 ;
        RECT 99.710 208.665 100.045 208.995 ;
        RECT 100.215 208.665 100.385 209.165 ;
        RECT 100.555 208.740 100.905 210.135 ;
        RECT 101.075 209.870 106.420 210.305 ;
        RECT 97.395 207.925 97.980 208.495 ;
        RECT 98.230 208.325 99.625 208.495 ;
        RECT 98.230 207.980 98.560 208.325 ;
        RECT 98.775 207.755 99.150 208.155 ;
        RECT 99.330 207.980 99.625 208.325 ;
        RECT 99.795 207.755 100.465 208.495 ;
        RECT 100.635 207.925 100.905 208.740 ;
        RECT 102.660 208.300 103.000 209.130 ;
        RECT 104.480 208.620 104.830 209.870 ;
        RECT 107.515 209.140 107.805 210.305 ;
        RECT 107.975 209.870 113.320 210.305 ;
        RECT 113.495 209.870 118.840 210.305 ;
        RECT 119.015 209.870 124.360 210.305 ;
        RECT 124.535 209.870 129.880 210.305 ;
        RECT 101.075 207.755 106.420 208.300 ;
        RECT 107.515 207.755 107.805 208.480 ;
        RECT 109.560 208.300 109.900 209.130 ;
        RECT 111.380 208.620 111.730 209.870 ;
        RECT 115.080 208.300 115.420 209.130 ;
        RECT 116.900 208.620 117.250 209.870 ;
        RECT 120.600 208.300 120.940 209.130 ;
        RECT 122.420 208.620 122.770 209.870 ;
        RECT 126.120 208.300 126.460 209.130 ;
        RECT 127.940 208.620 128.290 209.870 ;
        RECT 130.055 209.215 132.645 210.305 ;
        RECT 130.055 208.525 131.265 209.045 ;
        RECT 131.435 208.695 132.645 209.215 ;
        RECT 133.275 209.140 133.565 210.305 ;
        RECT 133.735 209.870 139.080 210.305 ;
        RECT 139.255 209.870 144.600 210.305 ;
        RECT 107.975 207.755 113.320 208.300 ;
        RECT 113.495 207.755 118.840 208.300 ;
        RECT 119.015 207.755 124.360 208.300 ;
        RECT 124.535 207.755 129.880 208.300 ;
        RECT 130.055 207.755 132.645 208.525 ;
        RECT 133.275 207.755 133.565 208.480 ;
        RECT 135.320 208.300 135.660 209.130 ;
        RECT 137.140 208.620 137.490 209.870 ;
        RECT 140.840 208.300 141.180 209.130 ;
        RECT 142.660 208.620 143.010 209.870 ;
        RECT 145.695 209.215 146.905 210.305 ;
        RECT 145.695 208.675 146.215 209.215 ;
        RECT 146.385 208.505 146.905 209.045 ;
        RECT 133.735 207.755 139.080 208.300 ;
        RECT 139.255 207.755 144.600 208.300 ;
        RECT 145.695 207.755 146.905 208.505 ;
        RECT 17.270 207.585 146.990 207.755 ;
        RECT 17.355 206.835 18.565 207.585 ;
        RECT 18.735 207.040 24.080 207.585 ;
        RECT 24.255 207.040 29.600 207.585 ;
        RECT 29.775 207.040 35.120 207.585 ;
        RECT 35.295 207.040 40.640 207.585 ;
        RECT 17.355 206.295 17.875 206.835 ;
        RECT 18.045 206.125 18.565 206.665 ;
        RECT 20.320 206.210 20.660 207.040 ;
        RECT 17.355 205.035 18.565 206.125 ;
        RECT 22.140 205.470 22.490 206.720 ;
        RECT 25.840 206.210 26.180 207.040 ;
        RECT 27.660 205.470 28.010 206.720 ;
        RECT 31.360 206.210 31.700 207.040 ;
        RECT 33.180 205.470 33.530 206.720 ;
        RECT 36.880 206.210 37.220 207.040 ;
        RECT 40.815 206.815 42.485 207.585 ;
        RECT 43.115 206.860 43.405 207.585 ;
        RECT 43.575 207.040 48.920 207.585 ;
        RECT 38.700 205.470 39.050 206.720 ;
        RECT 40.815 206.295 41.565 206.815 ;
        RECT 41.735 206.125 42.485 206.645 ;
        RECT 45.160 206.210 45.500 207.040 ;
        RECT 49.095 206.835 50.305 207.585 ;
        RECT 18.735 205.035 24.080 205.470 ;
        RECT 24.255 205.035 29.600 205.470 ;
        RECT 29.775 205.035 35.120 205.470 ;
        RECT 35.295 205.035 40.640 205.470 ;
        RECT 40.815 205.035 42.485 206.125 ;
        RECT 43.115 205.035 43.405 206.200 ;
        RECT 46.980 205.470 47.330 206.720 ;
        RECT 49.095 206.295 49.615 206.835 ;
        RECT 50.495 206.775 50.735 207.585 ;
        RECT 50.905 206.775 51.235 207.415 ;
        RECT 51.405 206.775 51.675 207.585 ;
        RECT 51.855 206.815 54.445 207.585 ;
        RECT 49.785 206.125 50.305 206.665 ;
        RECT 50.475 206.345 50.825 206.595 ;
        RECT 50.995 206.175 51.165 206.775 ;
        RECT 51.335 206.345 51.685 206.595 ;
        RECT 51.855 206.295 53.065 206.815 ;
        RECT 55.135 206.765 55.345 207.585 ;
        RECT 55.515 206.785 55.845 207.415 ;
        RECT 43.575 205.035 48.920 205.470 ;
        RECT 49.095 205.035 50.305 206.125 ;
        RECT 50.485 206.005 51.165 206.175 ;
        RECT 50.485 205.220 50.815 206.005 ;
        RECT 51.345 205.035 51.675 206.175 ;
        RECT 53.235 206.125 54.445 206.645 ;
        RECT 55.515 206.185 55.765 206.785 ;
        RECT 56.015 206.765 56.245 207.585 ;
        RECT 56.455 207.040 61.800 207.585 ;
        RECT 55.935 206.345 56.265 206.595 ;
        RECT 58.040 206.210 58.380 207.040 ;
        RECT 61.975 206.815 63.645 207.585 ;
        RECT 63.885 207.185 64.215 207.585 ;
        RECT 64.385 207.015 64.555 207.285 ;
        RECT 64.725 207.185 65.055 207.585 ;
        RECT 65.225 207.015 65.480 207.285 ;
        RECT 51.855 205.035 54.445 206.125 ;
        RECT 55.135 205.035 55.345 206.175 ;
        RECT 55.515 205.205 55.845 206.185 ;
        RECT 56.015 205.035 56.245 206.175 ;
        RECT 59.860 205.470 60.210 206.720 ;
        RECT 61.975 206.295 62.725 206.815 ;
        RECT 62.895 206.125 63.645 206.645 ;
        RECT 56.455 205.035 61.800 205.470 ;
        RECT 61.975 205.035 63.645 206.125 ;
        RECT 63.815 206.005 64.085 207.015 ;
        RECT 64.255 206.845 65.480 207.015 ;
        RECT 66.575 206.935 66.835 207.415 ;
        RECT 67.005 207.045 67.255 207.585 ;
        RECT 64.255 206.175 64.425 206.845 ;
        RECT 64.595 206.345 64.975 206.675 ;
        RECT 65.145 206.345 65.480 206.675 ;
        RECT 64.255 206.005 64.570 206.175 ;
        RECT 63.820 205.035 64.135 205.835 ;
        RECT 64.400 205.390 64.570 206.005 ;
        RECT 64.740 205.665 64.975 206.345 ;
        RECT 65.145 205.390 65.480 206.175 ;
        RECT 64.400 205.220 65.480 205.390 ;
        RECT 66.575 205.905 66.745 206.935 ;
        RECT 67.425 206.880 67.645 207.365 ;
        RECT 66.915 206.285 67.145 206.680 ;
        RECT 67.315 206.455 67.645 206.880 ;
        RECT 67.815 207.205 68.705 207.375 ;
        RECT 67.815 206.480 67.985 207.205 ;
        RECT 68.155 206.650 68.705 207.035 ;
        RECT 68.875 206.860 69.165 207.585 ;
        RECT 69.340 206.745 69.600 207.585 ;
        RECT 69.775 206.840 70.030 207.415 ;
        RECT 70.200 207.205 70.530 207.585 ;
        RECT 70.745 207.035 70.915 207.415 ;
        RECT 71.175 207.040 76.520 207.585 ;
        RECT 76.695 207.040 82.040 207.585 ;
        RECT 70.200 206.865 70.915 207.035 ;
        RECT 67.815 206.410 68.705 206.480 ;
        RECT 67.810 206.385 68.705 206.410 ;
        RECT 67.800 206.370 68.705 206.385 ;
        RECT 67.795 206.355 68.705 206.370 ;
        RECT 67.785 206.350 68.705 206.355 ;
        RECT 67.780 206.340 68.705 206.350 ;
        RECT 67.775 206.330 68.705 206.340 ;
        RECT 67.765 206.325 68.705 206.330 ;
        RECT 67.755 206.315 68.705 206.325 ;
        RECT 67.745 206.310 68.705 206.315 ;
        RECT 67.745 206.305 68.080 206.310 ;
        RECT 67.730 206.300 68.080 206.305 ;
        RECT 67.715 206.290 68.080 206.300 ;
        RECT 67.690 206.285 68.080 206.290 ;
        RECT 66.915 206.280 68.080 206.285 ;
        RECT 66.915 206.245 68.050 206.280 ;
        RECT 66.915 206.220 68.015 206.245 ;
        RECT 66.915 206.190 67.985 206.220 ;
        RECT 66.915 206.160 67.965 206.190 ;
        RECT 66.915 206.130 67.945 206.160 ;
        RECT 66.915 206.120 67.875 206.130 ;
        RECT 66.915 206.110 67.850 206.120 ;
        RECT 66.915 206.095 67.830 206.110 ;
        RECT 66.915 206.080 67.810 206.095 ;
        RECT 67.020 206.070 67.805 206.080 ;
        RECT 67.020 206.035 67.790 206.070 ;
        RECT 66.575 205.205 66.850 205.905 ;
        RECT 67.020 205.785 67.775 206.035 ;
        RECT 67.945 205.715 68.275 205.960 ;
        RECT 68.445 205.860 68.705 206.310 ;
        RECT 68.090 205.690 68.275 205.715 ;
        RECT 68.090 205.590 68.705 205.690 ;
        RECT 67.020 205.035 67.275 205.580 ;
        RECT 67.445 205.205 67.925 205.545 ;
        RECT 68.100 205.035 68.705 205.590 ;
        RECT 68.875 205.035 69.165 206.200 ;
        RECT 69.340 205.035 69.600 206.185 ;
        RECT 69.775 206.110 69.945 206.840 ;
        RECT 70.200 206.675 70.370 206.865 ;
        RECT 70.115 206.345 70.370 206.675 ;
        RECT 70.200 206.135 70.370 206.345 ;
        RECT 70.650 206.315 71.005 206.685 ;
        RECT 72.760 206.210 73.100 207.040 ;
        RECT 69.775 205.205 70.030 206.110 ;
        RECT 70.200 205.965 70.915 206.135 ;
        RECT 70.200 205.035 70.530 205.795 ;
        RECT 70.745 205.205 70.915 205.965 ;
        RECT 74.580 205.470 74.930 206.720 ;
        RECT 78.280 206.210 78.620 207.040 ;
        RECT 82.215 206.815 84.805 207.585 ;
        RECT 80.100 205.470 80.450 206.720 ;
        RECT 82.215 206.295 83.425 206.815 ;
        RECT 83.595 206.125 84.805 206.645 ;
        RECT 71.175 205.035 76.520 205.470 ;
        RECT 76.695 205.035 82.040 205.470 ;
        RECT 82.215 205.035 84.805 206.125 ;
        RECT 85.435 206.640 85.775 207.415 ;
        RECT 85.945 207.125 86.115 207.585 ;
        RECT 86.355 207.150 86.715 207.415 ;
        RECT 86.355 207.145 86.710 207.150 ;
        RECT 86.355 207.135 86.705 207.145 ;
        RECT 86.355 207.130 86.700 207.135 ;
        RECT 86.355 207.120 86.695 207.130 ;
        RECT 87.345 207.125 87.515 207.585 ;
        RECT 86.355 207.115 86.690 207.120 ;
        RECT 86.355 207.105 86.680 207.115 ;
        RECT 86.355 207.095 86.670 207.105 ;
        RECT 86.355 206.955 86.655 207.095 ;
        RECT 85.945 206.765 86.655 206.955 ;
        RECT 86.845 206.955 87.175 207.035 ;
        RECT 87.685 206.955 88.025 207.415 ;
        RECT 88.195 207.040 93.540 207.585 ;
        RECT 86.845 206.765 88.025 206.955 ;
        RECT 85.435 205.205 85.715 206.640 ;
        RECT 85.945 206.195 86.230 206.765 ;
        RECT 86.415 206.365 86.885 206.595 ;
        RECT 87.055 206.575 87.385 206.595 ;
        RECT 87.055 206.395 87.505 206.575 ;
        RECT 87.695 206.395 88.025 206.595 ;
        RECT 85.945 205.980 87.095 206.195 ;
        RECT 85.885 205.035 86.595 205.810 ;
        RECT 86.765 205.205 87.095 205.980 ;
        RECT 87.290 205.280 87.505 206.395 ;
        RECT 87.795 206.055 88.025 206.395 ;
        RECT 89.780 206.210 90.120 207.040 ;
        RECT 94.635 206.860 94.925 207.585 ;
        RECT 95.115 206.775 95.355 207.585 ;
        RECT 95.525 206.775 95.855 207.415 ;
        RECT 96.025 206.775 96.295 207.585 ;
        RECT 96.475 207.040 101.820 207.585 ;
        RECT 101.995 207.040 107.340 207.585 ;
        RECT 87.685 205.035 88.015 205.755 ;
        RECT 91.600 205.470 91.950 206.720 ;
        RECT 95.095 206.345 95.445 206.595 ;
        RECT 88.195 205.035 93.540 205.470 ;
        RECT 94.635 205.035 94.925 206.200 ;
        RECT 95.615 206.175 95.785 206.775 ;
        RECT 95.955 206.345 96.305 206.595 ;
        RECT 98.060 206.210 98.400 207.040 ;
        RECT 95.105 206.005 95.785 206.175 ;
        RECT 95.105 205.220 95.435 206.005 ;
        RECT 95.965 205.035 96.295 206.175 ;
        RECT 99.880 205.470 100.230 206.720 ;
        RECT 103.580 206.210 103.920 207.040 ;
        RECT 107.515 206.815 110.105 207.585 ;
        RECT 110.850 206.955 111.135 207.415 ;
        RECT 111.305 207.125 111.575 207.585 ;
        RECT 105.400 205.470 105.750 206.720 ;
        RECT 107.515 206.295 108.725 206.815 ;
        RECT 110.850 206.785 111.805 206.955 ;
        RECT 108.895 206.125 110.105 206.645 ;
        RECT 96.475 205.035 101.820 205.470 ;
        RECT 101.995 205.035 107.340 205.470 ;
        RECT 107.515 205.035 110.105 206.125 ;
        RECT 110.735 206.055 111.425 206.615 ;
        RECT 111.595 205.885 111.805 206.785 ;
        RECT 110.850 205.665 111.805 205.885 ;
        RECT 111.975 206.615 112.375 207.415 ;
        RECT 112.565 206.955 112.845 207.415 ;
        RECT 113.365 207.125 113.690 207.585 ;
        RECT 112.565 206.785 113.690 206.955 ;
        RECT 113.860 206.845 114.245 207.415 ;
        RECT 114.415 207.040 119.760 207.585 ;
        RECT 113.240 206.675 113.690 206.785 ;
        RECT 111.975 206.055 113.070 206.615 ;
        RECT 113.240 206.345 113.795 206.675 ;
        RECT 110.850 205.205 111.135 205.665 ;
        RECT 111.305 205.035 111.575 205.495 ;
        RECT 111.975 205.205 112.375 206.055 ;
        RECT 113.240 205.885 113.690 206.345 ;
        RECT 113.965 206.175 114.245 206.845 ;
        RECT 116.000 206.210 116.340 207.040 ;
        RECT 120.395 206.860 120.685 207.585 ;
        RECT 120.855 207.040 126.200 207.585 ;
        RECT 126.375 207.040 131.720 207.585 ;
        RECT 131.895 207.040 137.240 207.585 ;
        RECT 137.415 207.040 142.760 207.585 ;
        RECT 112.565 205.665 113.690 205.885 ;
        RECT 112.565 205.205 112.845 205.665 ;
        RECT 113.365 205.035 113.690 205.495 ;
        RECT 113.860 205.205 114.245 206.175 ;
        RECT 117.820 205.470 118.170 206.720 ;
        RECT 122.440 206.210 122.780 207.040 ;
        RECT 114.415 205.035 119.760 205.470 ;
        RECT 120.395 205.035 120.685 206.200 ;
        RECT 124.260 205.470 124.610 206.720 ;
        RECT 127.960 206.210 128.300 207.040 ;
        RECT 129.780 205.470 130.130 206.720 ;
        RECT 133.480 206.210 133.820 207.040 ;
        RECT 135.300 205.470 135.650 206.720 ;
        RECT 139.000 206.210 139.340 207.040 ;
        RECT 142.935 206.815 145.525 207.585 ;
        RECT 145.695 206.835 146.905 207.585 ;
        RECT 140.820 205.470 141.170 206.720 ;
        RECT 142.935 206.295 144.145 206.815 ;
        RECT 144.315 206.125 145.525 206.645 ;
        RECT 120.855 205.035 126.200 205.470 ;
        RECT 126.375 205.035 131.720 205.470 ;
        RECT 131.895 205.035 137.240 205.470 ;
        RECT 137.415 205.035 142.760 205.470 ;
        RECT 142.935 205.035 145.525 206.125 ;
        RECT 145.695 206.125 146.215 206.665 ;
        RECT 146.385 206.295 146.905 206.835 ;
        RECT 145.695 205.035 146.905 206.125 ;
        RECT 17.270 204.865 146.990 205.035 ;
        RECT 17.355 203.775 18.565 204.865 ;
        RECT 18.735 204.430 24.080 204.865 ;
        RECT 17.355 203.065 17.875 203.605 ;
        RECT 18.045 203.235 18.565 203.775 ;
        RECT 17.355 202.315 18.565 203.065 ;
        RECT 20.320 202.860 20.660 203.690 ;
        RECT 22.140 203.180 22.490 204.430 ;
        RECT 24.255 203.775 25.925 204.865 ;
        RECT 24.255 203.085 25.005 203.605 ;
        RECT 25.175 203.255 25.925 203.775 ;
        RECT 26.105 203.895 26.435 204.695 ;
        RECT 26.605 204.065 26.835 204.865 ;
        RECT 27.005 203.895 27.335 204.695 ;
        RECT 26.105 203.725 27.335 203.895 ;
        RECT 27.505 203.725 27.760 204.865 ;
        RECT 27.935 203.775 29.605 204.865 ;
        RECT 26.095 203.225 26.405 203.555 ;
        RECT 18.735 202.315 24.080 202.860 ;
        RECT 24.255 202.315 25.925 203.085 ;
        RECT 26.105 202.825 26.435 203.055 ;
        RECT 26.610 202.995 26.985 203.555 ;
        RECT 27.155 202.825 27.335 203.725 ;
        RECT 27.520 202.975 27.740 203.555 ;
        RECT 27.935 203.085 28.685 203.605 ;
        RECT 28.855 203.255 29.605 203.775 ;
        RECT 30.235 203.700 30.525 204.865 ;
        RECT 30.695 204.430 36.040 204.865 ;
        RECT 26.105 202.485 27.335 202.825 ;
        RECT 27.505 202.315 27.760 202.805 ;
        RECT 27.935 202.315 29.605 203.085 ;
        RECT 30.235 202.315 30.525 203.040 ;
        RECT 32.280 202.860 32.620 203.690 ;
        RECT 34.100 203.180 34.450 204.430 ;
        RECT 36.215 203.775 38.805 204.865 ;
        RECT 36.215 203.085 37.425 203.605 ;
        RECT 37.595 203.255 38.805 203.775 ;
        RECT 38.975 203.895 39.245 204.665 ;
        RECT 39.415 204.085 39.745 204.865 ;
        RECT 39.950 204.260 40.135 204.665 ;
        RECT 40.305 204.440 40.640 204.865 ;
        RECT 40.815 204.430 46.160 204.865 ;
        RECT 46.335 204.430 51.680 204.865 ;
        RECT 39.950 204.085 40.615 204.260 ;
        RECT 38.975 203.725 40.105 203.895 ;
        RECT 30.695 202.315 36.040 202.860 ;
        RECT 36.215 202.315 38.805 203.085 ;
        RECT 38.975 202.815 39.145 203.725 ;
        RECT 39.315 202.975 39.675 203.555 ;
        RECT 39.855 203.225 40.105 203.725 ;
        RECT 40.275 203.055 40.615 204.085 ;
        RECT 39.930 202.885 40.615 203.055 ;
        RECT 38.975 202.485 39.235 202.815 ;
        RECT 39.445 202.315 39.720 202.795 ;
        RECT 39.930 202.485 40.135 202.885 ;
        RECT 42.400 202.860 42.740 203.690 ;
        RECT 44.220 203.180 44.570 204.430 ;
        RECT 47.920 202.860 48.260 203.690 ;
        RECT 49.740 203.180 50.090 204.430 ;
        RECT 51.855 203.775 53.525 204.865 ;
        RECT 51.855 203.085 52.605 203.605 ;
        RECT 52.775 203.255 53.525 203.775 ;
        RECT 53.880 203.895 54.270 204.070 ;
        RECT 54.755 204.065 55.085 204.865 ;
        RECT 55.255 204.075 55.790 204.695 ;
        RECT 53.880 203.725 55.305 203.895 ;
        RECT 40.305 202.315 40.640 202.715 ;
        RECT 40.815 202.315 46.160 202.860 ;
        RECT 46.335 202.315 51.680 202.860 ;
        RECT 51.855 202.315 53.525 203.085 ;
        RECT 53.755 202.995 54.110 203.555 ;
        RECT 54.280 202.825 54.450 203.725 ;
        RECT 54.620 202.995 54.885 203.555 ;
        RECT 55.135 203.225 55.305 203.725 ;
        RECT 55.475 203.055 55.790 204.075 ;
        RECT 55.995 203.700 56.285 204.865 ;
        RECT 56.465 204.145 56.795 204.865 ;
        RECT 56.455 203.505 56.685 203.845 ;
        RECT 56.975 203.505 57.190 204.620 ;
        RECT 57.385 203.920 57.715 204.695 ;
        RECT 57.885 204.090 58.595 204.865 ;
        RECT 57.385 203.705 58.535 203.920 ;
        RECT 56.455 203.305 56.785 203.505 ;
        RECT 56.975 203.325 57.425 203.505 ;
        RECT 57.095 203.305 57.425 203.325 ;
        RECT 57.595 203.305 58.065 203.535 ;
        RECT 58.250 203.135 58.535 203.705 ;
        RECT 58.765 203.260 59.045 204.695 ;
        RECT 59.225 203.915 59.500 204.685 ;
        RECT 59.670 204.255 60.000 204.685 ;
        RECT 60.170 204.425 60.365 204.865 ;
        RECT 60.545 204.255 60.875 204.685 ;
        RECT 61.055 204.430 66.400 204.865 ;
        RECT 66.575 204.430 71.920 204.865 ;
        RECT 72.095 204.430 77.440 204.865 ;
        RECT 59.670 204.085 60.875 204.255 ;
        RECT 59.225 203.725 59.810 203.915 ;
        RECT 59.980 203.755 60.875 204.085 ;
        RECT 53.860 202.315 54.100 202.825 ;
        RECT 54.280 202.495 54.560 202.825 ;
        RECT 54.790 202.315 55.005 202.825 ;
        RECT 55.175 202.485 55.790 203.055 ;
        RECT 55.995 202.315 56.285 203.040 ;
        RECT 56.455 202.945 57.635 203.135 ;
        RECT 56.455 202.485 56.795 202.945 ;
        RECT 57.305 202.865 57.635 202.945 ;
        RECT 57.825 202.945 58.535 203.135 ;
        RECT 57.825 202.805 58.125 202.945 ;
        RECT 57.810 202.795 58.125 202.805 ;
        RECT 57.800 202.785 58.125 202.795 ;
        RECT 57.790 202.780 58.125 202.785 ;
        RECT 56.965 202.315 57.135 202.775 ;
        RECT 57.785 202.770 58.125 202.780 ;
        RECT 57.780 202.765 58.125 202.770 ;
        RECT 57.775 202.755 58.125 202.765 ;
        RECT 57.770 202.750 58.125 202.755 ;
        RECT 57.765 202.485 58.125 202.750 ;
        RECT 58.365 202.315 58.535 202.775 ;
        RECT 58.705 202.485 59.045 203.260 ;
        RECT 59.225 202.905 59.465 203.555 ;
        RECT 59.635 203.055 59.810 203.725 ;
        RECT 59.980 203.225 60.395 203.555 ;
        RECT 60.575 203.225 60.870 203.555 ;
        RECT 59.635 202.875 59.965 203.055 ;
        RECT 59.240 202.315 59.570 202.705 ;
        RECT 59.740 202.495 59.965 202.875 ;
        RECT 60.165 202.605 60.395 203.225 ;
        RECT 60.575 202.315 60.875 203.045 ;
        RECT 62.640 202.860 62.980 203.690 ;
        RECT 64.460 203.180 64.810 204.430 ;
        RECT 68.160 202.860 68.500 203.690 ;
        RECT 69.980 203.180 70.330 204.430 ;
        RECT 73.680 202.860 74.020 203.690 ;
        RECT 75.500 203.180 75.850 204.430 ;
        RECT 77.615 203.775 79.285 204.865 ;
        RECT 77.615 203.085 78.365 203.605 ;
        RECT 78.535 203.255 79.285 203.775 ;
        RECT 79.920 203.725 80.240 204.865 ;
        RECT 80.420 203.555 80.615 204.605 ;
        RECT 80.795 204.015 81.125 204.695 ;
        RECT 81.325 204.065 81.580 204.865 ;
        RECT 80.795 203.735 81.145 204.015 ;
        RECT 79.980 203.505 80.240 203.555 ;
        RECT 79.975 203.335 80.240 203.505 ;
        RECT 79.980 203.225 80.240 203.335 ;
        RECT 80.420 203.225 80.805 203.555 ;
        RECT 80.975 203.355 81.145 203.735 ;
        RECT 81.335 203.525 81.580 203.885 ;
        RECT 81.755 203.700 82.045 204.865 ;
        RECT 82.305 204.195 82.475 204.695 ;
        RECT 82.645 204.365 82.975 204.865 ;
        RECT 82.305 204.025 82.970 204.195 ;
        RECT 80.975 203.185 81.495 203.355 ;
        RECT 82.220 203.205 82.570 203.855 ;
        RECT 61.055 202.315 66.400 202.860 ;
        RECT 66.575 202.315 71.920 202.860 ;
        RECT 72.095 202.315 77.440 202.860 ;
        RECT 77.615 202.315 79.285 203.085 ;
        RECT 79.920 202.845 81.135 203.015 ;
        RECT 79.920 202.495 80.210 202.845 ;
        RECT 80.405 202.315 80.735 202.675 ;
        RECT 80.905 202.540 81.135 202.845 ;
        RECT 81.325 202.825 81.495 203.185 ;
        RECT 81.325 202.655 81.525 202.825 ;
        RECT 81.325 202.620 81.495 202.655 ;
        RECT 81.755 202.315 82.045 203.040 ;
        RECT 82.740 203.035 82.970 204.025 ;
        RECT 82.305 202.865 82.970 203.035 ;
        RECT 82.305 202.575 82.475 202.865 ;
        RECT 82.645 202.315 82.975 202.695 ;
        RECT 83.145 202.575 83.330 204.695 ;
        RECT 83.570 204.405 83.835 204.865 ;
        RECT 84.005 204.270 84.255 204.695 ;
        RECT 84.465 204.420 85.570 204.590 ;
        RECT 83.950 204.140 84.255 204.270 ;
        RECT 83.500 202.945 83.780 203.895 ;
        RECT 83.950 203.035 84.120 204.140 ;
        RECT 84.290 203.355 84.530 203.950 ;
        RECT 84.700 203.885 85.230 204.250 ;
        RECT 84.700 203.185 84.870 203.885 ;
        RECT 85.400 203.805 85.570 204.420 ;
        RECT 85.740 204.065 85.910 204.865 ;
        RECT 86.080 204.365 86.330 204.695 ;
        RECT 86.555 204.395 87.440 204.565 ;
        RECT 85.400 203.715 85.910 203.805 ;
        RECT 83.950 202.905 84.175 203.035 ;
        RECT 84.345 202.965 84.870 203.185 ;
        RECT 85.040 203.545 85.910 203.715 ;
        RECT 83.585 202.315 83.835 202.775 ;
        RECT 84.005 202.765 84.175 202.905 ;
        RECT 85.040 202.765 85.210 203.545 ;
        RECT 85.740 203.475 85.910 203.545 ;
        RECT 85.420 203.295 85.620 203.325 ;
        RECT 86.080 203.295 86.250 204.365 ;
        RECT 86.420 203.475 86.610 204.195 ;
        RECT 85.420 202.995 86.250 203.295 ;
        RECT 86.780 203.265 87.100 204.225 ;
        RECT 84.005 202.595 84.340 202.765 ;
        RECT 84.535 202.595 85.210 202.765 ;
        RECT 85.530 202.315 85.900 202.815 ;
        RECT 86.080 202.765 86.250 202.995 ;
        RECT 86.635 202.935 87.100 203.265 ;
        RECT 87.270 203.555 87.440 204.395 ;
        RECT 87.620 204.365 87.935 204.865 ;
        RECT 88.165 204.135 88.505 204.695 ;
        RECT 87.610 203.760 88.505 204.135 ;
        RECT 88.675 203.855 88.845 204.865 ;
        RECT 88.315 203.555 88.505 203.760 ;
        RECT 89.015 203.805 89.345 204.650 ;
        RECT 89.015 203.725 89.405 203.805 ;
        RECT 89.190 203.675 89.405 203.725 ;
        RECT 87.270 203.225 88.145 203.555 ;
        RECT 88.315 203.225 89.065 203.555 ;
        RECT 87.270 202.765 87.440 203.225 ;
        RECT 88.315 203.055 88.515 203.225 ;
        RECT 89.235 203.095 89.405 203.675 ;
        RECT 89.180 203.055 89.405 203.095 ;
        RECT 86.080 202.595 86.485 202.765 ;
        RECT 86.655 202.595 87.440 202.765 ;
        RECT 87.715 202.315 87.925 202.845 ;
        RECT 88.185 202.530 88.515 203.055 ;
        RECT 89.025 202.970 89.405 203.055 ;
        RECT 89.575 203.725 89.960 204.695 ;
        RECT 90.130 204.405 90.455 204.865 ;
        RECT 90.975 204.235 91.255 204.695 ;
        RECT 90.130 204.015 91.255 204.235 ;
        RECT 89.575 203.055 89.855 203.725 ;
        RECT 90.130 203.555 90.580 204.015 ;
        RECT 91.445 203.845 91.845 204.695 ;
        RECT 92.245 204.405 92.515 204.865 ;
        RECT 92.685 204.235 92.970 204.695 ;
        RECT 90.025 203.225 90.580 203.555 ;
        RECT 90.750 203.285 91.845 203.845 ;
        RECT 90.130 203.115 90.580 203.225 ;
        RECT 88.685 202.315 88.855 202.925 ;
        RECT 89.025 202.535 89.355 202.970 ;
        RECT 89.575 202.485 89.960 203.055 ;
        RECT 90.130 202.945 91.255 203.115 ;
        RECT 90.130 202.315 90.455 202.775 ;
        RECT 90.975 202.485 91.255 202.945 ;
        RECT 91.445 202.485 91.845 203.285 ;
        RECT 92.015 204.015 92.970 204.235 ;
        RECT 92.015 203.115 92.225 204.015 ;
        RECT 92.395 203.285 93.085 203.845 ;
        RECT 93.255 203.725 93.530 204.695 ;
        RECT 93.740 204.065 94.020 204.865 ;
        RECT 94.190 204.355 95.805 204.685 ;
        RECT 94.190 204.015 95.365 204.185 ;
        RECT 94.190 203.895 94.360 204.015 ;
        RECT 93.700 203.725 94.360 203.895 ;
        RECT 92.015 202.945 92.970 203.115 ;
        RECT 92.245 202.315 92.515 202.775 ;
        RECT 92.685 202.485 92.970 202.945 ;
        RECT 93.255 202.990 93.425 203.725 ;
        RECT 93.700 203.555 93.870 203.725 ;
        RECT 94.620 203.555 94.865 203.845 ;
        RECT 95.035 203.725 95.365 204.015 ;
        RECT 95.625 203.555 95.795 204.115 ;
        RECT 96.045 203.725 96.305 204.865 ;
        RECT 96.565 204.195 96.735 204.695 ;
        RECT 96.905 204.365 97.235 204.865 ;
        RECT 96.565 204.025 97.230 204.195 ;
        RECT 93.595 203.225 93.870 203.555 ;
        RECT 94.040 203.225 94.865 203.555 ;
        RECT 95.080 203.225 95.795 203.555 ;
        RECT 95.965 203.305 96.300 203.555 ;
        RECT 93.700 203.055 93.870 203.225 ;
        RECT 95.545 203.135 95.795 203.225 ;
        RECT 96.480 203.205 96.830 203.855 ;
        RECT 93.255 202.645 93.530 202.990 ;
        RECT 93.700 202.885 95.365 203.055 ;
        RECT 93.720 202.315 94.095 202.715 ;
        RECT 94.265 202.535 94.435 202.885 ;
        RECT 94.605 202.315 94.935 202.715 ;
        RECT 95.105 202.485 95.365 202.885 ;
        RECT 95.545 202.715 95.875 203.135 ;
        RECT 96.045 202.315 96.305 203.135 ;
        RECT 97.000 203.035 97.230 204.025 ;
        RECT 96.565 202.865 97.230 203.035 ;
        RECT 96.565 202.575 96.735 202.865 ;
        RECT 96.905 202.315 97.235 202.695 ;
        RECT 97.405 202.575 97.590 204.695 ;
        RECT 97.830 204.405 98.095 204.865 ;
        RECT 98.265 204.270 98.515 204.695 ;
        RECT 98.725 204.420 99.830 204.590 ;
        RECT 98.210 204.140 98.515 204.270 ;
        RECT 97.760 202.945 98.040 203.895 ;
        RECT 98.210 203.035 98.380 204.140 ;
        RECT 98.550 203.355 98.790 203.950 ;
        RECT 98.960 203.885 99.490 204.250 ;
        RECT 98.960 203.185 99.130 203.885 ;
        RECT 99.660 203.805 99.830 204.420 ;
        RECT 100.000 204.065 100.170 204.865 ;
        RECT 100.340 204.365 100.590 204.695 ;
        RECT 100.815 204.395 101.700 204.565 ;
        RECT 99.660 203.715 100.170 203.805 ;
        RECT 98.210 202.905 98.435 203.035 ;
        RECT 98.605 202.965 99.130 203.185 ;
        RECT 99.300 203.545 100.170 203.715 ;
        RECT 97.845 202.315 98.095 202.775 ;
        RECT 98.265 202.765 98.435 202.905 ;
        RECT 99.300 202.765 99.470 203.545 ;
        RECT 100.000 203.475 100.170 203.545 ;
        RECT 99.680 203.295 99.880 203.325 ;
        RECT 100.340 203.295 100.510 204.365 ;
        RECT 100.680 203.475 100.870 204.195 ;
        RECT 99.680 202.995 100.510 203.295 ;
        RECT 101.040 203.265 101.360 204.225 ;
        RECT 98.265 202.595 98.600 202.765 ;
        RECT 98.795 202.595 99.470 202.765 ;
        RECT 99.790 202.315 100.160 202.815 ;
        RECT 100.340 202.765 100.510 202.995 ;
        RECT 100.895 202.935 101.360 203.265 ;
        RECT 101.530 203.555 101.700 204.395 ;
        RECT 101.880 204.365 102.195 204.865 ;
        RECT 102.425 204.135 102.765 204.695 ;
        RECT 101.870 203.760 102.765 204.135 ;
        RECT 102.935 203.855 103.105 204.865 ;
        RECT 102.575 203.555 102.765 203.760 ;
        RECT 103.275 203.805 103.605 204.650 ;
        RECT 103.275 203.725 103.665 203.805 ;
        RECT 103.450 203.675 103.665 203.725 ;
        RECT 101.530 203.225 102.405 203.555 ;
        RECT 102.575 203.225 103.325 203.555 ;
        RECT 101.530 202.765 101.700 203.225 ;
        RECT 102.575 203.055 102.775 203.225 ;
        RECT 103.495 203.095 103.665 203.675 ;
        RECT 103.440 203.055 103.665 203.095 ;
        RECT 100.340 202.595 100.745 202.765 ;
        RECT 100.915 202.595 101.700 202.765 ;
        RECT 101.975 202.315 102.185 202.845 ;
        RECT 102.445 202.530 102.775 203.055 ;
        RECT 103.285 202.970 103.665 203.055 ;
        RECT 103.835 203.725 104.220 204.695 ;
        RECT 104.390 204.405 104.715 204.865 ;
        RECT 105.235 204.235 105.515 204.695 ;
        RECT 104.390 204.015 105.515 204.235 ;
        RECT 103.835 203.055 104.115 203.725 ;
        RECT 104.390 203.555 104.840 204.015 ;
        RECT 105.705 203.845 106.105 204.695 ;
        RECT 106.505 204.405 106.775 204.865 ;
        RECT 106.945 204.235 107.230 204.695 ;
        RECT 104.285 203.225 104.840 203.555 ;
        RECT 105.010 203.285 106.105 203.845 ;
        RECT 104.390 203.115 104.840 203.225 ;
        RECT 102.945 202.315 103.115 202.925 ;
        RECT 103.285 202.535 103.615 202.970 ;
        RECT 103.835 202.485 104.220 203.055 ;
        RECT 104.390 202.945 105.515 203.115 ;
        RECT 104.390 202.315 104.715 202.775 ;
        RECT 105.235 202.485 105.515 202.945 ;
        RECT 105.705 202.485 106.105 203.285 ;
        RECT 106.275 204.015 107.230 204.235 ;
        RECT 106.275 203.115 106.485 204.015 ;
        RECT 106.655 203.285 107.345 203.845 ;
        RECT 107.515 203.700 107.805 204.865 ;
        RECT 108.495 203.805 108.825 204.650 ;
        RECT 108.995 203.855 109.165 204.865 ;
        RECT 109.335 204.135 109.675 204.695 ;
        RECT 109.905 204.365 110.220 204.865 ;
        RECT 110.400 204.395 111.285 204.565 ;
        RECT 108.435 203.725 108.825 203.805 ;
        RECT 109.335 203.760 110.230 204.135 ;
        RECT 108.435 203.675 108.650 203.725 ;
        RECT 106.275 202.945 107.230 203.115 ;
        RECT 108.435 203.095 108.605 203.675 ;
        RECT 109.335 203.555 109.525 203.760 ;
        RECT 110.400 203.555 110.570 204.395 ;
        RECT 111.510 204.365 111.760 204.695 ;
        RECT 108.775 203.225 109.525 203.555 ;
        RECT 109.695 203.225 110.570 203.555 ;
        RECT 108.435 203.055 108.660 203.095 ;
        RECT 109.325 203.055 109.525 203.225 ;
        RECT 106.505 202.315 106.775 202.775 ;
        RECT 106.945 202.485 107.230 202.945 ;
        RECT 107.515 202.315 107.805 203.040 ;
        RECT 108.435 202.970 108.815 203.055 ;
        RECT 108.485 202.535 108.815 202.970 ;
        RECT 108.985 202.315 109.155 202.925 ;
        RECT 109.325 202.530 109.655 203.055 ;
        RECT 109.915 202.315 110.125 202.845 ;
        RECT 110.400 202.765 110.570 203.225 ;
        RECT 110.740 203.265 111.060 204.225 ;
        RECT 111.230 203.475 111.420 204.195 ;
        RECT 111.590 203.295 111.760 204.365 ;
        RECT 111.930 204.065 112.100 204.865 ;
        RECT 112.270 204.420 113.375 204.590 ;
        RECT 112.270 203.805 112.440 204.420 ;
        RECT 113.585 204.270 113.835 204.695 ;
        RECT 114.005 204.405 114.270 204.865 ;
        RECT 112.610 203.885 113.140 204.250 ;
        RECT 113.585 204.140 113.890 204.270 ;
        RECT 111.930 203.715 112.440 203.805 ;
        RECT 111.930 203.545 112.800 203.715 ;
        RECT 111.930 203.475 112.100 203.545 ;
        RECT 112.220 203.295 112.420 203.325 ;
        RECT 110.740 202.935 111.205 203.265 ;
        RECT 111.590 202.995 112.420 203.295 ;
        RECT 111.590 202.765 111.760 202.995 ;
        RECT 110.400 202.595 111.185 202.765 ;
        RECT 111.355 202.595 111.760 202.765 ;
        RECT 111.940 202.315 112.310 202.815 ;
        RECT 112.630 202.765 112.800 203.545 ;
        RECT 112.970 203.185 113.140 203.885 ;
        RECT 113.310 203.355 113.550 203.950 ;
        RECT 112.970 202.965 113.495 203.185 ;
        RECT 113.720 203.035 113.890 204.140 ;
        RECT 113.665 202.905 113.890 203.035 ;
        RECT 114.060 202.945 114.340 203.895 ;
        RECT 113.665 202.765 113.835 202.905 ;
        RECT 112.630 202.595 113.305 202.765 ;
        RECT 113.500 202.595 113.835 202.765 ;
        RECT 114.005 202.315 114.255 202.775 ;
        RECT 114.510 202.575 114.695 204.695 ;
        RECT 114.865 204.365 115.195 204.865 ;
        RECT 115.365 204.195 115.535 204.695 ;
        RECT 115.795 204.430 121.140 204.865 ;
        RECT 121.315 204.430 126.660 204.865 ;
        RECT 126.835 204.430 132.180 204.865 ;
        RECT 114.870 204.025 115.535 204.195 ;
        RECT 114.870 203.035 115.100 204.025 ;
        RECT 115.270 203.205 115.620 203.855 ;
        RECT 114.870 202.865 115.535 203.035 ;
        RECT 114.865 202.315 115.195 202.695 ;
        RECT 115.365 202.575 115.535 202.865 ;
        RECT 117.380 202.860 117.720 203.690 ;
        RECT 119.200 203.180 119.550 204.430 ;
        RECT 122.900 202.860 123.240 203.690 ;
        RECT 124.720 203.180 125.070 204.430 ;
        RECT 128.420 202.860 128.760 203.690 ;
        RECT 130.240 203.180 130.590 204.430 ;
        RECT 133.275 203.700 133.565 204.865 ;
        RECT 133.735 204.430 139.080 204.865 ;
        RECT 139.255 204.430 144.600 204.865 ;
        RECT 115.795 202.315 121.140 202.860 ;
        RECT 121.315 202.315 126.660 202.860 ;
        RECT 126.835 202.315 132.180 202.860 ;
        RECT 133.275 202.315 133.565 203.040 ;
        RECT 135.320 202.860 135.660 203.690 ;
        RECT 137.140 203.180 137.490 204.430 ;
        RECT 140.840 202.860 141.180 203.690 ;
        RECT 142.660 203.180 143.010 204.430 ;
        RECT 145.695 203.775 146.905 204.865 ;
        RECT 145.695 203.235 146.215 203.775 ;
        RECT 146.385 203.065 146.905 203.605 ;
        RECT 133.735 202.315 139.080 202.860 ;
        RECT 139.255 202.315 144.600 202.860 ;
        RECT 145.695 202.315 146.905 203.065 ;
        RECT 17.270 202.145 146.990 202.315 ;
        RECT 17.355 201.395 18.565 202.145 ;
        RECT 18.825 201.595 18.995 201.975 ;
        RECT 19.175 201.765 19.505 202.145 ;
        RECT 18.825 201.425 19.490 201.595 ;
        RECT 19.685 201.470 19.945 201.975 ;
        RECT 17.355 200.855 17.875 201.395 ;
        RECT 18.045 200.685 18.565 201.225 ;
        RECT 18.755 200.875 19.085 201.245 ;
        RECT 19.320 201.170 19.490 201.425 ;
        RECT 19.320 200.840 19.605 201.170 ;
        RECT 19.320 200.695 19.490 200.840 ;
        RECT 17.355 199.595 18.565 200.685 ;
        RECT 18.825 200.525 19.490 200.695 ;
        RECT 19.775 200.670 19.945 201.470 ;
        RECT 20.115 201.395 21.325 202.145 ;
        RECT 21.500 201.640 21.835 202.145 ;
        RECT 22.005 201.575 22.245 201.950 ;
        RECT 22.525 201.815 22.695 201.960 ;
        RECT 22.525 201.620 22.900 201.815 ;
        RECT 23.260 201.650 23.655 202.145 ;
        RECT 20.115 200.855 20.635 201.395 ;
        RECT 20.805 200.685 21.325 201.225 ;
        RECT 18.825 199.765 18.995 200.525 ;
        RECT 19.175 199.595 19.505 200.355 ;
        RECT 19.675 199.765 19.945 200.670 ;
        RECT 20.115 199.595 21.325 200.685 ;
        RECT 21.555 200.615 21.855 201.465 ;
        RECT 22.025 201.425 22.245 201.575 ;
        RECT 22.025 201.095 22.560 201.425 ;
        RECT 22.730 201.285 22.900 201.620 ;
        RECT 23.825 201.455 24.065 201.975 ;
        RECT 22.025 200.445 22.260 201.095 ;
        RECT 22.730 200.925 23.715 201.285 ;
        RECT 21.585 200.215 22.260 200.445 ;
        RECT 22.430 200.905 23.715 200.925 ;
        RECT 22.430 200.755 23.290 200.905 ;
        RECT 21.585 199.785 21.755 200.215 ;
        RECT 21.925 199.595 22.255 200.045 ;
        RECT 22.430 199.810 22.715 200.755 ;
        RECT 23.890 200.650 24.065 201.455 ;
        RECT 25.265 201.595 25.435 201.885 ;
        RECT 25.605 201.765 25.935 202.145 ;
        RECT 25.265 201.425 25.930 201.595 ;
        RECT 22.890 200.275 23.585 200.585 ;
        RECT 22.895 199.595 23.580 200.065 ;
        RECT 23.760 199.865 24.065 200.650 ;
        RECT 25.180 200.605 25.530 201.255 ;
        RECT 25.700 200.435 25.930 201.425 ;
        RECT 25.265 200.265 25.930 200.435 ;
        RECT 25.265 199.765 25.435 200.265 ;
        RECT 25.605 199.595 25.935 200.095 ;
        RECT 26.105 199.765 26.290 201.885 ;
        RECT 26.545 201.685 26.795 202.145 ;
        RECT 26.965 201.695 27.300 201.865 ;
        RECT 27.495 201.695 28.170 201.865 ;
        RECT 26.965 201.555 27.135 201.695 ;
        RECT 26.460 200.565 26.740 201.515 ;
        RECT 26.910 201.425 27.135 201.555 ;
        RECT 26.910 200.320 27.080 201.425 ;
        RECT 27.305 201.275 27.830 201.495 ;
        RECT 27.250 200.510 27.490 201.105 ;
        RECT 27.660 200.575 27.830 201.275 ;
        RECT 28.000 200.915 28.170 201.695 ;
        RECT 28.490 201.645 28.860 202.145 ;
        RECT 29.040 201.695 29.445 201.865 ;
        RECT 29.615 201.695 30.400 201.865 ;
        RECT 29.040 201.465 29.210 201.695 ;
        RECT 28.380 201.165 29.210 201.465 ;
        RECT 29.595 201.195 30.060 201.525 ;
        RECT 28.380 201.135 28.580 201.165 ;
        RECT 28.700 200.915 28.870 200.985 ;
        RECT 28.000 200.745 28.870 200.915 ;
        RECT 28.360 200.655 28.870 200.745 ;
        RECT 26.910 200.190 27.215 200.320 ;
        RECT 27.660 200.210 28.190 200.575 ;
        RECT 26.530 199.595 26.795 200.055 ;
        RECT 26.965 199.765 27.215 200.190 ;
        RECT 28.360 200.040 28.530 200.655 ;
        RECT 27.425 199.870 28.530 200.040 ;
        RECT 28.700 199.595 28.870 200.395 ;
        RECT 29.040 200.095 29.210 201.165 ;
        RECT 29.380 200.265 29.570 200.985 ;
        RECT 29.740 200.235 30.060 201.195 ;
        RECT 30.230 201.235 30.400 201.695 ;
        RECT 30.675 201.615 30.885 202.145 ;
        RECT 31.145 201.405 31.475 201.930 ;
        RECT 31.645 201.535 31.815 202.145 ;
        RECT 31.985 201.490 32.315 201.925 ;
        RECT 32.625 201.595 32.795 201.885 ;
        RECT 32.965 201.765 33.295 202.145 ;
        RECT 31.985 201.405 32.365 201.490 ;
        RECT 32.625 201.425 33.290 201.595 ;
        RECT 31.275 201.235 31.475 201.405 ;
        RECT 32.140 201.365 32.365 201.405 ;
        RECT 30.230 200.905 31.105 201.235 ;
        RECT 31.275 200.905 32.025 201.235 ;
        RECT 29.040 199.765 29.290 200.095 ;
        RECT 30.230 200.065 30.400 200.905 ;
        RECT 31.275 200.700 31.465 200.905 ;
        RECT 32.195 200.785 32.365 201.365 ;
        RECT 32.150 200.735 32.365 200.785 ;
        RECT 30.570 200.325 31.465 200.700 ;
        RECT 31.975 200.655 32.365 200.735 ;
        RECT 29.515 199.895 30.400 200.065 ;
        RECT 30.580 199.595 30.895 200.095 ;
        RECT 31.125 199.765 31.465 200.325 ;
        RECT 31.635 199.595 31.805 200.605 ;
        RECT 31.975 199.810 32.305 200.655 ;
        RECT 32.540 200.605 32.890 201.255 ;
        RECT 33.060 200.435 33.290 201.425 ;
        RECT 32.625 200.265 33.290 200.435 ;
        RECT 32.625 199.765 32.795 200.265 ;
        RECT 32.965 199.595 33.295 200.095 ;
        RECT 33.465 199.765 33.650 201.885 ;
        RECT 33.905 201.685 34.155 202.145 ;
        RECT 34.325 201.695 34.660 201.865 ;
        RECT 34.855 201.695 35.530 201.865 ;
        RECT 34.325 201.555 34.495 201.695 ;
        RECT 33.820 200.565 34.100 201.515 ;
        RECT 34.270 201.425 34.495 201.555 ;
        RECT 34.270 200.320 34.440 201.425 ;
        RECT 34.665 201.275 35.190 201.495 ;
        RECT 34.610 200.510 34.850 201.105 ;
        RECT 35.020 200.575 35.190 201.275 ;
        RECT 35.360 200.915 35.530 201.695 ;
        RECT 35.850 201.645 36.220 202.145 ;
        RECT 36.400 201.695 36.805 201.865 ;
        RECT 36.975 201.695 37.760 201.865 ;
        RECT 36.400 201.465 36.570 201.695 ;
        RECT 35.740 201.165 36.570 201.465 ;
        RECT 36.955 201.195 37.420 201.525 ;
        RECT 35.740 201.135 35.940 201.165 ;
        RECT 36.060 200.915 36.230 200.985 ;
        RECT 35.360 200.745 36.230 200.915 ;
        RECT 35.720 200.655 36.230 200.745 ;
        RECT 34.270 200.190 34.575 200.320 ;
        RECT 35.020 200.210 35.550 200.575 ;
        RECT 33.890 199.595 34.155 200.055 ;
        RECT 34.325 199.765 34.575 200.190 ;
        RECT 35.720 200.040 35.890 200.655 ;
        RECT 34.785 199.870 35.890 200.040 ;
        RECT 36.060 199.595 36.230 200.395 ;
        RECT 36.400 200.095 36.570 201.165 ;
        RECT 36.740 200.265 36.930 200.985 ;
        RECT 37.100 200.235 37.420 201.195 ;
        RECT 37.590 201.235 37.760 201.695 ;
        RECT 38.035 201.615 38.245 202.145 ;
        RECT 38.505 201.405 38.835 201.930 ;
        RECT 39.005 201.535 39.175 202.145 ;
        RECT 39.345 201.490 39.675 201.925 ;
        RECT 39.345 201.405 39.725 201.490 ;
        RECT 38.635 201.235 38.835 201.405 ;
        RECT 39.500 201.365 39.725 201.405 ;
        RECT 37.590 200.905 38.465 201.235 ;
        RECT 38.635 200.905 39.385 201.235 ;
        RECT 36.400 199.765 36.650 200.095 ;
        RECT 37.590 200.065 37.760 200.905 ;
        RECT 38.635 200.700 38.825 200.905 ;
        RECT 39.555 200.785 39.725 201.365 ;
        RECT 39.915 201.335 40.155 202.145 ;
        RECT 40.325 201.335 40.655 201.975 ;
        RECT 40.825 201.335 41.095 202.145 ;
        RECT 39.895 200.905 40.245 201.155 ;
        RECT 39.510 200.735 39.725 200.785 ;
        RECT 40.415 200.735 40.585 201.335 ;
        RECT 41.280 201.305 41.540 202.145 ;
        RECT 41.715 201.400 41.970 201.975 ;
        RECT 42.140 201.765 42.470 202.145 ;
        RECT 42.685 201.595 42.855 201.975 ;
        RECT 42.140 201.425 42.855 201.595 ;
        RECT 40.755 200.905 41.105 201.155 ;
        RECT 37.930 200.325 38.825 200.700 ;
        RECT 39.335 200.655 39.725 200.735 ;
        RECT 36.875 199.895 37.760 200.065 ;
        RECT 37.940 199.595 38.255 200.095 ;
        RECT 38.485 199.765 38.825 200.325 ;
        RECT 38.995 199.595 39.165 200.605 ;
        RECT 39.335 199.810 39.665 200.655 ;
        RECT 39.905 200.565 40.585 200.735 ;
        RECT 39.905 199.780 40.235 200.565 ;
        RECT 40.765 199.595 41.095 200.735 ;
        RECT 41.280 199.595 41.540 200.745 ;
        RECT 41.715 200.670 41.885 201.400 ;
        RECT 42.140 201.235 42.310 201.425 ;
        RECT 43.115 201.420 43.405 202.145 ;
        RECT 43.815 201.675 43.985 202.145 ;
        RECT 44.655 201.675 44.825 202.145 ;
        RECT 45.090 201.755 46.320 201.975 ;
        RECT 44.155 201.505 44.485 201.585 ;
        RECT 45.515 201.505 45.845 201.585 ;
        RECT 43.575 201.325 45.845 201.505 ;
        RECT 46.070 201.505 46.320 201.755 ;
        RECT 46.490 201.675 46.660 202.145 ;
        RECT 46.830 201.505 47.160 201.975 ;
        RECT 47.430 201.675 47.600 202.145 ;
        RECT 46.070 201.325 47.160 201.505 ;
        RECT 47.770 201.505 48.100 201.975 ;
        RECT 48.270 201.675 48.440 202.145 ;
        RECT 48.610 201.505 48.940 201.975 ;
        RECT 49.110 201.675 49.280 202.145 ;
        RECT 47.770 201.325 49.350 201.505 ;
        RECT 42.055 200.905 42.310 201.235 ;
        RECT 42.140 200.695 42.310 200.905 ;
        RECT 42.590 200.875 42.945 201.245 ;
        RECT 43.575 200.815 43.985 201.325 ;
        RECT 44.195 200.985 44.855 201.155 ;
        RECT 41.715 199.765 41.970 200.670 ;
        RECT 42.140 200.525 42.855 200.695 ;
        RECT 42.140 199.595 42.470 200.355 ;
        RECT 42.685 199.765 42.855 200.525 ;
        RECT 43.115 199.595 43.405 200.760 ;
        RECT 43.575 200.605 44.445 200.815 ;
        RECT 44.685 200.785 44.855 200.985 ;
        RECT 45.380 200.955 46.050 201.155 ;
        RECT 46.240 200.955 47.760 201.155 ;
        RECT 47.930 200.955 48.425 201.155 ;
        RECT 48.595 200.955 48.925 201.155 ;
        RECT 47.590 200.785 47.760 200.955 ;
        RECT 48.595 200.785 48.765 200.955 ;
        RECT 44.685 200.615 47.420 200.785 ;
        RECT 47.590 200.615 48.765 200.785 ;
        RECT 43.775 199.935 44.025 200.435 ;
        RECT 44.195 200.105 44.445 200.605 ;
        RECT 47.250 200.445 47.420 200.615 ;
        RECT 49.180 200.445 49.350 201.325 ;
        RECT 49.555 201.395 50.765 202.145 ;
        RECT 50.935 201.635 51.275 202.145 ;
        RECT 49.555 200.855 50.075 201.395 ;
        RECT 50.245 200.685 50.765 201.225 ;
        RECT 50.945 200.905 51.285 201.465 ;
        RECT 51.455 201.235 51.705 201.965 ;
        RECT 52.030 201.605 52.215 201.965 ;
        RECT 52.395 201.775 52.725 202.145 ;
        RECT 52.905 201.605 53.130 201.965 ;
        RECT 53.780 201.645 54.275 201.975 ;
        RECT 52.030 201.415 53.510 201.605 ;
        RECT 51.455 200.905 52.095 201.235 ;
        RECT 52.275 200.905 52.605 201.235 ;
        RECT 44.615 200.275 47.080 200.445 ;
        RECT 47.250 200.275 49.350 200.445 ;
        RECT 44.615 199.935 45.385 200.275 ;
        RECT 43.775 199.765 45.385 199.935 ;
        RECT 45.555 199.595 45.860 200.095 ;
        RECT 46.030 199.765 46.280 200.275 ;
        RECT 46.870 200.105 47.080 200.275 ;
        RECT 47.810 200.105 48.060 200.275 ;
        RECT 46.450 199.595 46.700 200.095 ;
        RECT 46.870 199.765 47.185 200.105 ;
        RECT 48.235 200.095 48.405 200.105 ;
        RECT 49.155 200.095 49.325 200.105 ;
        RECT 47.390 199.935 47.640 200.095 ;
        RECT 48.230 199.935 48.480 200.095 ;
        RECT 47.390 199.765 48.480 199.935 ;
        RECT 48.650 199.595 48.900 200.095 ;
        RECT 49.070 199.765 49.350 200.095 ;
        RECT 49.555 199.595 50.765 200.685 ;
        RECT 51.100 200.505 52.205 200.705 ;
        RECT 51.100 199.775 51.350 200.505 ;
        RECT 51.520 199.595 51.850 200.325 ;
        RECT 52.020 199.775 52.205 200.505 ;
        RECT 52.375 199.775 52.605 200.905 ;
        RECT 52.785 200.615 53.085 201.235 ;
        RECT 53.295 200.445 53.510 201.415 ;
        RECT 52.785 199.775 53.510 200.445 ;
        RECT 53.695 200.155 53.935 201.465 ;
        RECT 54.105 200.735 54.275 201.645 ;
        RECT 54.495 200.905 54.845 201.870 ;
        RECT 55.025 200.905 55.325 201.875 ;
        RECT 55.505 200.905 55.785 201.875 ;
        RECT 55.965 201.345 56.235 202.145 ;
        RECT 56.405 201.425 56.745 201.935 ;
        RECT 56.915 201.645 57.255 202.145 ;
        RECT 55.980 200.905 56.310 201.155 ;
        RECT 55.980 200.735 56.295 200.905 ;
        RECT 54.105 200.565 56.295 200.735 ;
        RECT 53.700 199.595 54.035 199.975 ;
        RECT 54.205 199.765 54.455 200.565 ;
        RECT 54.675 199.595 55.005 200.315 ;
        RECT 55.190 199.765 55.440 200.565 ;
        RECT 55.905 199.595 56.235 200.395 ;
        RECT 56.485 200.025 56.745 201.425 ;
        RECT 56.915 200.905 57.255 201.475 ;
        RECT 57.425 201.235 57.670 201.925 ;
        RECT 57.865 201.645 58.195 202.145 ;
        RECT 58.395 201.575 58.565 201.925 ;
        RECT 58.740 201.745 59.070 202.145 ;
        RECT 59.240 201.575 59.410 201.925 ;
        RECT 59.580 201.745 59.960 202.145 ;
        RECT 58.395 201.405 59.980 201.575 ;
        RECT 60.150 201.470 60.425 201.815 ;
        RECT 59.810 201.235 59.980 201.405 ;
        RECT 57.425 200.905 58.080 201.235 ;
        RECT 56.405 199.765 56.745 200.025 ;
        RECT 56.915 199.595 57.255 200.670 ;
        RECT 57.425 200.310 57.665 200.905 ;
        RECT 57.860 200.445 58.180 200.735 ;
        RECT 58.350 200.615 59.090 201.235 ;
        RECT 59.260 200.905 59.640 201.235 ;
        RECT 59.810 200.905 60.085 201.235 ;
        RECT 59.810 200.735 59.980 200.905 ;
        RECT 60.255 200.735 60.425 201.470 ;
        RECT 59.320 200.565 59.980 200.735 ;
        RECT 59.320 200.445 59.490 200.565 ;
        RECT 57.860 200.275 59.490 200.445 ;
        RECT 57.435 199.935 59.490 200.105 ;
        RECT 57.440 199.815 59.490 199.935 ;
        RECT 59.660 199.595 59.940 200.395 ;
        RECT 60.150 199.765 60.425 200.735 ;
        RECT 60.595 201.200 60.935 201.975 ;
        RECT 61.105 201.685 61.275 202.145 ;
        RECT 61.515 201.710 61.875 201.975 ;
        RECT 61.515 201.705 61.870 201.710 ;
        RECT 61.515 201.695 61.865 201.705 ;
        RECT 61.515 201.690 61.860 201.695 ;
        RECT 61.515 201.680 61.855 201.690 ;
        RECT 62.505 201.685 62.675 202.145 ;
        RECT 61.515 201.675 61.850 201.680 ;
        RECT 61.515 201.665 61.840 201.675 ;
        RECT 61.515 201.655 61.830 201.665 ;
        RECT 61.515 201.515 61.815 201.655 ;
        RECT 61.105 201.325 61.815 201.515 ;
        RECT 62.005 201.515 62.335 201.595 ;
        RECT 62.845 201.515 63.185 201.975 ;
        RECT 62.005 201.325 63.185 201.515 ;
        RECT 63.415 201.325 63.625 202.145 ;
        RECT 63.795 201.345 64.125 201.975 ;
        RECT 60.595 199.765 60.875 201.200 ;
        RECT 61.105 200.755 61.390 201.325 ;
        RECT 61.575 200.925 62.045 201.155 ;
        RECT 62.215 201.135 62.545 201.155 ;
        RECT 62.215 200.955 62.665 201.135 ;
        RECT 62.855 200.955 63.185 201.155 ;
        RECT 61.105 200.540 62.255 200.755 ;
        RECT 61.045 199.595 61.755 200.370 ;
        RECT 61.925 199.765 62.255 200.540 ;
        RECT 62.450 199.840 62.665 200.955 ;
        RECT 62.955 200.615 63.185 200.955 ;
        RECT 63.795 200.745 64.045 201.345 ;
        RECT 64.295 201.325 64.525 202.145 ;
        RECT 64.735 201.375 68.245 202.145 ;
        RECT 68.875 201.420 69.165 202.145 ;
        RECT 69.795 201.405 70.180 201.975 ;
        RECT 70.350 201.685 70.675 202.145 ;
        RECT 71.195 201.515 71.475 201.975 ;
        RECT 64.215 200.905 64.545 201.155 ;
        RECT 64.735 200.855 66.385 201.375 ;
        RECT 62.845 199.595 63.175 200.315 ;
        RECT 63.415 199.595 63.625 200.735 ;
        RECT 63.795 199.765 64.125 200.745 ;
        RECT 64.295 199.595 64.525 200.735 ;
        RECT 66.555 200.685 68.245 201.205 ;
        RECT 64.735 199.595 68.245 200.685 ;
        RECT 68.875 199.595 69.165 200.760 ;
        RECT 69.795 200.735 70.075 201.405 ;
        RECT 70.350 201.345 71.475 201.515 ;
        RECT 70.350 201.235 70.800 201.345 ;
        RECT 70.245 200.905 70.800 201.235 ;
        RECT 71.665 201.175 72.065 201.975 ;
        RECT 72.465 201.685 72.735 202.145 ;
        RECT 72.905 201.515 73.190 201.975 ;
        RECT 69.795 199.765 70.180 200.735 ;
        RECT 70.350 200.445 70.800 200.905 ;
        RECT 70.970 200.615 72.065 201.175 ;
        RECT 70.350 200.225 71.475 200.445 ;
        RECT 70.350 199.595 70.675 200.055 ;
        RECT 71.195 199.765 71.475 200.225 ;
        RECT 71.665 199.765 72.065 200.615 ;
        RECT 72.235 201.345 73.190 201.515 ;
        RECT 73.475 201.685 74.035 201.975 ;
        RECT 74.205 201.685 74.455 202.145 ;
        RECT 72.235 200.445 72.445 201.345 ;
        RECT 72.615 200.615 73.305 201.175 ;
        RECT 72.235 200.225 73.190 200.445 ;
        RECT 72.465 199.595 72.735 200.055 ;
        RECT 72.905 199.765 73.190 200.225 ;
        RECT 73.475 200.315 73.725 201.685 ;
        RECT 75.075 201.515 75.405 201.875 ;
        RECT 76.480 201.665 76.780 202.145 ;
        RECT 74.015 201.325 75.405 201.515 ;
        RECT 76.950 201.495 77.210 201.950 ;
        RECT 77.380 201.665 77.640 202.145 ;
        RECT 77.810 201.495 78.070 201.950 ;
        RECT 78.240 201.665 78.500 202.145 ;
        RECT 78.670 201.495 78.930 201.950 ;
        RECT 79.100 201.665 79.360 202.145 ;
        RECT 79.530 201.495 79.790 201.950 ;
        RECT 79.960 201.620 80.220 202.145 ;
        RECT 76.480 201.325 79.790 201.495 ;
        RECT 74.015 201.235 74.185 201.325 ;
        RECT 73.895 200.905 74.185 201.235 ;
        RECT 74.355 200.905 74.695 201.155 ;
        RECT 74.915 200.905 75.590 201.155 ;
        RECT 74.015 200.655 74.185 200.905 ;
        RECT 74.015 200.485 74.955 200.655 ;
        RECT 75.325 200.545 75.590 200.905 ;
        RECT 76.480 200.735 77.450 201.325 ;
        RECT 80.390 201.155 80.640 201.965 ;
        RECT 80.820 201.685 81.065 202.145 ;
        RECT 77.620 200.905 80.640 201.155 ;
        RECT 80.810 200.905 81.125 201.515 ;
        RECT 81.355 201.325 81.565 202.145 ;
        RECT 81.735 201.345 82.065 201.975 ;
        RECT 76.480 200.495 79.790 200.735 ;
        RECT 73.475 199.765 73.935 200.315 ;
        RECT 74.125 199.595 74.455 200.315 ;
        RECT 74.655 199.935 74.955 200.485 ;
        RECT 75.125 199.595 75.405 200.265 ;
        RECT 76.485 199.595 76.780 200.325 ;
        RECT 76.950 199.770 77.210 200.495 ;
        RECT 77.380 199.595 77.640 200.325 ;
        RECT 77.810 199.770 78.070 200.495 ;
        RECT 78.240 199.595 78.500 200.325 ;
        RECT 78.670 199.770 78.930 200.495 ;
        RECT 79.100 199.595 79.360 200.325 ;
        RECT 79.530 199.770 79.790 200.495 ;
        RECT 79.960 199.595 80.220 200.705 ;
        RECT 80.390 199.770 80.640 200.905 ;
        RECT 81.735 200.745 81.985 201.345 ;
        RECT 82.235 201.325 82.465 202.145 ;
        RECT 82.790 201.515 83.075 201.975 ;
        RECT 83.245 201.685 83.515 202.145 ;
        RECT 82.790 201.345 83.745 201.515 ;
        RECT 82.155 200.905 82.485 201.155 ;
        RECT 80.820 199.595 81.115 200.705 ;
        RECT 81.355 199.595 81.565 200.735 ;
        RECT 81.735 199.765 82.065 200.745 ;
        RECT 82.235 199.595 82.465 200.735 ;
        RECT 82.675 200.615 83.365 201.175 ;
        RECT 83.535 200.445 83.745 201.345 ;
        RECT 82.790 200.225 83.745 200.445 ;
        RECT 83.915 201.175 84.315 201.975 ;
        RECT 84.505 201.515 84.785 201.975 ;
        RECT 85.305 201.685 85.630 202.145 ;
        RECT 84.505 201.345 85.630 201.515 ;
        RECT 85.800 201.405 86.185 201.975 ;
        RECT 87.365 201.595 87.535 201.885 ;
        RECT 87.705 201.765 88.035 202.145 ;
        RECT 87.365 201.425 88.030 201.595 ;
        RECT 85.180 201.235 85.630 201.345 ;
        RECT 83.915 200.615 85.010 201.175 ;
        RECT 85.180 200.905 85.735 201.235 ;
        RECT 82.790 199.765 83.075 200.225 ;
        RECT 83.245 199.595 83.515 200.055 ;
        RECT 83.915 199.765 84.315 200.615 ;
        RECT 85.180 200.445 85.630 200.905 ;
        RECT 85.905 200.735 86.185 201.405 ;
        RECT 84.505 200.225 85.630 200.445 ;
        RECT 84.505 199.765 84.785 200.225 ;
        RECT 85.305 199.595 85.630 200.055 ;
        RECT 85.800 199.765 86.185 200.735 ;
        RECT 87.280 200.605 87.630 201.255 ;
        RECT 87.800 200.435 88.030 201.425 ;
        RECT 87.365 200.265 88.030 200.435 ;
        RECT 87.365 199.765 87.535 200.265 ;
        RECT 87.705 199.595 88.035 200.095 ;
        RECT 88.205 199.765 88.390 201.885 ;
        RECT 88.645 201.685 88.895 202.145 ;
        RECT 89.065 201.695 89.400 201.865 ;
        RECT 89.595 201.695 90.270 201.865 ;
        RECT 89.065 201.555 89.235 201.695 ;
        RECT 88.560 200.565 88.840 201.515 ;
        RECT 89.010 201.425 89.235 201.555 ;
        RECT 89.010 200.320 89.180 201.425 ;
        RECT 89.405 201.275 89.930 201.495 ;
        RECT 89.350 200.510 89.590 201.105 ;
        RECT 89.760 200.575 89.930 201.275 ;
        RECT 90.100 200.915 90.270 201.695 ;
        RECT 90.590 201.645 90.960 202.145 ;
        RECT 91.140 201.695 91.545 201.865 ;
        RECT 91.715 201.695 92.500 201.865 ;
        RECT 91.140 201.465 91.310 201.695 ;
        RECT 90.480 201.165 91.310 201.465 ;
        RECT 91.695 201.195 92.160 201.525 ;
        RECT 90.480 201.135 90.680 201.165 ;
        RECT 90.800 200.915 90.970 200.985 ;
        RECT 90.100 200.745 90.970 200.915 ;
        RECT 90.460 200.655 90.970 200.745 ;
        RECT 89.010 200.190 89.315 200.320 ;
        RECT 89.760 200.210 90.290 200.575 ;
        RECT 88.630 199.595 88.895 200.055 ;
        RECT 89.065 199.765 89.315 200.190 ;
        RECT 90.460 200.040 90.630 200.655 ;
        RECT 89.525 199.870 90.630 200.040 ;
        RECT 90.800 199.595 90.970 200.395 ;
        RECT 91.140 200.095 91.310 201.165 ;
        RECT 91.480 200.265 91.670 200.985 ;
        RECT 91.840 200.235 92.160 201.195 ;
        RECT 92.330 201.235 92.500 201.695 ;
        RECT 92.775 201.615 92.985 202.145 ;
        RECT 93.245 201.405 93.575 201.930 ;
        RECT 93.745 201.535 93.915 202.145 ;
        RECT 94.085 201.490 94.415 201.925 ;
        RECT 94.085 201.405 94.465 201.490 ;
        RECT 94.635 201.420 94.925 202.145 ;
        RECT 93.375 201.235 93.575 201.405 ;
        RECT 94.240 201.365 94.465 201.405 ;
        RECT 92.330 200.905 93.205 201.235 ;
        RECT 93.375 200.905 94.125 201.235 ;
        RECT 91.140 199.765 91.390 200.095 ;
        RECT 92.330 200.065 92.500 200.905 ;
        RECT 93.375 200.700 93.565 200.905 ;
        RECT 94.295 200.785 94.465 201.365 ;
        RECT 94.250 200.735 94.465 200.785 ;
        RECT 95.100 201.405 95.355 201.975 ;
        RECT 95.525 201.745 95.855 202.145 ;
        RECT 96.280 201.610 96.810 201.975 ;
        RECT 96.280 201.575 96.455 201.610 ;
        RECT 95.525 201.405 96.455 201.575 ;
        RECT 97.000 201.465 97.275 201.975 ;
        RECT 92.670 200.325 93.565 200.700 ;
        RECT 94.075 200.655 94.465 200.735 ;
        RECT 91.615 199.895 92.500 200.065 ;
        RECT 92.680 199.595 92.995 200.095 ;
        RECT 93.225 199.765 93.565 200.325 ;
        RECT 93.735 199.595 93.905 200.605 ;
        RECT 94.075 199.810 94.405 200.655 ;
        RECT 94.635 199.595 94.925 200.760 ;
        RECT 95.100 200.735 95.270 201.405 ;
        RECT 95.525 201.235 95.695 201.405 ;
        RECT 95.440 200.905 95.695 201.235 ;
        RECT 95.920 200.905 96.115 201.235 ;
        RECT 95.100 199.765 95.435 200.735 ;
        RECT 95.605 199.595 95.775 200.735 ;
        RECT 95.945 199.935 96.115 200.905 ;
        RECT 96.285 200.275 96.455 201.405 ;
        RECT 96.625 200.615 96.795 201.415 ;
        RECT 96.995 201.295 97.275 201.465 ;
        RECT 97.000 200.815 97.275 201.295 ;
        RECT 97.445 200.615 97.635 201.975 ;
        RECT 97.815 201.610 98.325 202.145 ;
        RECT 98.545 201.335 98.790 201.940 ;
        RECT 99.235 201.405 99.745 201.975 ;
        RECT 99.915 201.585 100.085 202.145 ;
        RECT 100.290 201.575 100.620 201.975 ;
        RECT 100.795 201.745 101.125 202.145 ;
        RECT 101.360 201.765 102.745 201.975 ;
        RECT 101.360 201.575 101.690 201.765 ;
        RECT 100.290 201.405 101.690 201.575 ;
        RECT 101.860 201.405 102.285 201.595 ;
        RECT 102.455 201.495 102.745 201.765 ;
        RECT 97.835 201.165 99.065 201.335 ;
        RECT 96.625 200.445 97.635 200.615 ;
        RECT 97.805 200.600 98.555 200.790 ;
        RECT 96.285 200.105 97.410 200.275 ;
        RECT 97.805 199.935 97.975 200.600 ;
        RECT 98.725 200.355 99.065 201.165 ;
        RECT 95.945 199.765 97.975 199.935 ;
        RECT 98.145 199.595 98.315 200.355 ;
        RECT 98.550 199.945 99.065 200.355 ;
        RECT 99.235 200.735 99.410 201.405 ;
        RECT 99.595 201.155 99.785 201.235 ;
        RECT 100.155 201.155 100.325 201.235 ;
        RECT 99.595 200.905 99.960 201.155 ;
        RECT 100.155 200.905 100.405 201.155 ;
        RECT 100.615 200.905 100.960 201.235 ;
        RECT 99.790 200.735 99.960 200.905 ;
        RECT 99.235 199.775 99.620 200.735 ;
        RECT 99.790 200.565 100.465 200.735 ;
        RECT 99.835 199.595 100.125 200.395 ;
        RECT 100.295 199.935 100.465 200.565 ;
        RECT 100.635 200.105 100.960 200.905 ;
        RECT 101.130 200.570 101.405 201.235 ;
        RECT 101.590 200.570 101.945 201.235 ;
        RECT 102.115 200.395 102.285 201.405 ;
        RECT 102.925 201.420 103.255 201.930 ;
        RECT 103.425 201.745 103.755 202.145 ;
        RECT 104.805 201.575 105.135 201.915 ;
        RECT 105.305 201.745 105.635 202.145 ;
        RECT 102.470 200.905 102.745 201.235 ;
        RECT 101.330 200.145 102.285 200.395 ;
        RECT 101.330 199.935 101.660 200.145 ;
        RECT 100.295 199.765 101.660 199.935 ;
        RECT 102.455 199.595 102.745 200.735 ;
        RECT 102.925 200.655 103.115 201.420 ;
        RECT 103.425 201.405 105.790 201.575 ;
        RECT 103.425 201.235 103.595 201.405 ;
        RECT 103.285 200.905 103.595 201.235 ;
        RECT 103.765 200.905 104.070 201.235 ;
        RECT 102.925 199.805 103.255 200.655 ;
        RECT 103.425 199.595 103.675 200.735 ;
        RECT 103.855 200.575 104.070 200.905 ;
        RECT 104.245 200.575 104.530 201.235 ;
        RECT 104.725 200.575 104.990 201.235 ;
        RECT 105.205 200.575 105.450 201.235 ;
        RECT 105.620 200.405 105.790 201.405 ;
        RECT 106.175 201.325 106.405 202.145 ;
        RECT 106.575 201.345 106.905 201.975 ;
        RECT 106.155 200.905 106.485 201.155 ;
        RECT 106.655 200.745 106.905 201.345 ;
        RECT 107.075 201.325 107.285 202.145 ;
        RECT 107.515 201.375 111.025 202.145 ;
        RECT 107.515 200.855 109.165 201.375 ;
        RECT 111.470 201.335 111.715 201.940 ;
        RECT 111.935 201.610 112.445 202.145 ;
        RECT 103.865 200.235 105.155 200.405 ;
        RECT 103.865 199.815 104.115 200.235 ;
        RECT 104.345 199.595 104.675 200.065 ;
        RECT 104.905 199.815 105.155 200.235 ;
        RECT 105.335 200.235 105.790 200.405 ;
        RECT 105.335 199.805 105.665 200.235 ;
        RECT 106.175 199.595 106.405 200.735 ;
        RECT 106.575 199.765 106.905 200.745 ;
        RECT 107.075 199.595 107.285 200.735 ;
        RECT 109.335 200.685 111.025 201.205 ;
        RECT 107.515 199.595 111.025 200.685 ;
        RECT 111.195 201.165 112.425 201.335 ;
        RECT 111.195 200.355 111.535 201.165 ;
        RECT 111.705 200.600 112.455 200.790 ;
        RECT 111.195 199.945 111.710 200.355 ;
        RECT 111.945 199.595 112.115 200.355 ;
        RECT 112.285 199.935 112.455 200.600 ;
        RECT 112.625 200.615 112.815 201.975 ;
        RECT 112.985 201.125 113.260 201.975 ;
        RECT 113.450 201.610 113.980 201.975 ;
        RECT 114.405 201.745 114.735 202.145 ;
        RECT 113.805 201.575 113.980 201.610 ;
        RECT 112.985 200.955 113.265 201.125 ;
        RECT 112.985 200.815 113.260 200.955 ;
        RECT 113.465 200.615 113.635 201.415 ;
        RECT 112.625 200.445 113.635 200.615 ;
        RECT 113.805 201.405 114.735 201.575 ;
        RECT 114.905 201.405 115.160 201.975 ;
        RECT 113.805 200.275 113.975 201.405 ;
        RECT 114.565 201.235 114.735 201.405 ;
        RECT 112.850 200.105 113.975 200.275 ;
        RECT 114.145 200.905 114.340 201.235 ;
        RECT 114.565 200.905 114.820 201.235 ;
        RECT 114.145 199.935 114.315 200.905 ;
        RECT 114.990 200.735 115.160 201.405 ;
        RECT 115.335 201.375 118.845 202.145 ;
        RECT 119.015 201.395 120.225 202.145 ;
        RECT 120.395 201.420 120.685 202.145 ;
        RECT 120.855 201.600 126.200 202.145 ;
        RECT 126.375 201.600 131.720 202.145 ;
        RECT 131.895 201.600 137.240 202.145 ;
        RECT 137.415 201.600 142.760 202.145 ;
        RECT 115.335 200.855 116.985 201.375 ;
        RECT 112.285 199.765 114.315 199.935 ;
        RECT 114.485 199.595 114.655 200.735 ;
        RECT 114.825 199.765 115.160 200.735 ;
        RECT 117.155 200.685 118.845 201.205 ;
        RECT 119.015 200.855 119.535 201.395 ;
        RECT 119.705 200.685 120.225 201.225 ;
        RECT 122.440 200.770 122.780 201.600 ;
        RECT 115.335 199.595 118.845 200.685 ;
        RECT 119.015 199.595 120.225 200.685 ;
        RECT 120.395 199.595 120.685 200.760 ;
        RECT 124.260 200.030 124.610 201.280 ;
        RECT 127.960 200.770 128.300 201.600 ;
        RECT 129.780 200.030 130.130 201.280 ;
        RECT 133.480 200.770 133.820 201.600 ;
        RECT 135.300 200.030 135.650 201.280 ;
        RECT 139.000 200.770 139.340 201.600 ;
        RECT 142.935 201.375 145.525 202.145 ;
        RECT 145.695 201.395 146.905 202.145 ;
        RECT 140.820 200.030 141.170 201.280 ;
        RECT 142.935 200.855 144.145 201.375 ;
        RECT 144.315 200.685 145.525 201.205 ;
        RECT 120.855 199.595 126.200 200.030 ;
        RECT 126.375 199.595 131.720 200.030 ;
        RECT 131.895 199.595 137.240 200.030 ;
        RECT 137.415 199.595 142.760 200.030 ;
        RECT 142.935 199.595 145.525 200.685 ;
        RECT 145.695 200.685 146.215 201.225 ;
        RECT 146.385 200.855 146.905 201.395 ;
        RECT 145.695 199.595 146.905 200.685 ;
        RECT 17.270 199.425 146.990 199.595 ;
        RECT 17.355 198.335 18.565 199.425 ;
        RECT 18.735 198.335 21.325 199.425 ;
        RECT 21.585 198.755 21.755 199.255 ;
        RECT 21.925 198.925 22.255 199.425 ;
        RECT 21.585 198.585 22.250 198.755 ;
        RECT 17.355 197.625 17.875 198.165 ;
        RECT 18.045 197.795 18.565 198.335 ;
        RECT 18.735 197.645 19.945 198.165 ;
        RECT 20.115 197.815 21.325 198.335 ;
        RECT 21.500 197.765 21.850 198.415 ;
        RECT 17.355 196.875 18.565 197.625 ;
        RECT 18.735 196.875 21.325 197.645 ;
        RECT 22.020 197.595 22.250 198.585 ;
        RECT 21.585 197.425 22.250 197.595 ;
        RECT 21.585 197.135 21.755 197.425 ;
        RECT 21.925 196.875 22.255 197.255 ;
        RECT 22.425 197.135 22.610 199.255 ;
        RECT 22.850 198.965 23.115 199.425 ;
        RECT 23.285 198.830 23.535 199.255 ;
        RECT 23.745 198.980 24.850 199.150 ;
        RECT 23.230 198.700 23.535 198.830 ;
        RECT 22.780 197.505 23.060 198.455 ;
        RECT 23.230 197.595 23.400 198.700 ;
        RECT 23.570 197.915 23.810 198.510 ;
        RECT 23.980 198.445 24.510 198.810 ;
        RECT 23.980 197.745 24.150 198.445 ;
        RECT 24.680 198.365 24.850 198.980 ;
        RECT 25.020 198.625 25.190 199.425 ;
        RECT 25.360 198.925 25.610 199.255 ;
        RECT 25.835 198.955 26.720 199.125 ;
        RECT 24.680 198.275 25.190 198.365 ;
        RECT 23.230 197.465 23.455 197.595 ;
        RECT 23.625 197.525 24.150 197.745 ;
        RECT 24.320 198.105 25.190 198.275 ;
        RECT 22.865 196.875 23.115 197.335 ;
        RECT 23.285 197.325 23.455 197.465 ;
        RECT 24.320 197.325 24.490 198.105 ;
        RECT 25.020 198.035 25.190 198.105 ;
        RECT 24.700 197.855 24.900 197.885 ;
        RECT 25.360 197.855 25.530 198.925 ;
        RECT 25.700 198.035 25.890 198.755 ;
        RECT 24.700 197.555 25.530 197.855 ;
        RECT 26.060 197.825 26.380 198.785 ;
        RECT 23.285 197.155 23.620 197.325 ;
        RECT 23.815 197.155 24.490 197.325 ;
        RECT 24.810 196.875 25.180 197.375 ;
        RECT 25.360 197.325 25.530 197.555 ;
        RECT 25.915 197.495 26.380 197.825 ;
        RECT 26.550 198.115 26.720 198.955 ;
        RECT 26.900 198.925 27.215 199.425 ;
        RECT 27.445 198.695 27.785 199.255 ;
        RECT 26.890 198.320 27.785 198.695 ;
        RECT 27.955 198.415 28.125 199.425 ;
        RECT 27.595 198.115 27.785 198.320 ;
        RECT 28.295 198.365 28.625 199.210 ;
        RECT 28.295 198.285 28.685 198.365 ;
        RECT 28.855 198.285 29.135 199.425 ;
        RECT 28.470 198.235 28.685 198.285 ;
        RECT 29.305 198.275 29.635 199.255 ;
        RECT 29.805 198.285 30.065 199.425 ;
        RECT 26.550 197.785 27.425 198.115 ;
        RECT 27.595 197.785 28.345 198.115 ;
        RECT 26.550 197.325 26.720 197.785 ;
        RECT 27.595 197.615 27.795 197.785 ;
        RECT 28.515 197.655 28.685 198.235 ;
        RECT 28.865 197.845 29.200 198.115 ;
        RECT 29.370 197.675 29.540 198.275 ;
        RECT 30.235 198.260 30.525 199.425 ;
        RECT 29.710 197.865 30.045 198.115 ;
        RECT 28.460 197.615 28.685 197.655 ;
        RECT 25.360 197.155 25.765 197.325 ;
        RECT 25.935 197.155 26.720 197.325 ;
        RECT 26.995 196.875 27.205 197.405 ;
        RECT 27.465 197.090 27.795 197.615 ;
        RECT 28.305 197.530 28.685 197.615 ;
        RECT 27.965 196.875 28.135 197.485 ;
        RECT 28.305 197.095 28.635 197.530 ;
        RECT 28.855 196.875 29.165 197.675 ;
        RECT 29.370 197.045 30.065 197.675 ;
        RECT 30.235 196.875 30.525 197.600 ;
        RECT 30.705 197.055 30.965 199.245 ;
        RECT 31.135 198.695 31.475 199.425 ;
        RECT 31.655 198.515 31.925 199.245 ;
        RECT 31.155 198.295 31.925 198.515 ;
        RECT 32.105 198.535 32.335 199.245 ;
        RECT 32.505 198.715 32.835 199.425 ;
        RECT 33.005 198.535 33.265 199.245 ;
        RECT 32.105 198.295 33.265 198.535 ;
        RECT 33.640 198.455 34.030 198.630 ;
        RECT 34.515 198.625 34.845 199.425 ;
        RECT 35.015 198.635 35.550 199.255 ;
        RECT 31.155 197.625 31.445 198.295 ;
        RECT 33.640 198.285 35.065 198.455 ;
        RECT 31.625 197.805 32.090 198.115 ;
        RECT 32.270 197.805 32.795 198.115 ;
        RECT 31.155 197.425 32.385 197.625 ;
        RECT 31.225 196.875 31.895 197.245 ;
        RECT 32.075 197.055 32.385 197.425 ;
        RECT 32.565 197.165 32.795 197.805 ;
        RECT 32.975 197.785 33.275 198.115 ;
        RECT 32.975 196.875 33.265 197.605 ;
        RECT 33.515 197.555 33.870 198.115 ;
        RECT 34.040 197.385 34.210 198.285 ;
        RECT 34.380 197.555 34.645 198.115 ;
        RECT 34.895 197.785 35.065 198.285 ;
        RECT 35.235 197.615 35.550 198.635 ;
        RECT 33.620 196.875 33.860 197.385 ;
        RECT 34.040 197.055 34.320 197.385 ;
        RECT 34.550 196.875 34.765 197.385 ;
        RECT 34.935 197.045 35.550 197.615 ;
        RECT 35.755 198.555 36.030 199.255 ;
        RECT 36.200 198.880 36.455 199.425 ;
        RECT 36.625 198.915 37.105 199.255 ;
        RECT 37.280 198.870 37.885 199.425 ;
        RECT 37.270 198.770 37.885 198.870 ;
        RECT 37.270 198.745 37.455 198.770 ;
        RECT 35.755 197.525 35.925 198.555 ;
        RECT 36.200 198.425 36.955 198.675 ;
        RECT 37.125 198.500 37.455 198.745 ;
        RECT 36.200 198.390 36.970 198.425 ;
        RECT 36.200 198.380 36.985 198.390 ;
        RECT 36.095 198.365 36.990 198.380 ;
        RECT 36.095 198.350 37.010 198.365 ;
        RECT 36.095 198.340 37.030 198.350 ;
        RECT 36.095 198.330 37.055 198.340 ;
        RECT 36.095 198.300 37.125 198.330 ;
        RECT 36.095 198.270 37.145 198.300 ;
        RECT 36.095 198.240 37.165 198.270 ;
        RECT 36.095 198.215 37.195 198.240 ;
        RECT 36.095 198.180 37.230 198.215 ;
        RECT 36.095 198.175 37.260 198.180 ;
        RECT 36.095 197.780 36.325 198.175 ;
        RECT 36.870 198.170 37.260 198.175 ;
        RECT 36.895 198.160 37.260 198.170 ;
        RECT 36.910 198.155 37.260 198.160 ;
        RECT 36.925 198.150 37.260 198.155 ;
        RECT 37.625 198.150 37.885 198.600 ;
        RECT 38.985 198.445 39.315 199.255 ;
        RECT 39.485 198.625 39.725 199.425 ;
        RECT 38.985 198.275 39.700 198.445 ;
        RECT 36.925 198.145 37.885 198.150 ;
        RECT 36.935 198.135 37.885 198.145 ;
        RECT 36.945 198.130 37.885 198.135 ;
        RECT 36.955 198.120 37.885 198.130 ;
        RECT 36.960 198.110 37.885 198.120 ;
        RECT 36.965 198.105 37.885 198.110 ;
        RECT 36.975 198.090 37.885 198.105 ;
        RECT 36.980 198.075 37.885 198.090 ;
        RECT 36.990 198.050 37.885 198.075 ;
        RECT 36.495 197.580 36.825 198.005 ;
        RECT 36.575 197.555 36.825 197.580 ;
        RECT 35.755 197.045 36.015 197.525 ;
        RECT 36.185 196.875 36.435 197.415 ;
        RECT 36.605 197.095 36.825 197.555 ;
        RECT 36.995 197.980 37.885 198.050 ;
        RECT 36.995 197.255 37.165 197.980 ;
        RECT 38.980 197.865 39.360 198.105 ;
        RECT 39.530 198.035 39.700 198.275 ;
        RECT 39.905 198.405 40.075 199.255 ;
        RECT 40.245 198.625 40.575 199.425 ;
        RECT 40.745 198.405 40.915 199.255 ;
        RECT 39.905 198.235 40.915 198.405 ;
        RECT 41.085 198.275 41.415 199.425 ;
        RECT 42.220 198.455 42.520 198.650 ;
        RECT 42.690 198.625 42.945 199.425 ;
        RECT 43.145 198.795 43.475 199.255 ;
        RECT 43.645 198.965 44.220 199.425 ;
        RECT 44.390 198.795 44.745 199.255 ;
        RECT 43.145 198.625 44.745 198.795 ;
        RECT 42.220 198.285 43.470 198.455 ;
        RECT 40.420 198.065 40.915 198.235 ;
        RECT 39.530 197.865 40.030 198.035 ;
        RECT 40.415 197.895 40.915 198.065 ;
        RECT 37.335 197.425 37.885 197.810 ;
        RECT 39.530 197.695 39.700 197.865 ;
        RECT 40.420 197.695 40.915 197.895 ;
        RECT 39.065 197.525 39.700 197.695 ;
        RECT 39.905 197.525 40.915 197.695 ;
        RECT 36.995 197.085 37.885 197.255 ;
        RECT 39.065 197.045 39.235 197.525 ;
        RECT 39.415 196.875 39.655 197.355 ;
        RECT 39.905 197.045 40.075 197.525 ;
        RECT 40.245 196.875 40.575 197.355 ;
        RECT 40.745 197.045 40.915 197.525 ;
        RECT 41.085 196.875 41.415 197.675 ;
        RECT 42.220 197.630 42.390 198.285 ;
        RECT 42.565 197.785 42.910 198.115 ;
        RECT 43.140 197.865 43.470 198.285 ;
        RECT 43.640 197.695 43.920 198.625 ;
        RECT 44.100 198.405 44.290 198.445 ;
        RECT 44.095 198.235 44.290 198.405 ;
        RECT 44.470 198.285 44.745 198.625 ;
        RECT 44.915 198.285 45.245 199.425 ;
        RECT 45.600 198.455 45.990 198.630 ;
        RECT 46.475 198.625 46.805 199.425 ;
        RECT 46.975 198.635 47.510 199.255 ;
        RECT 45.600 198.285 47.025 198.455 ;
        RECT 44.555 198.235 44.725 198.285 ;
        RECT 44.100 198.065 44.290 198.235 ;
        RECT 44.100 197.865 45.245 198.065 ;
        RECT 42.220 197.300 42.455 197.630 ;
        RECT 42.625 196.875 42.955 197.615 ;
        RECT 43.190 197.255 43.465 197.695 ;
        RECT 43.640 197.595 43.965 197.695 ;
        RECT 43.635 197.425 43.965 197.595 ;
        RECT 44.135 197.485 45.245 197.695 ;
        RECT 45.475 197.555 45.830 198.115 ;
        RECT 44.135 197.255 44.385 197.485 ;
        RECT 43.190 197.045 44.385 197.255 ;
        RECT 44.555 196.875 44.725 197.315 ;
        RECT 44.895 197.045 45.245 197.485 ;
        RECT 46.000 197.385 46.170 198.285 ;
        RECT 46.340 197.555 46.605 198.115 ;
        RECT 46.855 197.785 47.025 198.285 ;
        RECT 47.195 197.615 47.510 198.635 ;
        RECT 48.645 198.475 48.920 199.245 ;
        RECT 49.090 198.815 49.420 199.245 ;
        RECT 49.590 198.985 49.785 199.425 ;
        RECT 49.965 198.815 50.295 199.245 ;
        RECT 49.090 198.645 50.295 198.815 ;
        RECT 50.675 198.755 50.955 199.425 ;
        RECT 48.645 198.285 49.230 198.475 ;
        RECT 49.400 198.315 50.295 198.645 ;
        RECT 51.125 198.535 51.425 199.085 ;
        RECT 51.625 198.705 51.955 199.425 ;
        RECT 52.145 198.705 52.605 199.255 ;
        RECT 53.075 198.785 53.405 199.215 ;
        RECT 45.580 196.875 45.820 197.385 ;
        RECT 46.000 197.055 46.280 197.385 ;
        RECT 46.510 196.875 46.725 197.385 ;
        RECT 46.895 197.045 47.510 197.615 ;
        RECT 48.645 197.465 48.885 198.115 ;
        RECT 49.055 197.615 49.230 198.285 ;
        RECT 50.490 198.115 50.755 198.475 ;
        RECT 51.125 198.365 52.065 198.535 ;
        RECT 51.895 198.115 52.065 198.365 ;
        RECT 49.400 197.785 49.815 198.115 ;
        RECT 49.995 197.785 50.290 198.115 ;
        RECT 50.490 197.865 51.165 198.115 ;
        RECT 51.385 197.865 51.725 198.115 ;
        RECT 51.895 197.785 52.185 198.115 ;
        RECT 49.055 197.435 49.385 197.615 ;
        RECT 48.660 196.875 48.990 197.265 ;
        RECT 49.160 197.055 49.385 197.435 ;
        RECT 49.585 197.165 49.815 197.785 ;
        RECT 51.895 197.695 52.065 197.785 ;
        RECT 49.995 196.875 50.295 197.605 ;
        RECT 50.675 197.505 52.065 197.695 ;
        RECT 50.675 197.145 51.005 197.505 ;
        RECT 52.355 197.335 52.605 198.705 ;
        RECT 52.950 198.615 53.405 198.785 ;
        RECT 53.585 198.785 53.835 199.205 ;
        RECT 54.065 198.955 54.395 199.425 ;
        RECT 54.625 198.785 54.875 199.205 ;
        RECT 53.585 198.615 54.875 198.785 ;
        RECT 52.950 197.615 53.120 198.615 ;
        RECT 53.290 197.785 53.535 198.445 ;
        RECT 53.750 197.785 54.015 198.445 ;
        RECT 54.210 197.785 54.495 198.445 ;
        RECT 54.670 198.115 54.885 198.445 ;
        RECT 55.065 198.285 55.315 199.425 ;
        RECT 55.485 198.365 55.815 199.215 ;
        RECT 54.670 197.785 54.975 198.115 ;
        RECT 55.145 197.785 55.455 198.115 ;
        RECT 55.145 197.615 55.315 197.785 ;
        RECT 52.950 197.445 55.315 197.615 ;
        RECT 55.625 197.600 55.815 198.365 ;
        RECT 55.995 198.260 56.285 199.425 ;
        RECT 56.515 198.285 56.725 199.425 ;
        RECT 56.895 198.275 57.225 199.255 ;
        RECT 57.395 198.285 57.625 199.425 ;
        RECT 57.835 198.925 58.095 199.255 ;
        RECT 58.405 199.045 58.735 199.425 ;
        RECT 51.625 196.875 51.875 197.335 ;
        RECT 52.045 197.045 52.605 197.335 ;
        RECT 53.105 196.875 53.435 197.275 ;
        RECT 53.605 197.105 53.935 197.445 ;
        RECT 54.985 196.875 55.315 197.275 ;
        RECT 55.485 197.090 55.815 197.600 ;
        RECT 55.995 196.875 56.285 197.600 ;
        RECT 56.515 196.875 56.725 197.695 ;
        RECT 56.895 197.675 57.145 198.275 ;
        RECT 57.835 198.245 58.005 198.925 ;
        RECT 58.975 198.875 59.165 199.255 ;
        RECT 59.415 199.045 59.745 199.425 ;
        RECT 59.955 198.875 60.125 199.255 ;
        RECT 60.320 199.045 60.650 199.425 ;
        RECT 60.910 198.875 61.080 199.255 ;
        RECT 61.505 199.045 61.835 199.425 ;
        RECT 58.175 198.415 58.525 198.745 ;
        RECT 58.975 198.705 59.715 198.875 ;
        RECT 58.795 198.365 59.375 198.535 ;
        RECT 58.795 198.245 58.965 198.365 ;
        RECT 57.315 197.865 57.645 198.115 ;
        RECT 57.835 198.075 58.965 198.245 ;
        RECT 59.545 198.195 59.715 198.705 ;
        RECT 56.895 197.045 57.225 197.675 ;
        RECT 57.395 196.875 57.625 197.695 ;
        RECT 57.835 197.375 58.005 198.075 ;
        RECT 59.145 198.025 59.715 198.195 ;
        RECT 59.885 198.705 61.835 198.875 ;
        RECT 58.355 197.735 58.975 197.905 ;
        RECT 58.355 197.555 58.565 197.735 ;
        RECT 59.145 197.545 59.315 198.025 ;
        RECT 59.885 197.715 60.055 198.705 ;
        RECT 60.645 198.115 60.830 198.425 ;
        RECT 61.100 198.115 61.295 198.425 ;
        RECT 57.835 197.045 58.095 197.375 ;
        RECT 58.405 196.875 58.735 197.255 ;
        RECT 58.915 197.215 59.315 197.545 ;
        RECT 59.505 197.385 60.055 197.715 ;
        RECT 60.225 197.215 60.395 198.115 ;
        RECT 58.915 197.045 60.395 197.215 ;
        RECT 60.645 197.785 60.875 198.115 ;
        RECT 61.100 197.785 61.355 198.115 ;
        RECT 61.665 197.785 61.835 198.705 ;
        RECT 60.645 197.205 60.830 197.785 ;
        RECT 61.100 197.210 61.295 197.785 ;
        RECT 61.505 196.875 61.835 197.255 ;
        RECT 62.005 197.045 62.265 199.255 ;
        RECT 62.435 198.285 62.710 199.255 ;
        RECT 62.920 198.625 63.200 199.425 ;
        RECT 63.370 198.915 64.985 199.245 ;
        RECT 63.370 198.575 64.545 198.745 ;
        RECT 63.370 198.455 63.540 198.575 ;
        RECT 62.880 198.285 63.540 198.455 ;
        RECT 62.435 197.550 62.605 198.285 ;
        RECT 62.880 198.115 63.050 198.285 ;
        RECT 63.800 198.115 64.045 198.405 ;
        RECT 64.215 198.285 64.545 198.575 ;
        RECT 64.805 198.115 64.975 198.675 ;
        RECT 65.225 198.285 65.485 199.425 ;
        RECT 65.660 198.285 65.980 199.425 ;
        RECT 66.160 198.115 66.355 199.165 ;
        RECT 66.535 198.575 66.865 199.255 ;
        RECT 67.065 198.625 67.320 199.425 ;
        RECT 66.535 198.295 66.885 198.575 ;
        RECT 62.775 197.785 63.050 198.115 ;
        RECT 63.220 197.785 64.045 198.115 ;
        RECT 64.260 197.785 64.975 198.115 ;
        RECT 65.145 197.865 65.480 198.115 ;
        RECT 65.720 198.065 65.980 198.115 ;
        RECT 65.715 197.895 65.980 198.065 ;
        RECT 65.720 197.785 65.980 197.895 ;
        RECT 66.160 197.785 66.545 198.115 ;
        RECT 66.715 197.915 66.885 198.295 ;
        RECT 67.075 198.085 67.320 198.445 ;
        RECT 67.495 198.335 68.705 199.425 ;
        RECT 62.880 197.615 63.050 197.785 ;
        RECT 64.725 197.695 64.975 197.785 ;
        RECT 66.715 197.745 67.235 197.915 ;
        RECT 62.435 197.205 62.710 197.550 ;
        RECT 62.880 197.445 64.545 197.615 ;
        RECT 62.900 196.875 63.275 197.275 ;
        RECT 63.445 197.095 63.615 197.445 ;
        RECT 63.785 196.875 64.115 197.275 ;
        RECT 64.285 197.045 64.545 197.445 ;
        RECT 64.725 197.275 65.055 197.695 ;
        RECT 65.225 196.875 65.485 197.695 ;
        RECT 65.660 197.405 66.875 197.575 ;
        RECT 65.660 197.055 65.950 197.405 ;
        RECT 66.145 196.875 66.475 197.235 ;
        RECT 66.645 197.100 66.875 197.405 ;
        RECT 67.065 197.180 67.235 197.745 ;
        RECT 67.495 197.625 68.015 198.165 ;
        RECT 68.185 197.795 68.705 198.335 ;
        RECT 68.885 198.455 69.215 199.240 ;
        RECT 68.885 198.285 69.565 198.455 ;
        RECT 69.745 198.285 70.075 199.425 ;
        RECT 70.345 198.755 70.515 199.255 ;
        RECT 70.685 198.925 71.015 199.425 ;
        RECT 70.345 198.585 71.010 198.755 ;
        RECT 68.875 197.865 69.225 198.115 ;
        RECT 69.395 197.685 69.565 198.285 ;
        RECT 69.735 197.865 70.085 198.115 ;
        RECT 70.260 197.765 70.610 198.415 ;
        RECT 67.495 196.875 68.705 197.625 ;
        RECT 68.895 196.875 69.135 197.685 ;
        RECT 69.305 197.045 69.635 197.685 ;
        RECT 69.805 196.875 70.075 197.685 ;
        RECT 70.780 197.595 71.010 198.585 ;
        RECT 70.345 197.425 71.010 197.595 ;
        RECT 70.345 197.135 70.515 197.425 ;
        RECT 70.685 196.875 71.015 197.255 ;
        RECT 71.185 197.135 71.370 199.255 ;
        RECT 71.610 198.965 71.875 199.425 ;
        RECT 72.045 198.830 72.295 199.255 ;
        RECT 72.505 198.980 73.610 199.150 ;
        RECT 71.990 198.700 72.295 198.830 ;
        RECT 71.540 197.505 71.820 198.455 ;
        RECT 71.990 197.595 72.160 198.700 ;
        RECT 72.330 197.915 72.570 198.510 ;
        RECT 72.740 198.445 73.270 198.810 ;
        RECT 72.740 197.745 72.910 198.445 ;
        RECT 73.440 198.365 73.610 198.980 ;
        RECT 73.780 198.625 73.950 199.425 ;
        RECT 74.120 198.925 74.370 199.255 ;
        RECT 74.595 198.955 75.480 199.125 ;
        RECT 73.440 198.275 73.950 198.365 ;
        RECT 71.990 197.465 72.215 197.595 ;
        RECT 72.385 197.525 72.910 197.745 ;
        RECT 73.080 198.105 73.950 198.275 ;
        RECT 71.625 196.875 71.875 197.335 ;
        RECT 72.045 197.325 72.215 197.465 ;
        RECT 73.080 197.325 73.250 198.105 ;
        RECT 73.780 198.035 73.950 198.105 ;
        RECT 73.460 197.855 73.660 197.885 ;
        RECT 74.120 197.855 74.290 198.925 ;
        RECT 74.460 198.035 74.650 198.755 ;
        RECT 73.460 197.555 74.290 197.855 ;
        RECT 74.820 197.825 75.140 198.785 ;
        RECT 72.045 197.155 72.380 197.325 ;
        RECT 72.575 197.155 73.250 197.325 ;
        RECT 73.570 196.875 73.940 197.375 ;
        RECT 74.120 197.325 74.290 197.555 ;
        RECT 74.675 197.495 75.140 197.825 ;
        RECT 75.310 198.115 75.480 198.955 ;
        RECT 75.660 198.925 75.975 199.425 ;
        RECT 76.205 198.695 76.545 199.255 ;
        RECT 75.650 198.320 76.545 198.695 ;
        RECT 76.715 198.415 76.885 199.425 ;
        RECT 76.355 198.115 76.545 198.320 ;
        RECT 77.055 198.365 77.385 199.210 ;
        RECT 77.685 198.420 77.940 199.225 ;
        RECT 78.110 198.590 78.370 199.425 ;
        RECT 78.540 198.420 78.800 199.225 ;
        RECT 78.970 198.590 79.225 199.425 ;
        RECT 77.055 198.285 77.445 198.365 ;
        RECT 77.230 198.235 77.445 198.285 ;
        RECT 77.685 198.250 79.285 198.420 ;
        RECT 79.455 198.335 81.125 199.425 ;
        RECT 75.310 197.785 76.185 198.115 ;
        RECT 76.355 197.785 77.105 198.115 ;
        RECT 75.310 197.325 75.480 197.785 ;
        RECT 76.355 197.615 76.555 197.785 ;
        RECT 77.275 197.655 77.445 198.235 ;
        RECT 77.615 197.855 78.835 198.080 ;
        RECT 79.005 197.685 79.285 198.250 ;
        RECT 77.220 197.615 77.445 197.655 ;
        RECT 74.120 197.155 74.525 197.325 ;
        RECT 74.695 197.155 75.480 197.325 ;
        RECT 75.755 196.875 75.965 197.405 ;
        RECT 76.225 197.090 76.555 197.615 ;
        RECT 77.065 197.530 77.445 197.615 ;
        RECT 76.725 196.875 76.895 197.485 ;
        RECT 77.065 197.095 77.395 197.530 ;
        RECT 78.555 197.515 79.285 197.685 ;
        RECT 79.455 197.645 80.205 198.165 ;
        RECT 80.375 197.815 81.125 198.335 ;
        RECT 81.755 198.260 82.045 199.425 ;
        RECT 82.215 198.335 83.885 199.425 ;
        RECT 82.215 197.645 82.965 198.165 ;
        RECT 83.135 197.815 83.885 198.335 ;
        RECT 78.090 196.875 78.385 197.400 ;
        RECT 78.555 197.070 78.780 197.515 ;
        RECT 78.950 196.875 79.280 197.345 ;
        RECT 79.455 196.875 81.125 197.645 ;
        RECT 81.755 196.875 82.045 197.600 ;
        RECT 82.215 196.875 83.885 197.645 ;
        RECT 84.065 197.055 84.325 199.245 ;
        RECT 84.495 198.695 84.835 199.425 ;
        RECT 85.015 198.515 85.285 199.245 ;
        RECT 84.515 198.295 85.285 198.515 ;
        RECT 85.465 198.535 85.695 199.245 ;
        RECT 85.865 198.715 86.195 199.425 ;
        RECT 86.365 198.535 86.625 199.245 ;
        RECT 85.465 198.295 86.625 198.535 ;
        RECT 86.815 198.335 88.485 199.425 ;
        RECT 84.515 197.625 84.805 198.295 ;
        RECT 84.985 197.805 85.450 198.115 ;
        RECT 85.630 197.805 86.155 198.115 ;
        RECT 84.515 197.425 85.745 197.625 ;
        RECT 84.585 196.875 85.255 197.245 ;
        RECT 85.435 197.055 85.745 197.425 ;
        RECT 85.925 197.165 86.155 197.805 ;
        RECT 86.335 197.785 86.635 198.115 ;
        RECT 86.815 197.645 87.565 198.165 ;
        RECT 87.735 197.815 88.485 198.335 ;
        RECT 89.115 198.285 89.375 199.425 ;
        RECT 89.545 198.275 89.875 199.255 ;
        RECT 90.045 198.285 90.325 199.425 ;
        RECT 90.505 198.285 90.835 199.425 ;
        RECT 91.365 198.455 91.695 199.240 ;
        RECT 91.015 198.285 91.695 198.455 ;
        RECT 91.935 198.285 92.145 199.425 ;
        RECT 89.135 197.865 89.470 198.115 ;
        RECT 89.640 197.725 89.810 198.275 ;
        RECT 89.980 197.845 90.315 198.115 ;
        RECT 90.495 197.865 90.845 198.115 ;
        RECT 89.635 197.675 89.810 197.725 ;
        RECT 91.015 197.685 91.185 198.285 ;
        RECT 92.315 198.275 92.645 199.255 ;
        RECT 92.815 198.285 93.045 199.425 ;
        RECT 93.275 198.535 93.535 199.245 ;
        RECT 93.705 198.715 94.035 199.425 ;
        RECT 94.205 198.535 94.435 199.245 ;
        RECT 93.275 198.295 94.435 198.535 ;
        RECT 94.615 198.515 94.885 199.245 ;
        RECT 95.065 198.695 95.405 199.425 ;
        RECT 94.615 198.295 95.385 198.515 ;
        RECT 91.355 197.865 91.705 198.115 ;
        RECT 86.335 196.875 86.625 197.605 ;
        RECT 86.815 196.875 88.485 197.645 ;
        RECT 89.115 197.045 89.810 197.675 ;
        RECT 90.015 196.875 90.325 197.675 ;
        RECT 90.505 196.875 90.775 197.685 ;
        RECT 90.945 197.045 91.275 197.685 ;
        RECT 91.445 196.875 91.685 197.685 ;
        RECT 91.935 196.875 92.145 197.695 ;
        RECT 92.315 197.675 92.565 198.275 ;
        RECT 92.735 197.865 93.065 198.115 ;
        RECT 93.265 197.785 93.565 198.115 ;
        RECT 93.745 197.805 94.270 198.115 ;
        RECT 94.450 197.805 94.915 198.115 ;
        RECT 92.315 197.045 92.645 197.675 ;
        RECT 92.815 196.875 93.045 197.695 ;
        RECT 93.275 196.875 93.565 197.605 ;
        RECT 93.745 197.165 93.975 197.805 ;
        RECT 95.095 197.625 95.385 198.295 ;
        RECT 94.155 197.425 95.385 197.625 ;
        RECT 94.155 197.055 94.465 197.425 ;
        RECT 94.645 196.875 95.315 197.245 ;
        RECT 95.575 197.055 95.835 199.245 ;
        RECT 96.015 198.575 96.355 199.215 ;
        RECT 96.525 198.965 96.770 199.425 ;
        RECT 96.945 198.795 97.195 199.255 ;
        RECT 97.385 199.045 98.055 199.425 ;
        RECT 98.255 198.795 98.505 199.255 ;
        RECT 96.945 198.625 98.505 198.795 ;
        RECT 96.015 197.460 96.185 198.575 ;
        RECT 99.265 198.455 99.435 199.255 ;
        RECT 96.495 198.285 99.435 198.455 ;
        RECT 99.730 198.635 100.265 199.255 ;
        RECT 96.495 198.115 96.665 198.285 ;
        RECT 96.355 197.785 96.665 198.115 ;
        RECT 96.835 197.785 97.170 198.115 ;
        RECT 96.495 197.615 96.665 197.785 ;
        RECT 96.015 197.045 96.325 197.460 ;
        RECT 96.495 197.445 97.190 197.615 ;
        RECT 97.440 197.540 97.635 198.115 ;
        RECT 97.895 197.785 98.240 198.115 ;
        RECT 98.550 197.785 99.025 198.115 ;
        RECT 99.280 197.785 99.465 198.115 ;
        RECT 97.895 197.555 98.085 197.785 ;
        RECT 99.730 197.615 100.045 198.635 ;
        RECT 100.435 198.625 100.765 199.425 ;
        RECT 101.250 198.455 101.640 198.630 ;
        RECT 100.215 198.285 101.640 198.455 ;
        RECT 102.015 198.585 102.270 199.255 ;
        RECT 102.440 198.665 102.770 199.425 ;
        RECT 102.940 198.825 103.190 199.255 ;
        RECT 103.360 199.005 103.715 199.425 ;
        RECT 103.905 199.085 105.075 199.255 ;
        RECT 103.905 199.045 104.235 199.085 ;
        RECT 104.345 198.825 104.575 198.915 ;
        RECT 102.940 198.585 104.575 198.825 ;
        RECT 104.745 198.585 105.075 199.085 ;
        RECT 100.215 197.785 100.385 198.285 ;
        RECT 96.520 196.875 96.850 197.255 ;
        RECT 97.020 197.215 97.190 197.445 ;
        RECT 98.255 197.445 99.435 197.615 ;
        RECT 98.255 197.215 98.425 197.445 ;
        RECT 97.020 197.045 98.425 197.215 ;
        RECT 98.695 196.875 99.025 197.275 ;
        RECT 99.265 197.045 99.435 197.445 ;
        RECT 99.730 197.045 100.345 197.615 ;
        RECT 100.635 197.555 100.900 198.115 ;
        RECT 101.070 197.385 101.240 198.285 ;
        RECT 101.410 197.555 101.765 198.115 ;
        RECT 102.015 197.455 102.185 198.585 ;
        RECT 105.245 198.415 105.415 199.255 ;
        RECT 102.355 198.245 105.415 198.415 ;
        RECT 105.715 198.285 105.945 199.425 ;
        RECT 106.115 198.275 106.445 199.255 ;
        RECT 106.615 198.285 106.825 199.425 ;
        RECT 102.355 197.695 102.525 198.245 ;
        RECT 102.755 197.865 103.120 198.065 ;
        RECT 103.290 197.865 103.620 198.065 ;
        RECT 102.355 197.525 103.155 197.695 ;
        RECT 102.015 197.385 102.200 197.455 ;
        RECT 100.515 196.875 100.730 197.385 ;
        RECT 100.960 197.055 101.240 197.385 ;
        RECT 101.420 196.875 101.660 197.385 ;
        RECT 102.015 197.375 102.225 197.385 ;
        RECT 102.015 197.045 102.270 197.375 ;
        RECT 102.485 196.875 102.815 197.355 ;
        RECT 102.985 197.295 103.155 197.525 ;
        RECT 103.335 197.465 103.620 197.865 ;
        RECT 103.890 197.865 104.365 198.065 ;
        RECT 104.535 197.865 104.980 198.065 ;
        RECT 105.150 197.865 105.500 198.075 ;
        RECT 105.695 197.865 106.025 198.115 ;
        RECT 103.890 197.465 104.170 197.865 ;
        RECT 104.350 197.525 105.415 197.695 ;
        RECT 104.350 197.295 104.520 197.525 ;
        RECT 102.985 197.045 104.520 197.295 ;
        RECT 104.745 196.875 105.075 197.355 ;
        RECT 105.245 197.045 105.415 197.525 ;
        RECT 105.715 196.875 105.945 197.695 ;
        RECT 106.195 197.675 106.445 198.275 ;
        RECT 107.515 198.260 107.805 199.425 ;
        RECT 107.985 198.455 108.315 199.240 ;
        RECT 107.985 198.285 108.665 198.455 ;
        RECT 108.845 198.285 109.175 199.425 ;
        RECT 110.280 198.285 110.615 199.255 ;
        RECT 110.785 198.285 110.955 199.425 ;
        RECT 111.125 199.085 113.155 199.255 ;
        RECT 107.975 197.865 108.325 198.115 ;
        RECT 106.115 197.045 106.445 197.675 ;
        RECT 106.615 196.875 106.825 197.695 ;
        RECT 108.495 197.685 108.665 198.285 ;
        RECT 108.835 197.865 109.185 198.115 ;
        RECT 107.515 196.875 107.805 197.600 ;
        RECT 107.995 196.875 108.235 197.685 ;
        RECT 108.405 197.045 108.735 197.685 ;
        RECT 108.905 196.875 109.175 197.685 ;
        RECT 110.280 197.615 110.450 198.285 ;
        RECT 111.125 198.115 111.295 199.085 ;
        RECT 110.620 197.785 110.875 198.115 ;
        RECT 111.100 197.785 111.295 198.115 ;
        RECT 111.465 198.745 112.590 198.915 ;
        RECT 110.705 197.615 110.875 197.785 ;
        RECT 111.465 197.615 111.635 198.745 ;
        RECT 110.280 197.045 110.535 197.615 ;
        RECT 110.705 197.445 111.635 197.615 ;
        RECT 111.805 198.405 112.815 198.575 ;
        RECT 111.805 197.605 111.975 198.405 ;
        RECT 112.180 197.725 112.455 198.205 ;
        RECT 112.175 197.555 112.455 197.725 ;
        RECT 111.460 197.410 111.635 197.445 ;
        RECT 110.705 196.875 111.035 197.275 ;
        RECT 111.460 197.045 111.990 197.410 ;
        RECT 112.180 197.045 112.455 197.555 ;
        RECT 112.625 197.045 112.815 198.405 ;
        RECT 112.985 198.420 113.155 199.085 ;
        RECT 113.325 198.665 113.495 199.425 ;
        RECT 113.730 198.665 114.245 199.075 ;
        RECT 112.985 198.230 113.735 198.420 ;
        RECT 113.905 197.855 114.245 198.665 ;
        RECT 113.015 197.685 114.245 197.855 ;
        RECT 114.415 198.285 114.800 199.255 ;
        RECT 114.970 198.965 115.295 199.425 ;
        RECT 115.815 198.795 116.095 199.255 ;
        RECT 114.970 198.575 116.095 198.795 ;
        RECT 112.995 196.875 113.505 197.410 ;
        RECT 113.725 197.080 113.970 197.685 ;
        RECT 114.415 197.615 114.695 198.285 ;
        RECT 114.970 198.115 115.420 198.575 ;
        RECT 116.285 198.405 116.685 199.255 ;
        RECT 117.085 198.965 117.355 199.425 ;
        RECT 117.525 198.795 117.810 199.255 ;
        RECT 114.865 197.785 115.420 198.115 ;
        RECT 115.590 197.845 116.685 198.405 ;
        RECT 114.970 197.675 115.420 197.785 ;
        RECT 114.415 197.045 114.800 197.615 ;
        RECT 114.970 197.505 116.095 197.675 ;
        RECT 114.970 196.875 115.295 197.335 ;
        RECT 115.815 197.045 116.095 197.505 ;
        RECT 116.285 197.045 116.685 197.845 ;
        RECT 116.855 198.575 117.810 198.795 ;
        RECT 116.855 197.675 117.065 198.575 ;
        RECT 117.235 197.845 117.925 198.405 ;
        RECT 118.095 198.335 121.605 199.425 ;
        RECT 116.855 197.505 117.810 197.675 ;
        RECT 117.085 196.875 117.355 197.335 ;
        RECT 117.525 197.045 117.810 197.505 ;
        RECT 118.095 197.645 119.745 198.165 ;
        RECT 119.915 197.815 121.605 198.335 ;
        RECT 122.235 198.575 122.495 199.255 ;
        RECT 122.665 198.645 122.915 199.425 ;
        RECT 123.165 198.875 123.415 199.255 ;
        RECT 123.585 199.045 123.940 199.425 ;
        RECT 124.945 199.035 125.280 199.255 ;
        RECT 124.545 198.875 124.775 198.915 ;
        RECT 123.165 198.675 124.775 198.875 ;
        RECT 123.165 198.665 124.000 198.675 ;
        RECT 124.590 198.585 124.775 198.675 ;
        RECT 118.095 196.875 121.605 197.645 ;
        RECT 122.235 197.385 122.405 198.575 ;
        RECT 124.105 198.475 124.435 198.505 ;
        RECT 122.635 198.415 124.435 198.475 ;
        RECT 125.025 198.415 125.280 199.035 ;
        RECT 125.455 198.990 130.800 199.425 ;
        RECT 122.575 198.305 125.280 198.415 ;
        RECT 122.575 198.270 122.775 198.305 ;
        RECT 122.575 197.695 122.745 198.270 ;
        RECT 124.105 198.245 125.280 198.305 ;
        RECT 122.975 197.830 123.385 198.135 ;
        RECT 123.555 197.865 123.885 198.075 ;
        RECT 122.575 197.575 122.845 197.695 ;
        RECT 122.575 197.530 123.420 197.575 ;
        RECT 122.665 197.405 123.420 197.530 ;
        RECT 123.675 197.465 123.885 197.865 ;
        RECT 124.130 197.865 124.605 198.075 ;
        RECT 124.795 197.865 125.285 198.065 ;
        RECT 124.130 197.465 124.350 197.865 ;
        RECT 122.235 197.375 122.465 197.385 ;
        RECT 122.235 197.045 122.495 197.375 ;
        RECT 123.250 197.255 123.420 197.405 ;
        RECT 122.665 196.875 122.995 197.235 ;
        RECT 123.250 197.045 124.550 197.255 ;
        RECT 124.825 196.875 125.280 197.640 ;
        RECT 127.040 197.420 127.380 198.250 ;
        RECT 128.860 197.740 129.210 198.990 ;
        RECT 130.975 198.335 132.645 199.425 ;
        RECT 130.975 197.645 131.725 198.165 ;
        RECT 131.895 197.815 132.645 198.335 ;
        RECT 133.275 198.260 133.565 199.425 ;
        RECT 133.735 198.990 139.080 199.425 ;
        RECT 139.255 198.990 144.600 199.425 ;
        RECT 125.455 196.875 130.800 197.420 ;
        RECT 130.975 196.875 132.645 197.645 ;
        RECT 133.275 196.875 133.565 197.600 ;
        RECT 135.320 197.420 135.660 198.250 ;
        RECT 137.140 197.740 137.490 198.990 ;
        RECT 140.840 197.420 141.180 198.250 ;
        RECT 142.660 197.740 143.010 198.990 ;
        RECT 145.695 198.335 146.905 199.425 ;
        RECT 145.695 197.795 146.215 198.335 ;
        RECT 146.385 197.625 146.905 198.165 ;
        RECT 133.735 196.875 139.080 197.420 ;
        RECT 139.255 196.875 144.600 197.420 ;
        RECT 145.695 196.875 146.905 197.625 ;
        RECT 17.270 196.705 146.990 196.875 ;
        RECT 17.355 195.955 18.565 196.705 ;
        RECT 19.245 196.050 19.575 196.485 ;
        RECT 19.745 196.095 19.915 196.705 ;
        RECT 19.195 195.965 19.575 196.050 ;
        RECT 20.085 195.965 20.415 196.490 ;
        RECT 20.675 196.175 20.885 196.705 ;
        RECT 21.160 196.255 21.945 196.425 ;
        RECT 22.115 196.255 22.520 196.425 ;
        RECT 17.355 195.415 17.875 195.955 ;
        RECT 19.195 195.925 19.420 195.965 ;
        RECT 18.045 195.245 18.565 195.785 ;
        RECT 17.355 194.155 18.565 195.245 ;
        RECT 19.195 195.345 19.365 195.925 ;
        RECT 20.085 195.795 20.285 195.965 ;
        RECT 21.160 195.795 21.330 196.255 ;
        RECT 19.535 195.465 20.285 195.795 ;
        RECT 20.455 195.465 21.330 195.795 ;
        RECT 19.195 195.295 19.410 195.345 ;
        RECT 19.195 195.215 19.585 195.295 ;
        RECT 19.255 194.370 19.585 195.215 ;
        RECT 20.095 195.260 20.285 195.465 ;
        RECT 19.755 194.155 19.925 195.165 ;
        RECT 20.095 194.885 20.990 195.260 ;
        RECT 20.095 194.325 20.435 194.885 ;
        RECT 20.665 194.155 20.980 194.655 ;
        RECT 21.160 194.625 21.330 195.465 ;
        RECT 21.500 195.755 21.965 196.085 ;
        RECT 22.350 196.025 22.520 196.255 ;
        RECT 22.700 196.205 23.070 196.705 ;
        RECT 23.390 196.255 24.065 196.425 ;
        RECT 24.260 196.255 24.595 196.425 ;
        RECT 21.500 194.795 21.820 195.755 ;
        RECT 22.350 195.725 23.180 196.025 ;
        RECT 21.990 194.825 22.180 195.545 ;
        RECT 22.350 194.655 22.520 195.725 ;
        RECT 22.980 195.695 23.180 195.725 ;
        RECT 22.690 195.475 22.860 195.545 ;
        RECT 23.390 195.475 23.560 196.255 ;
        RECT 24.425 196.115 24.595 196.255 ;
        RECT 24.765 196.245 25.015 196.705 ;
        RECT 22.690 195.305 23.560 195.475 ;
        RECT 23.730 195.835 24.255 196.055 ;
        RECT 24.425 195.985 24.650 196.115 ;
        RECT 22.690 195.215 23.200 195.305 ;
        RECT 21.160 194.455 22.045 194.625 ;
        RECT 22.270 194.325 22.520 194.655 ;
        RECT 22.690 194.155 22.860 194.955 ;
        RECT 23.030 194.600 23.200 195.215 ;
        RECT 23.730 195.135 23.900 195.835 ;
        RECT 23.370 194.770 23.900 195.135 ;
        RECT 24.070 195.070 24.310 195.665 ;
        RECT 24.480 194.880 24.650 195.985 ;
        RECT 24.820 195.125 25.100 196.075 ;
        RECT 24.345 194.750 24.650 194.880 ;
        RECT 23.030 194.430 24.135 194.600 ;
        RECT 24.345 194.325 24.595 194.750 ;
        RECT 24.765 194.155 25.030 194.615 ;
        RECT 25.270 194.325 25.455 196.445 ;
        RECT 25.625 196.325 25.955 196.705 ;
        RECT 26.125 196.155 26.295 196.445 ;
        RECT 25.630 195.985 26.295 196.155 ;
        RECT 26.555 195.985 26.895 196.495 ;
        RECT 25.630 194.995 25.860 195.985 ;
        RECT 26.030 195.165 26.380 195.815 ;
        RECT 25.630 194.825 26.295 194.995 ;
        RECT 25.625 194.155 25.955 194.655 ;
        RECT 26.125 194.325 26.295 194.825 ;
        RECT 26.555 194.585 26.815 195.985 ;
        RECT 27.065 195.905 27.335 196.705 ;
        RECT 26.990 195.465 27.320 195.715 ;
        RECT 27.515 195.465 27.795 196.435 ;
        RECT 27.975 195.465 28.275 196.435 ;
        RECT 28.455 195.465 28.805 196.430 ;
        RECT 29.025 196.205 29.520 196.535 ;
        RECT 27.005 195.295 27.320 195.465 ;
        RECT 29.025 195.295 29.195 196.205 ;
        RECT 27.005 195.125 29.195 195.295 ;
        RECT 26.555 194.325 26.895 194.585 ;
        RECT 27.065 194.155 27.395 194.955 ;
        RECT 27.860 194.325 28.110 195.125 ;
        RECT 28.295 194.155 28.625 194.875 ;
        RECT 28.845 194.325 29.095 195.125 ;
        RECT 29.365 194.715 29.605 196.025 ;
        RECT 29.785 195.980 30.115 196.490 ;
        RECT 30.285 196.305 30.615 196.705 ;
        RECT 31.665 196.135 31.995 196.475 ;
        RECT 32.165 196.305 32.495 196.705 ;
        RECT 33.470 196.135 33.725 196.485 ;
        RECT 33.895 196.305 34.225 196.705 ;
        RECT 34.395 196.135 34.565 196.485 ;
        RECT 34.735 196.305 35.115 196.705 ;
        RECT 29.785 195.215 29.975 195.980 ;
        RECT 30.285 195.965 32.650 196.135 ;
        RECT 33.470 195.965 35.135 196.135 ;
        RECT 35.305 196.030 35.580 196.375 ;
        RECT 30.285 195.795 30.455 195.965 ;
        RECT 30.145 195.465 30.455 195.795 ;
        RECT 30.625 195.465 30.930 195.795 ;
        RECT 29.265 194.155 29.600 194.535 ;
        RECT 29.785 194.365 30.115 195.215 ;
        RECT 30.285 194.155 30.535 195.295 ;
        RECT 30.715 195.135 30.930 195.465 ;
        RECT 31.105 195.135 31.390 195.795 ;
        RECT 31.585 195.135 31.850 195.795 ;
        RECT 32.065 195.135 32.310 195.795 ;
        RECT 32.480 194.965 32.650 195.965 ;
        RECT 34.965 195.795 35.135 195.965 ;
        RECT 33.455 195.465 33.800 195.795 ;
        RECT 33.970 195.465 34.795 195.795 ;
        RECT 34.965 195.465 35.240 195.795 ;
        RECT 30.725 194.795 32.015 194.965 ;
        RECT 30.725 194.375 30.975 194.795 ;
        RECT 31.205 194.155 31.535 194.625 ;
        RECT 31.765 194.375 32.015 194.795 ;
        RECT 32.195 194.795 32.650 194.965 ;
        RECT 33.475 195.005 33.800 195.295 ;
        RECT 33.970 195.175 34.165 195.465 ;
        RECT 34.965 195.295 35.135 195.465 ;
        RECT 35.410 195.295 35.580 196.030 ;
        RECT 35.755 196.095 36.095 196.510 ;
        RECT 36.265 196.265 36.435 196.705 ;
        RECT 36.605 196.315 37.855 196.495 ;
        RECT 36.605 196.095 36.935 196.315 ;
        RECT 38.125 196.245 38.295 196.705 ;
        RECT 35.755 195.925 36.935 196.095 ;
        RECT 37.105 196.075 37.470 196.145 ;
        RECT 37.105 195.895 38.355 196.075 ;
        RECT 35.755 195.515 36.220 195.715 ;
        RECT 36.395 195.465 36.725 195.715 ;
        RECT 36.895 195.685 37.360 195.715 ;
        RECT 36.895 195.515 37.365 195.685 ;
        RECT 36.895 195.465 37.360 195.515 ;
        RECT 37.555 195.465 37.910 195.715 ;
        RECT 36.395 195.345 36.575 195.465 ;
        RECT 34.475 195.125 35.135 195.295 ;
        RECT 34.475 195.005 34.645 195.125 ;
        RECT 33.475 194.835 34.645 195.005 ;
        RECT 32.195 194.365 32.525 194.795 ;
        RECT 33.455 194.375 34.645 194.665 ;
        RECT 34.815 194.155 35.095 194.955 ;
        RECT 35.305 194.325 35.580 195.295 ;
        RECT 35.755 194.155 36.075 195.335 ;
        RECT 36.245 195.175 36.575 195.345 ;
        RECT 38.080 195.295 38.355 195.895 ;
        RECT 36.245 194.385 36.445 195.175 ;
        RECT 36.745 195.085 38.355 195.295 ;
        RECT 36.745 194.985 37.155 195.085 ;
        RECT 36.770 194.325 37.155 194.985 ;
        RECT 37.550 194.155 38.335 194.915 ;
        RECT 38.525 194.325 38.805 196.425 ;
        RECT 38.980 195.940 39.435 196.705 ;
        RECT 39.710 196.325 41.010 196.535 ;
        RECT 41.265 196.345 41.595 196.705 ;
        RECT 40.840 196.175 41.010 196.325 ;
        RECT 41.765 196.205 42.025 196.535 ;
        RECT 39.910 195.715 40.130 196.115 ;
        RECT 38.975 195.515 39.465 195.715 ;
        RECT 39.655 195.505 40.130 195.715 ;
        RECT 40.375 195.715 40.585 196.115 ;
        RECT 40.840 196.050 41.595 196.175 ;
        RECT 40.840 196.005 41.685 196.050 ;
        RECT 41.415 195.885 41.685 196.005 ;
        RECT 40.375 195.505 40.705 195.715 ;
        RECT 40.875 195.445 41.285 195.750 ;
        RECT 38.980 195.275 40.155 195.335 ;
        RECT 41.515 195.310 41.685 195.885 ;
        RECT 41.485 195.275 41.685 195.310 ;
        RECT 38.980 195.165 41.685 195.275 ;
        RECT 38.980 194.545 39.235 195.165 ;
        RECT 39.825 195.105 41.625 195.165 ;
        RECT 39.825 195.075 40.155 195.105 ;
        RECT 41.855 195.005 42.025 196.205 ;
        RECT 43.115 195.980 43.405 196.705 ;
        RECT 43.580 196.055 43.850 196.265 ;
        RECT 44.070 196.245 44.400 196.705 ;
        RECT 44.910 196.245 45.660 196.535 ;
        RECT 45.880 196.305 46.215 196.705 ;
        RECT 43.580 195.885 44.915 196.055 ;
        RECT 44.745 195.715 44.915 195.885 ;
        RECT 43.580 195.475 43.930 195.715 ;
        RECT 44.100 195.475 44.575 195.715 ;
        RECT 44.745 195.465 45.120 195.715 ;
        RECT 39.485 194.905 39.670 194.995 ;
        RECT 40.260 194.905 41.095 194.915 ;
        RECT 39.485 194.705 41.095 194.905 ;
        RECT 39.485 194.665 39.715 194.705 ;
        RECT 38.980 194.325 39.315 194.545 ;
        RECT 40.320 194.155 40.675 194.535 ;
        RECT 40.845 194.325 41.095 194.705 ;
        RECT 41.345 194.155 41.595 194.935 ;
        RECT 41.765 194.325 42.025 195.005 ;
        RECT 43.115 194.155 43.405 195.320 ;
        RECT 44.745 195.295 44.915 195.465 ;
        RECT 43.580 195.125 44.915 195.295 ;
        RECT 43.580 194.965 43.860 195.125 ;
        RECT 45.290 194.955 45.660 196.245 ;
        RECT 46.385 196.135 46.590 196.535 ;
        RECT 46.800 196.225 47.075 196.705 ;
        RECT 47.285 196.205 47.545 196.535 ;
        RECT 44.070 194.155 44.320 194.955 ;
        RECT 44.490 194.785 45.660 194.955 ;
        RECT 45.905 195.965 46.590 196.135 ;
        RECT 45.905 194.935 46.245 195.965 ;
        RECT 46.415 195.295 46.665 195.795 ;
        RECT 46.845 195.465 47.205 196.045 ;
        RECT 47.375 195.295 47.545 196.205 ;
        RECT 47.715 195.935 50.305 196.705 ;
        RECT 47.715 195.415 48.925 195.935 ;
        RECT 50.935 195.905 51.245 196.705 ;
        RECT 51.450 195.905 52.145 196.535 ;
        RECT 52.330 196.135 52.585 196.485 ;
        RECT 52.755 196.305 53.085 196.705 ;
        RECT 53.255 196.135 53.425 196.485 ;
        RECT 53.595 196.305 53.975 196.705 ;
        RECT 52.330 195.965 53.995 196.135 ;
        RECT 54.165 196.030 54.440 196.375 ;
        RECT 46.415 195.125 47.545 195.295 ;
        RECT 49.095 195.245 50.305 195.765 ;
        RECT 50.945 195.465 51.280 195.735 ;
        RECT 51.450 195.305 51.620 195.905 ;
        RECT 53.825 195.795 53.995 195.965 ;
        RECT 51.790 195.465 52.125 195.715 ;
        RECT 52.315 195.465 52.660 195.795 ;
        RECT 52.830 195.465 53.655 195.795 ;
        RECT 53.825 195.465 54.100 195.795 ;
        RECT 44.490 194.325 44.820 194.785 ;
        RECT 45.905 194.760 46.570 194.935 ;
        RECT 44.990 194.155 45.205 194.615 ;
        RECT 45.880 194.155 46.215 194.580 ;
        RECT 46.385 194.355 46.570 194.760 ;
        RECT 46.775 194.155 47.105 194.935 ;
        RECT 47.275 194.355 47.545 195.125 ;
        RECT 47.715 194.155 50.305 195.245 ;
        RECT 50.935 194.155 51.215 195.295 ;
        RECT 51.385 194.325 51.715 195.305 ;
        RECT 51.885 194.155 52.145 195.295 ;
        RECT 52.335 195.005 52.660 195.295 ;
        RECT 52.830 195.175 53.025 195.465 ;
        RECT 53.825 195.295 53.995 195.465 ;
        RECT 54.270 195.295 54.440 196.030 ;
        RECT 53.335 195.125 53.995 195.295 ;
        RECT 53.335 195.005 53.505 195.125 ;
        RECT 52.335 194.835 53.505 195.005 ;
        RECT 52.315 194.375 53.505 194.665 ;
        RECT 53.675 194.155 53.955 194.955 ;
        RECT 54.165 194.325 54.440 195.295 ;
        RECT 54.615 194.325 54.895 196.425 ;
        RECT 55.125 196.245 55.295 196.705 ;
        RECT 55.565 196.315 56.815 196.495 ;
        RECT 55.950 196.075 56.315 196.145 ;
        RECT 55.065 195.895 56.315 196.075 ;
        RECT 56.485 196.095 56.815 196.315 ;
        RECT 56.985 196.265 57.155 196.705 ;
        RECT 57.325 196.095 57.665 196.510 ;
        RECT 56.485 195.925 57.665 196.095 ;
        RECT 58.040 195.925 58.540 196.535 ;
        RECT 55.065 195.295 55.340 195.895 ;
        RECT 55.510 195.465 55.865 195.715 ;
        RECT 56.060 195.685 56.525 195.715 ;
        RECT 56.055 195.515 56.525 195.685 ;
        RECT 56.060 195.465 56.525 195.515 ;
        RECT 56.695 195.465 57.025 195.715 ;
        RECT 57.200 195.515 57.665 195.715 ;
        RECT 57.835 195.465 58.185 195.715 ;
        RECT 56.845 195.345 57.025 195.465 ;
        RECT 55.065 195.085 56.675 195.295 ;
        RECT 56.845 195.175 57.175 195.345 ;
        RECT 56.265 194.985 56.675 195.085 ;
        RECT 55.085 194.155 55.870 194.915 ;
        RECT 56.265 194.325 56.650 194.985 ;
        RECT 56.975 194.385 57.175 195.175 ;
        RECT 57.345 194.155 57.665 195.335 ;
        RECT 58.370 195.295 58.540 195.925 ;
        RECT 59.170 196.055 59.500 196.535 ;
        RECT 59.670 196.245 59.895 196.705 ;
        RECT 60.065 196.055 60.395 196.535 ;
        RECT 59.170 195.885 60.395 196.055 ;
        RECT 60.585 195.905 60.835 196.705 ;
        RECT 61.005 195.905 61.345 196.535 ;
        RECT 61.535 195.975 61.825 196.705 ;
        RECT 58.710 195.515 59.040 195.715 ;
        RECT 59.210 195.515 59.540 195.715 ;
        RECT 59.710 195.515 60.130 195.715 ;
        RECT 60.305 195.545 61.000 195.715 ;
        RECT 60.305 195.295 60.475 195.545 ;
        RECT 61.170 195.295 61.345 195.905 ;
        RECT 61.525 195.465 61.825 195.795 ;
        RECT 62.005 195.775 62.235 196.415 ;
        RECT 62.415 196.155 62.725 196.525 ;
        RECT 62.905 196.335 63.575 196.705 ;
        RECT 62.415 195.955 63.645 196.155 ;
        RECT 62.005 195.465 62.530 195.775 ;
        RECT 62.710 195.465 63.175 195.775 ;
        RECT 58.040 195.125 60.475 195.295 ;
        RECT 58.040 194.325 58.370 195.125 ;
        RECT 58.540 194.155 58.870 194.955 ;
        RECT 59.170 194.325 59.500 195.125 ;
        RECT 60.145 194.155 60.395 194.955 ;
        RECT 60.665 194.155 60.835 195.295 ;
        RECT 61.005 194.325 61.345 195.295 ;
        RECT 63.355 195.285 63.645 195.955 ;
        RECT 61.535 195.045 62.695 195.285 ;
        RECT 61.535 194.335 61.795 195.045 ;
        RECT 61.965 194.155 62.295 194.865 ;
        RECT 62.465 194.335 62.695 195.045 ;
        RECT 62.875 195.065 63.645 195.285 ;
        RECT 62.875 194.335 63.145 195.065 ;
        RECT 63.325 194.155 63.665 194.885 ;
        RECT 63.835 194.335 64.095 196.525 ;
        RECT 64.275 195.935 67.785 196.705 ;
        RECT 68.875 195.980 69.165 196.705 ;
        RECT 69.335 195.935 71.005 196.705 ;
        RECT 71.180 196.135 71.435 196.405 ;
        RECT 71.605 196.305 71.935 196.705 ;
        RECT 72.105 196.135 72.275 196.405 ;
        RECT 72.445 196.305 72.775 196.705 ;
        RECT 71.180 195.965 72.405 196.135 ;
        RECT 64.275 195.415 65.925 195.935 ;
        RECT 66.095 195.245 67.785 195.765 ;
        RECT 69.335 195.415 70.085 195.935 ;
        RECT 64.275 194.155 67.785 195.245 ;
        RECT 68.875 194.155 69.165 195.320 ;
        RECT 70.255 195.245 71.005 195.765 ;
        RECT 71.180 195.465 71.515 195.795 ;
        RECT 71.685 195.465 72.065 195.795 ;
        RECT 69.335 194.155 71.005 195.245 ;
        RECT 71.180 194.510 71.515 195.295 ;
        RECT 71.685 194.785 71.920 195.465 ;
        RECT 72.235 195.295 72.405 195.965 ;
        RECT 72.090 195.125 72.405 195.295 ;
        RECT 72.575 195.125 72.845 196.135 ;
        RECT 73.065 196.050 73.395 196.485 ;
        RECT 73.565 196.095 73.735 196.705 ;
        RECT 73.015 195.965 73.395 196.050 ;
        RECT 73.905 195.965 74.235 196.490 ;
        RECT 74.495 196.175 74.705 196.705 ;
        RECT 74.980 196.255 75.765 196.425 ;
        RECT 75.935 196.255 76.340 196.425 ;
        RECT 73.015 195.925 73.240 195.965 ;
        RECT 73.015 195.345 73.185 195.925 ;
        RECT 73.905 195.795 74.105 195.965 ;
        RECT 74.980 195.795 75.150 196.255 ;
        RECT 73.355 195.465 74.105 195.795 ;
        RECT 74.275 195.465 75.150 195.795 ;
        RECT 73.015 195.295 73.230 195.345 ;
        RECT 73.015 195.215 73.405 195.295 ;
        RECT 72.090 194.510 72.260 195.125 ;
        RECT 71.180 194.340 72.260 194.510 ;
        RECT 72.525 194.155 72.840 194.955 ;
        RECT 73.075 194.370 73.405 195.215 ;
        RECT 73.915 195.260 74.105 195.465 ;
        RECT 73.575 194.155 73.745 195.165 ;
        RECT 73.915 194.885 74.810 195.260 ;
        RECT 73.915 194.325 74.255 194.885 ;
        RECT 74.485 194.155 74.800 194.655 ;
        RECT 74.980 194.625 75.150 195.465 ;
        RECT 75.320 195.755 75.785 196.085 ;
        RECT 76.170 196.025 76.340 196.255 ;
        RECT 76.520 196.205 76.890 196.705 ;
        RECT 77.210 196.255 77.885 196.425 ;
        RECT 78.080 196.255 78.415 196.425 ;
        RECT 75.320 194.795 75.640 195.755 ;
        RECT 76.170 195.725 77.000 196.025 ;
        RECT 75.810 194.825 76.000 195.545 ;
        RECT 76.170 194.655 76.340 195.725 ;
        RECT 76.800 195.695 77.000 195.725 ;
        RECT 76.510 195.475 76.680 195.545 ;
        RECT 77.210 195.475 77.380 196.255 ;
        RECT 78.245 196.115 78.415 196.255 ;
        RECT 78.585 196.245 78.835 196.705 ;
        RECT 76.510 195.305 77.380 195.475 ;
        RECT 77.550 195.835 78.075 196.055 ;
        RECT 78.245 195.985 78.470 196.115 ;
        RECT 76.510 195.215 77.020 195.305 ;
        RECT 74.980 194.455 75.865 194.625 ;
        RECT 76.090 194.325 76.340 194.655 ;
        RECT 76.510 194.155 76.680 194.955 ;
        RECT 76.850 194.600 77.020 195.215 ;
        RECT 77.550 195.135 77.720 195.835 ;
        RECT 77.190 194.770 77.720 195.135 ;
        RECT 77.890 195.070 78.130 195.665 ;
        RECT 78.300 194.880 78.470 195.985 ;
        RECT 78.640 195.125 78.920 196.075 ;
        RECT 78.165 194.750 78.470 194.880 ;
        RECT 76.850 194.430 77.955 194.600 ;
        RECT 78.165 194.325 78.415 194.750 ;
        RECT 78.585 194.155 78.850 194.615 ;
        RECT 79.090 194.325 79.275 196.445 ;
        RECT 79.445 196.325 79.775 196.705 ;
        RECT 79.945 196.155 80.115 196.445 ;
        RECT 79.450 195.985 80.115 196.155 ;
        RECT 80.925 196.155 81.095 196.445 ;
        RECT 81.265 196.325 81.595 196.705 ;
        RECT 80.925 195.985 81.590 196.155 ;
        RECT 79.450 194.995 79.680 195.985 ;
        RECT 79.850 195.165 80.200 195.815 ;
        RECT 80.840 195.165 81.190 195.815 ;
        RECT 81.360 194.995 81.590 195.985 ;
        RECT 79.450 194.825 80.115 194.995 ;
        RECT 79.445 194.155 79.775 194.655 ;
        RECT 79.945 194.325 80.115 194.825 ;
        RECT 80.925 194.825 81.590 194.995 ;
        RECT 80.925 194.325 81.095 194.825 ;
        RECT 81.265 194.155 81.595 194.655 ;
        RECT 81.765 194.325 81.950 196.445 ;
        RECT 82.205 196.245 82.455 196.705 ;
        RECT 82.625 196.255 82.960 196.425 ;
        RECT 83.155 196.255 83.830 196.425 ;
        RECT 82.625 196.115 82.795 196.255 ;
        RECT 82.120 195.125 82.400 196.075 ;
        RECT 82.570 195.985 82.795 196.115 ;
        RECT 82.570 194.880 82.740 195.985 ;
        RECT 82.965 195.835 83.490 196.055 ;
        RECT 82.910 195.070 83.150 195.665 ;
        RECT 83.320 195.135 83.490 195.835 ;
        RECT 83.660 195.475 83.830 196.255 ;
        RECT 84.150 196.205 84.520 196.705 ;
        RECT 84.700 196.255 85.105 196.425 ;
        RECT 85.275 196.255 86.060 196.425 ;
        RECT 84.700 196.025 84.870 196.255 ;
        RECT 84.040 195.725 84.870 196.025 ;
        RECT 85.255 195.755 85.720 196.085 ;
        RECT 84.040 195.695 84.240 195.725 ;
        RECT 84.360 195.475 84.530 195.545 ;
        RECT 83.660 195.305 84.530 195.475 ;
        RECT 84.020 195.215 84.530 195.305 ;
        RECT 82.570 194.750 82.875 194.880 ;
        RECT 83.320 194.770 83.850 195.135 ;
        RECT 82.190 194.155 82.455 194.615 ;
        RECT 82.625 194.325 82.875 194.750 ;
        RECT 84.020 194.600 84.190 195.215 ;
        RECT 83.085 194.430 84.190 194.600 ;
        RECT 84.360 194.155 84.530 194.955 ;
        RECT 84.700 194.655 84.870 195.725 ;
        RECT 85.040 194.825 85.230 195.545 ;
        RECT 85.400 194.795 85.720 195.755 ;
        RECT 85.890 195.795 86.060 196.255 ;
        RECT 86.335 196.175 86.545 196.705 ;
        RECT 86.805 195.965 87.135 196.490 ;
        RECT 87.305 196.095 87.475 196.705 ;
        RECT 87.645 196.050 87.975 196.485 ;
        RECT 88.195 196.160 93.540 196.705 ;
        RECT 87.645 195.965 88.025 196.050 ;
        RECT 86.935 195.795 87.135 195.965 ;
        RECT 87.800 195.925 88.025 195.965 ;
        RECT 85.890 195.465 86.765 195.795 ;
        RECT 86.935 195.465 87.685 195.795 ;
        RECT 84.700 194.325 84.950 194.655 ;
        RECT 85.890 194.625 86.060 195.465 ;
        RECT 86.935 195.260 87.125 195.465 ;
        RECT 87.855 195.345 88.025 195.925 ;
        RECT 87.810 195.295 88.025 195.345 ;
        RECT 89.780 195.330 90.120 196.160 ;
        RECT 94.635 195.980 94.925 196.705 ;
        RECT 95.095 195.935 97.685 196.705 ;
        RECT 97.860 195.940 98.315 196.705 ;
        RECT 98.590 196.325 99.890 196.535 ;
        RECT 100.145 196.345 100.475 196.705 ;
        RECT 99.720 196.175 99.890 196.325 ;
        RECT 100.645 196.205 100.905 196.535 ;
        RECT 101.865 196.305 102.195 196.705 ;
        RECT 100.675 196.195 100.905 196.205 ;
        RECT 86.230 194.885 87.125 195.260 ;
        RECT 87.635 195.215 88.025 195.295 ;
        RECT 85.175 194.455 86.060 194.625 ;
        RECT 86.240 194.155 86.555 194.655 ;
        RECT 86.785 194.325 87.125 194.885 ;
        RECT 87.295 194.155 87.465 195.165 ;
        RECT 87.635 194.370 87.965 195.215 ;
        RECT 91.600 194.590 91.950 195.840 ;
        RECT 95.095 195.415 96.305 195.935 ;
        RECT 88.195 194.155 93.540 194.590 ;
        RECT 94.635 194.155 94.925 195.320 ;
        RECT 96.475 195.245 97.685 195.765 ;
        RECT 98.790 195.715 99.010 196.115 ;
        RECT 97.855 195.515 98.345 195.715 ;
        RECT 98.535 195.505 99.010 195.715 ;
        RECT 99.255 195.715 99.465 196.115 ;
        RECT 99.720 196.050 100.475 196.175 ;
        RECT 99.720 196.005 100.565 196.050 ;
        RECT 100.295 195.885 100.565 196.005 ;
        RECT 99.255 195.505 99.585 195.715 ;
        RECT 99.755 195.445 100.165 195.750 ;
        RECT 95.095 194.155 97.685 195.245 ;
        RECT 97.860 195.275 99.035 195.335 ;
        RECT 100.395 195.310 100.565 195.885 ;
        RECT 100.365 195.275 100.565 195.310 ;
        RECT 97.860 195.165 100.565 195.275 ;
        RECT 97.860 194.545 98.115 195.165 ;
        RECT 98.705 195.105 100.505 195.165 ;
        RECT 98.705 195.075 99.035 195.105 ;
        RECT 100.735 195.005 100.905 196.195 ;
        RECT 102.365 196.135 102.695 196.475 ;
        RECT 103.745 196.305 104.075 196.705 ;
        RECT 98.365 194.905 98.550 194.995 ;
        RECT 99.140 194.905 99.975 194.915 ;
        RECT 98.365 194.705 99.975 194.905 ;
        RECT 98.365 194.665 98.595 194.705 ;
        RECT 97.860 194.325 98.195 194.545 ;
        RECT 99.200 194.155 99.555 194.535 ;
        RECT 99.725 194.325 99.975 194.705 ;
        RECT 100.225 194.155 100.475 194.935 ;
        RECT 100.645 194.325 100.905 195.005 ;
        RECT 101.710 195.965 104.075 196.135 ;
        RECT 104.245 195.980 104.575 196.490 ;
        RECT 101.710 194.965 101.880 195.965 ;
        RECT 103.905 195.795 104.075 195.965 ;
        RECT 102.050 195.135 102.295 195.795 ;
        RECT 102.510 195.135 102.775 195.795 ;
        RECT 102.970 195.135 103.255 195.795 ;
        RECT 103.430 195.465 103.735 195.795 ;
        RECT 103.905 195.465 104.215 195.795 ;
        RECT 103.430 195.135 103.645 195.465 ;
        RECT 101.710 194.795 102.165 194.965 ;
        RECT 101.835 194.365 102.165 194.795 ;
        RECT 102.345 194.795 103.635 194.965 ;
        RECT 102.345 194.375 102.595 194.795 ;
        RECT 102.825 194.155 103.155 194.625 ;
        RECT 103.385 194.375 103.635 194.795 ;
        RECT 103.825 194.155 104.075 195.295 ;
        RECT 104.385 195.215 104.575 195.980 ;
        RECT 104.795 195.885 105.025 196.705 ;
        RECT 105.195 195.905 105.525 196.535 ;
        RECT 104.775 195.465 105.105 195.715 ;
        RECT 105.275 195.305 105.525 195.905 ;
        RECT 105.695 195.885 105.905 196.705 ;
        RECT 106.135 195.955 107.345 196.705 ;
        RECT 107.605 196.155 107.775 196.445 ;
        RECT 107.945 196.325 108.275 196.705 ;
        RECT 107.605 195.985 108.270 196.155 ;
        RECT 106.135 195.415 106.655 195.955 ;
        RECT 104.245 194.365 104.575 195.215 ;
        RECT 104.795 194.155 105.025 195.295 ;
        RECT 105.195 194.325 105.525 195.305 ;
        RECT 105.695 194.155 105.905 195.295 ;
        RECT 106.825 195.245 107.345 195.785 ;
        RECT 106.135 194.155 107.345 195.245 ;
        RECT 107.520 195.165 107.870 195.815 ;
        RECT 108.040 194.995 108.270 195.985 ;
        RECT 107.605 194.825 108.270 194.995 ;
        RECT 107.605 194.325 107.775 194.825 ;
        RECT 107.945 194.155 108.275 194.655 ;
        RECT 108.445 194.325 108.630 196.445 ;
        RECT 108.885 196.245 109.135 196.705 ;
        RECT 109.305 196.255 109.640 196.425 ;
        RECT 109.835 196.255 110.510 196.425 ;
        RECT 109.305 196.115 109.475 196.255 ;
        RECT 108.800 195.125 109.080 196.075 ;
        RECT 109.250 195.985 109.475 196.115 ;
        RECT 109.250 194.880 109.420 195.985 ;
        RECT 109.645 195.835 110.170 196.055 ;
        RECT 109.590 195.070 109.830 195.665 ;
        RECT 110.000 195.135 110.170 195.835 ;
        RECT 110.340 195.475 110.510 196.255 ;
        RECT 110.830 196.205 111.200 196.705 ;
        RECT 111.380 196.255 111.785 196.425 ;
        RECT 111.955 196.255 112.740 196.425 ;
        RECT 111.380 196.025 111.550 196.255 ;
        RECT 110.720 195.725 111.550 196.025 ;
        RECT 111.935 195.755 112.400 196.085 ;
        RECT 110.720 195.695 110.920 195.725 ;
        RECT 111.040 195.475 111.210 195.545 ;
        RECT 110.340 195.305 111.210 195.475 ;
        RECT 110.700 195.215 111.210 195.305 ;
        RECT 109.250 194.750 109.555 194.880 ;
        RECT 110.000 194.770 110.530 195.135 ;
        RECT 108.870 194.155 109.135 194.615 ;
        RECT 109.305 194.325 109.555 194.750 ;
        RECT 110.700 194.600 110.870 195.215 ;
        RECT 109.765 194.430 110.870 194.600 ;
        RECT 111.040 194.155 111.210 194.955 ;
        RECT 111.380 194.655 111.550 195.725 ;
        RECT 111.720 194.825 111.910 195.545 ;
        RECT 112.080 194.795 112.400 195.755 ;
        RECT 112.570 195.795 112.740 196.255 ;
        RECT 113.015 196.175 113.225 196.705 ;
        RECT 113.485 195.965 113.815 196.490 ;
        RECT 113.985 196.095 114.155 196.705 ;
        RECT 114.325 196.050 114.655 196.485 ;
        RECT 114.875 196.160 120.220 196.705 ;
        RECT 114.325 195.965 114.705 196.050 ;
        RECT 113.615 195.795 113.815 195.965 ;
        RECT 114.480 195.925 114.705 195.965 ;
        RECT 112.570 195.465 113.445 195.795 ;
        RECT 113.615 195.465 114.365 195.795 ;
        RECT 111.380 194.325 111.630 194.655 ;
        RECT 112.570 194.625 112.740 195.465 ;
        RECT 113.615 195.260 113.805 195.465 ;
        RECT 114.535 195.345 114.705 195.925 ;
        RECT 114.490 195.295 114.705 195.345 ;
        RECT 116.460 195.330 116.800 196.160 ;
        RECT 120.395 195.980 120.685 196.705 ;
        RECT 120.860 195.965 121.115 196.535 ;
        RECT 121.285 196.305 121.615 196.705 ;
        RECT 122.040 196.170 122.570 196.535 ;
        RECT 122.040 196.135 122.215 196.170 ;
        RECT 121.285 195.965 122.215 196.135 ;
        RECT 112.910 194.885 113.805 195.260 ;
        RECT 114.315 195.215 114.705 195.295 ;
        RECT 111.855 194.455 112.740 194.625 ;
        RECT 112.920 194.155 113.235 194.655 ;
        RECT 113.465 194.325 113.805 194.885 ;
        RECT 113.975 194.155 114.145 195.165 ;
        RECT 114.315 194.370 114.645 195.215 ;
        RECT 118.280 194.590 118.630 195.840 ;
        RECT 114.875 194.155 120.220 194.590 ;
        RECT 120.395 194.155 120.685 195.320 ;
        RECT 120.860 195.295 121.030 195.965 ;
        RECT 121.285 195.795 121.455 195.965 ;
        RECT 121.200 195.465 121.455 195.795 ;
        RECT 121.680 195.465 121.875 195.795 ;
        RECT 120.860 194.325 121.195 195.295 ;
        RECT 121.365 194.155 121.535 195.295 ;
        RECT 121.705 194.495 121.875 195.465 ;
        RECT 122.045 194.835 122.215 195.965 ;
        RECT 122.385 195.175 122.555 195.975 ;
        RECT 122.760 195.685 123.035 196.535 ;
        RECT 122.755 195.515 123.035 195.685 ;
        RECT 122.760 195.375 123.035 195.515 ;
        RECT 123.205 195.175 123.395 196.535 ;
        RECT 123.575 196.170 124.085 196.705 ;
        RECT 124.305 195.895 124.550 196.500 ;
        RECT 125.965 196.050 126.295 196.485 ;
        RECT 126.465 196.095 126.635 196.705 ;
        RECT 125.915 195.965 126.295 196.050 ;
        RECT 126.805 195.965 127.135 196.490 ;
        RECT 127.395 196.175 127.605 196.705 ;
        RECT 127.880 196.255 128.665 196.425 ;
        RECT 128.835 196.255 129.240 196.425 ;
        RECT 125.915 195.925 126.140 195.965 ;
        RECT 123.595 195.725 124.825 195.895 ;
        RECT 122.385 195.005 123.395 195.175 ;
        RECT 123.565 195.160 124.315 195.350 ;
        RECT 122.045 194.665 123.170 194.835 ;
        RECT 123.565 194.495 123.735 195.160 ;
        RECT 124.485 194.915 124.825 195.725 ;
        RECT 125.915 195.345 126.085 195.925 ;
        RECT 126.805 195.795 127.005 195.965 ;
        RECT 127.880 195.795 128.050 196.255 ;
        RECT 126.255 195.465 127.005 195.795 ;
        RECT 127.175 195.465 128.050 195.795 ;
        RECT 125.915 195.295 126.130 195.345 ;
        RECT 125.915 195.215 126.305 195.295 ;
        RECT 121.705 194.325 123.735 194.495 ;
        RECT 123.905 194.155 124.075 194.915 ;
        RECT 124.310 194.505 124.825 194.915 ;
        RECT 125.975 194.370 126.305 195.215 ;
        RECT 126.815 195.260 127.005 195.465 ;
        RECT 126.475 194.155 126.645 195.165 ;
        RECT 126.815 194.885 127.710 195.260 ;
        RECT 126.815 194.325 127.155 194.885 ;
        RECT 127.385 194.155 127.700 194.655 ;
        RECT 127.880 194.625 128.050 195.465 ;
        RECT 128.220 195.755 128.685 196.085 ;
        RECT 129.070 196.025 129.240 196.255 ;
        RECT 129.420 196.205 129.790 196.705 ;
        RECT 130.110 196.255 130.785 196.425 ;
        RECT 130.980 196.255 131.315 196.425 ;
        RECT 128.220 194.795 128.540 195.755 ;
        RECT 129.070 195.725 129.900 196.025 ;
        RECT 128.710 194.825 128.900 195.545 ;
        RECT 129.070 194.655 129.240 195.725 ;
        RECT 129.700 195.695 129.900 195.725 ;
        RECT 129.410 195.475 129.580 195.545 ;
        RECT 130.110 195.475 130.280 196.255 ;
        RECT 131.145 196.115 131.315 196.255 ;
        RECT 131.485 196.245 131.735 196.705 ;
        RECT 129.410 195.305 130.280 195.475 ;
        RECT 130.450 195.835 130.975 196.055 ;
        RECT 131.145 195.985 131.370 196.115 ;
        RECT 129.410 195.215 129.920 195.305 ;
        RECT 127.880 194.455 128.765 194.625 ;
        RECT 128.990 194.325 129.240 194.655 ;
        RECT 129.410 194.155 129.580 194.955 ;
        RECT 129.750 194.600 129.920 195.215 ;
        RECT 130.450 195.135 130.620 195.835 ;
        RECT 130.090 194.770 130.620 195.135 ;
        RECT 130.790 195.070 131.030 195.665 ;
        RECT 131.200 194.880 131.370 195.985 ;
        RECT 131.540 195.125 131.820 196.075 ;
        RECT 131.065 194.750 131.370 194.880 ;
        RECT 129.750 194.430 130.855 194.600 ;
        RECT 131.065 194.325 131.315 194.750 ;
        RECT 131.485 194.155 131.750 194.615 ;
        RECT 131.990 194.325 132.175 196.445 ;
        RECT 132.345 196.325 132.675 196.705 ;
        RECT 132.845 196.155 133.015 196.445 ;
        RECT 133.280 196.305 133.615 196.705 ;
        RECT 132.350 195.985 133.015 196.155 ;
        RECT 133.785 196.135 133.990 196.535 ;
        RECT 134.200 196.225 134.475 196.705 ;
        RECT 134.685 196.205 134.945 196.535 ;
        RECT 132.350 194.995 132.580 195.985 ;
        RECT 133.305 195.965 133.990 196.135 ;
        RECT 132.750 195.165 133.100 195.815 ;
        RECT 132.350 194.825 133.015 194.995 ;
        RECT 132.345 194.155 132.675 194.655 ;
        RECT 132.845 194.325 133.015 194.825 ;
        RECT 133.305 194.935 133.645 195.965 ;
        RECT 133.815 195.295 134.065 195.795 ;
        RECT 134.245 195.465 134.605 196.045 ;
        RECT 134.775 195.295 134.945 196.205 ;
        RECT 135.115 196.160 140.460 196.705 ;
        RECT 136.700 195.330 137.040 196.160 ;
        RECT 140.635 195.935 144.145 196.705 ;
        RECT 144.315 195.955 145.525 196.705 ;
        RECT 145.695 195.955 146.905 196.705 ;
        RECT 133.815 195.125 134.945 195.295 ;
        RECT 133.305 194.760 133.970 194.935 ;
        RECT 133.280 194.155 133.615 194.580 ;
        RECT 133.785 194.355 133.970 194.760 ;
        RECT 134.175 194.155 134.505 194.935 ;
        RECT 134.675 194.355 134.945 195.125 ;
        RECT 138.520 194.590 138.870 195.840 ;
        RECT 140.635 195.415 142.285 195.935 ;
        RECT 142.455 195.245 144.145 195.765 ;
        RECT 144.315 195.415 144.835 195.955 ;
        RECT 145.005 195.245 145.525 195.785 ;
        RECT 135.115 194.155 140.460 194.590 ;
        RECT 140.635 194.155 144.145 195.245 ;
        RECT 144.315 194.155 145.525 195.245 ;
        RECT 145.695 195.245 146.215 195.785 ;
        RECT 146.385 195.415 146.905 195.955 ;
        RECT 145.695 194.155 146.905 195.245 ;
        RECT 17.270 193.985 146.990 194.155 ;
        RECT 17.355 192.895 18.565 193.985 ;
        RECT 18.735 192.895 22.245 193.985 ;
        RECT 17.355 192.185 17.875 192.725 ;
        RECT 18.045 192.355 18.565 192.895 ;
        RECT 18.735 192.205 20.385 192.725 ;
        RECT 20.555 192.375 22.245 192.895 ;
        RECT 22.875 193.115 23.150 193.815 ;
        RECT 23.320 193.440 23.575 193.985 ;
        RECT 23.745 193.475 24.225 193.815 ;
        RECT 24.400 193.430 25.005 193.985 ;
        RECT 24.390 193.330 25.005 193.430 ;
        RECT 24.390 193.305 24.575 193.330 ;
        RECT 17.355 191.435 18.565 192.185 ;
        RECT 18.735 191.435 22.245 192.205 ;
        RECT 22.875 192.085 23.045 193.115 ;
        RECT 23.320 192.985 24.075 193.235 ;
        RECT 24.245 193.060 24.575 193.305 ;
        RECT 23.320 192.950 24.090 192.985 ;
        RECT 23.320 192.940 24.105 192.950 ;
        RECT 23.215 192.925 24.110 192.940 ;
        RECT 23.215 192.910 24.130 192.925 ;
        RECT 23.215 192.900 24.150 192.910 ;
        RECT 23.215 192.890 24.175 192.900 ;
        RECT 23.215 192.860 24.245 192.890 ;
        RECT 23.215 192.830 24.265 192.860 ;
        RECT 23.215 192.800 24.285 192.830 ;
        RECT 23.215 192.775 24.315 192.800 ;
        RECT 23.215 192.740 24.350 192.775 ;
        RECT 23.215 192.735 24.380 192.740 ;
        RECT 23.215 192.340 23.445 192.735 ;
        RECT 23.990 192.730 24.380 192.735 ;
        RECT 24.015 192.720 24.380 192.730 ;
        RECT 24.030 192.715 24.380 192.720 ;
        RECT 24.045 192.710 24.380 192.715 ;
        RECT 24.745 192.710 25.005 193.160 ;
        RECT 24.045 192.705 25.005 192.710 ;
        RECT 24.055 192.695 25.005 192.705 ;
        RECT 24.065 192.690 25.005 192.695 ;
        RECT 24.075 192.680 25.005 192.690 ;
        RECT 24.080 192.670 25.005 192.680 ;
        RECT 24.085 192.665 25.005 192.670 ;
        RECT 24.095 192.650 25.005 192.665 ;
        RECT 24.100 192.635 25.005 192.650 ;
        RECT 24.110 192.610 25.005 192.635 ;
        RECT 23.615 192.140 23.945 192.565 ;
        RECT 22.875 191.605 23.135 192.085 ;
        RECT 23.305 191.435 23.555 191.975 ;
        RECT 23.725 191.655 23.945 192.140 ;
        RECT 24.115 192.540 25.005 192.610 ;
        RECT 26.095 193.115 26.370 193.815 ;
        RECT 26.540 193.440 26.795 193.985 ;
        RECT 26.965 193.475 27.445 193.815 ;
        RECT 27.620 193.430 28.225 193.985 ;
        RECT 27.610 193.330 28.225 193.430 ;
        RECT 27.610 193.305 27.795 193.330 ;
        RECT 24.115 191.815 24.285 192.540 ;
        RECT 24.455 191.985 25.005 192.370 ;
        RECT 26.095 192.085 26.265 193.115 ;
        RECT 26.540 192.985 27.295 193.235 ;
        RECT 27.465 193.060 27.795 193.305 ;
        RECT 26.540 192.950 27.310 192.985 ;
        RECT 26.540 192.940 27.325 192.950 ;
        RECT 26.435 192.925 27.330 192.940 ;
        RECT 26.435 192.910 27.350 192.925 ;
        RECT 26.435 192.900 27.370 192.910 ;
        RECT 26.435 192.890 27.395 192.900 ;
        RECT 26.435 192.860 27.465 192.890 ;
        RECT 26.435 192.830 27.485 192.860 ;
        RECT 26.435 192.800 27.505 192.830 ;
        RECT 26.435 192.775 27.535 192.800 ;
        RECT 26.435 192.740 27.570 192.775 ;
        RECT 26.435 192.735 27.600 192.740 ;
        RECT 26.435 192.340 26.665 192.735 ;
        RECT 27.210 192.730 27.600 192.735 ;
        RECT 27.235 192.720 27.600 192.730 ;
        RECT 27.250 192.715 27.600 192.720 ;
        RECT 27.265 192.710 27.600 192.715 ;
        RECT 27.965 192.710 28.225 193.160 ;
        RECT 28.435 192.845 28.665 193.985 ;
        RECT 28.835 192.835 29.165 193.815 ;
        RECT 29.335 192.845 29.545 193.985 ;
        RECT 27.265 192.705 28.225 192.710 ;
        RECT 27.275 192.695 28.225 192.705 ;
        RECT 27.285 192.690 28.225 192.695 ;
        RECT 27.295 192.680 28.225 192.690 ;
        RECT 27.300 192.670 28.225 192.680 ;
        RECT 27.305 192.665 28.225 192.670 ;
        RECT 27.315 192.650 28.225 192.665 ;
        RECT 27.320 192.635 28.225 192.650 ;
        RECT 27.330 192.610 28.225 192.635 ;
        RECT 26.835 192.140 27.165 192.565 ;
        RECT 24.115 191.645 25.005 191.815 ;
        RECT 26.095 191.605 26.355 192.085 ;
        RECT 26.525 191.435 26.775 191.975 ;
        RECT 26.945 191.655 27.165 192.140 ;
        RECT 27.335 192.540 28.225 192.610 ;
        RECT 27.335 191.815 27.505 192.540 ;
        RECT 28.415 192.425 28.745 192.675 ;
        RECT 27.675 191.985 28.225 192.370 ;
        RECT 27.335 191.645 28.225 191.815 ;
        RECT 28.435 191.435 28.665 192.255 ;
        RECT 28.915 192.235 29.165 192.835 ;
        RECT 30.235 192.820 30.525 193.985 ;
        RECT 30.695 193.550 36.040 193.985 ;
        RECT 28.835 191.605 29.165 192.235 ;
        RECT 29.335 191.435 29.545 192.255 ;
        RECT 30.235 191.435 30.525 192.160 ;
        RECT 32.280 191.980 32.620 192.810 ;
        RECT 34.100 192.300 34.450 193.550 ;
        RECT 36.215 192.895 37.425 193.985 ;
        RECT 36.215 192.185 36.735 192.725 ;
        RECT 36.905 192.355 37.425 192.895 ;
        RECT 37.605 193.645 38.775 193.815 ;
        RECT 37.605 192.975 37.935 193.645 ;
        RECT 38.445 193.605 38.775 193.645 ;
        RECT 38.945 193.605 39.320 193.985 ;
        RECT 38.105 193.435 38.335 193.475 ;
        RECT 38.105 193.385 38.720 193.435 ;
        RECT 39.465 193.385 39.635 193.515 ;
        RECT 38.105 193.185 39.635 193.385 ;
        RECT 39.870 193.205 40.135 193.985 ;
        RECT 38.105 193.145 38.985 193.185 ;
        RECT 39.125 192.975 40.185 193.015 ;
        RECT 37.605 192.845 40.185 192.975 ;
        RECT 40.355 192.845 40.635 193.985 ;
        RECT 37.605 192.795 39.350 192.845 ;
        RECT 30.695 191.435 36.040 191.980 ;
        RECT 36.215 191.435 37.425 192.185 ;
        RECT 37.635 192.115 38.085 192.625 ;
        RECT 38.275 192.425 38.750 192.625 ;
        RECT 38.500 192.025 38.750 192.425 ;
        RECT 39.000 192.425 39.350 192.625 ;
        RECT 39.000 192.025 39.210 192.425 ;
        RECT 39.520 192.345 39.845 192.675 ;
        RECT 40.015 192.175 40.185 192.845 ;
        RECT 40.805 192.835 41.135 193.815 ;
        RECT 41.305 192.845 41.565 193.985 ;
        RECT 41.735 193.265 42.195 193.815 ;
        RECT 42.385 193.265 42.715 193.985 ;
        RECT 40.365 192.405 40.700 192.675 ;
        RECT 40.870 192.235 41.040 192.835 ;
        RECT 41.210 192.425 41.545 192.675 ;
        RECT 39.455 192.005 40.185 192.175 ;
        RECT 37.605 191.435 38.055 191.945 ;
        RECT 39.455 191.855 39.635 192.005 ;
        RECT 38.330 191.605 39.635 191.855 ;
        RECT 39.815 191.435 40.145 191.835 ;
        RECT 40.355 191.435 40.665 192.235 ;
        RECT 40.870 191.605 41.565 192.235 ;
        RECT 41.735 191.895 41.985 193.265 ;
        RECT 42.915 193.095 43.215 193.645 ;
        RECT 43.385 193.315 43.665 193.985 ;
        RECT 42.275 192.925 43.215 193.095 ;
        RECT 42.275 192.675 42.445 192.925 ;
        RECT 43.585 192.675 43.850 193.035 ;
        RECT 42.155 192.345 42.445 192.675 ;
        RECT 42.615 192.425 42.955 192.675 ;
        RECT 43.175 192.425 43.850 192.675 ;
        RECT 44.035 192.965 44.410 193.815 ;
        RECT 44.580 193.185 44.830 193.985 ;
        RECT 45.000 193.355 45.250 193.815 ;
        RECT 45.420 193.525 45.670 193.985 ;
        RECT 45.840 193.355 46.090 193.815 ;
        RECT 46.260 193.525 46.510 193.985 ;
        RECT 46.680 193.355 46.930 193.815 ;
        RECT 47.100 193.525 47.350 193.985 ;
        RECT 47.520 193.355 47.770 193.815 ;
        RECT 45.000 193.135 47.770 193.355 ;
        RECT 47.985 193.355 48.300 193.815 ;
        RECT 48.470 193.525 48.720 193.985 ;
        RECT 48.890 193.355 49.140 193.815 ;
        RECT 49.310 193.525 49.560 193.985 ;
        RECT 49.730 193.565 51.700 193.815 ;
        RECT 49.730 193.355 49.940 193.565 ;
        RECT 51.910 193.395 52.200 193.815 ;
        RECT 47.985 193.135 49.940 193.355 ;
        RECT 50.110 193.135 52.200 193.395 ;
        RECT 52.370 193.185 52.620 193.985 ;
        RECT 45.000 192.965 45.250 193.135 ;
        RECT 51.910 193.015 52.200 193.135 ;
        RECT 52.790 193.015 53.040 193.815 ;
        RECT 53.210 193.185 53.460 193.985 ;
        RECT 53.630 193.015 53.985 193.815 ;
        RECT 44.035 192.795 45.250 192.965 ;
        RECT 45.635 192.795 49.680 192.965 ;
        RECT 49.850 192.795 51.720 192.965 ;
        RECT 51.910 192.795 53.985 193.015 ;
        RECT 54.155 192.895 55.825 193.985 ;
        RECT 42.275 192.255 42.445 192.345 ;
        RECT 44.035 192.255 44.270 192.795 ;
        RECT 45.635 192.625 45.805 192.795 ;
        RECT 49.510 192.625 49.680 192.795 ;
        RECT 51.550 192.625 51.720 192.795 ;
        RECT 44.440 192.425 45.805 192.625 ;
        RECT 46.125 192.425 49.340 192.625 ;
        RECT 49.510 192.425 51.380 192.625 ;
        RECT 51.550 192.425 53.595 192.625 ;
        RECT 53.765 192.255 53.985 192.795 ;
        RECT 42.275 192.065 43.665 192.255 ;
        RECT 41.735 191.605 42.295 191.895 ;
        RECT 42.465 191.435 42.715 191.895 ;
        RECT 43.335 191.705 43.665 192.065 ;
        RECT 44.035 191.995 45.710 192.255 ;
        RECT 45.880 192.075 47.810 192.255 ;
        RECT 45.880 191.825 46.130 192.075 ;
        RECT 44.120 191.605 46.130 191.825 ;
        RECT 46.300 191.435 46.470 191.905 ;
        RECT 46.640 191.605 46.970 192.075 ;
        RECT 47.140 191.435 47.310 191.905 ;
        RECT 47.480 191.605 47.810 192.075 ;
        RECT 47.985 191.435 48.260 192.255 ;
        RECT 48.430 192.085 52.160 192.255 ;
        RECT 48.430 192.075 51.380 192.085 ;
        RECT 48.430 191.605 48.760 192.075 ;
        RECT 48.930 191.435 49.100 191.905 ;
        RECT 49.270 191.605 49.600 192.075 ;
        RECT 49.770 191.435 49.940 191.905 ;
        RECT 50.110 191.605 50.440 192.075 ;
        RECT 50.610 191.435 50.780 191.905 ;
        RECT 50.950 191.605 51.280 192.075 ;
        RECT 51.450 191.435 51.720 191.905 ;
        RECT 51.910 191.825 52.160 192.085 ;
        RECT 52.330 191.995 53.985 192.255 ;
        RECT 54.155 192.205 54.905 192.725 ;
        RECT 55.075 192.375 55.825 192.895 ;
        RECT 55.995 192.820 56.285 193.985 ;
        RECT 56.460 193.595 56.795 193.815 ;
        RECT 57.800 193.605 58.155 193.985 ;
        RECT 56.460 192.975 56.715 193.595 ;
        RECT 56.965 193.435 57.195 193.475 ;
        RECT 58.325 193.435 58.575 193.815 ;
        RECT 56.965 193.235 58.575 193.435 ;
        RECT 56.965 193.145 57.150 193.235 ;
        RECT 57.740 193.225 58.575 193.235 ;
        RECT 58.825 193.205 59.075 193.985 ;
        RECT 59.245 193.135 59.505 193.815 ;
        RECT 57.305 193.035 57.635 193.065 ;
        RECT 57.305 192.975 59.105 193.035 ;
        RECT 56.460 192.865 59.165 192.975 ;
        RECT 56.460 192.805 57.635 192.865 ;
        RECT 58.965 192.830 59.165 192.865 ;
        RECT 56.455 192.425 56.945 192.625 ;
        RECT 57.135 192.425 57.610 192.635 ;
        RECT 51.910 191.655 53.920 191.825 ;
        RECT 54.155 191.435 55.825 192.205 ;
        RECT 55.995 191.435 56.285 192.160 ;
        RECT 56.460 191.435 56.915 192.200 ;
        RECT 57.390 192.025 57.610 192.425 ;
        RECT 57.855 192.425 58.185 192.635 ;
        RECT 57.855 192.025 58.065 192.425 ;
        RECT 58.355 192.390 58.765 192.695 ;
        RECT 58.995 192.255 59.165 192.830 ;
        RECT 58.895 192.135 59.165 192.255 ;
        RECT 58.320 192.090 59.165 192.135 ;
        RECT 58.320 191.965 59.075 192.090 ;
        RECT 58.320 191.815 58.490 191.965 ;
        RECT 59.335 191.935 59.505 193.135 ;
        RECT 57.190 191.605 58.490 191.815 ;
        RECT 58.745 191.435 59.075 191.795 ;
        RECT 59.245 191.605 59.505 191.935 ;
        RECT 59.675 193.265 60.135 193.815 ;
        RECT 60.325 193.265 60.655 193.985 ;
        RECT 59.675 191.895 59.925 193.265 ;
        RECT 60.855 193.095 61.155 193.645 ;
        RECT 61.325 193.315 61.605 193.985 ;
        RECT 61.975 193.550 67.320 193.985 ;
        RECT 60.215 192.925 61.155 193.095 ;
        RECT 60.215 192.675 60.385 192.925 ;
        RECT 61.525 192.675 61.790 193.035 ;
        RECT 60.095 192.345 60.385 192.675 ;
        RECT 60.555 192.425 60.895 192.675 ;
        RECT 61.115 192.425 61.790 192.675 ;
        RECT 60.215 192.255 60.385 192.345 ;
        RECT 60.215 192.065 61.605 192.255 ;
        RECT 59.675 191.605 60.235 191.895 ;
        RECT 60.405 191.435 60.655 191.895 ;
        RECT 61.275 191.705 61.605 192.065 ;
        RECT 63.560 191.980 63.900 192.810 ;
        RECT 65.380 192.300 65.730 193.550 ;
        RECT 67.495 192.895 71.005 193.985 ;
        RECT 71.175 192.895 72.385 193.985 ;
        RECT 72.555 193.475 72.855 193.985 ;
        RECT 73.025 193.305 73.355 193.815 ;
        RECT 73.525 193.475 74.155 193.985 ;
        RECT 74.735 193.475 75.115 193.645 ;
        RECT 75.285 193.475 75.585 193.985 ;
        RECT 74.945 193.305 75.115 193.475 ;
        RECT 67.495 192.205 69.145 192.725 ;
        RECT 69.315 192.375 71.005 192.895 ;
        RECT 61.975 191.435 67.320 191.980 ;
        RECT 67.495 191.435 71.005 192.205 ;
        RECT 71.175 192.185 71.695 192.725 ;
        RECT 71.865 192.355 72.385 192.895 ;
        RECT 72.555 193.135 74.775 193.305 ;
        RECT 71.175 191.435 72.385 192.185 ;
        RECT 72.555 192.175 72.725 193.135 ;
        RECT 72.895 192.795 74.435 192.965 ;
        RECT 72.895 192.345 73.140 192.795 ;
        RECT 73.400 192.425 74.095 192.625 ;
        RECT 74.265 192.595 74.435 192.795 ;
        RECT 74.605 192.935 74.775 193.135 ;
        RECT 74.945 193.105 75.605 193.305 ;
        RECT 76.945 193.255 77.240 193.985 ;
        RECT 74.605 192.765 75.265 192.935 ;
        RECT 74.265 192.425 74.865 192.595 ;
        RECT 75.095 192.345 75.265 192.765 ;
        RECT 72.555 191.630 73.020 192.175 ;
        RECT 73.525 191.435 73.695 192.255 ;
        RECT 73.865 192.175 74.775 192.255 ;
        RECT 75.435 192.175 75.605 193.105 ;
        RECT 77.410 193.085 77.670 193.810 ;
        RECT 77.840 193.255 78.100 193.985 ;
        RECT 78.270 193.085 78.530 193.810 ;
        RECT 78.700 193.255 78.960 193.985 ;
        RECT 79.130 193.085 79.390 193.810 ;
        RECT 79.560 193.255 79.820 193.985 ;
        RECT 79.990 193.085 80.250 193.810 ;
        RECT 73.865 192.085 75.115 192.175 ;
        RECT 73.865 191.605 74.195 192.085 ;
        RECT 74.605 192.005 75.115 192.085 ;
        RECT 74.365 191.435 74.715 191.825 ;
        RECT 74.885 191.605 75.115 192.005 ;
        RECT 75.285 191.695 75.605 192.175 ;
        RECT 76.940 192.845 80.250 193.085 ;
        RECT 80.420 192.875 80.680 193.985 ;
        RECT 76.940 192.255 77.910 192.845 ;
        RECT 80.850 192.675 81.100 193.810 ;
        RECT 81.280 192.875 81.575 193.985 ;
        RECT 81.755 192.820 82.045 193.985 ;
        RECT 82.215 193.550 87.560 193.985 ;
        RECT 78.080 192.425 81.100 192.675 ;
        RECT 76.940 192.085 80.250 192.255 ;
        RECT 76.940 191.435 77.240 191.915 ;
        RECT 77.410 191.630 77.670 192.085 ;
        RECT 77.840 191.435 78.100 191.915 ;
        RECT 78.270 191.630 78.530 192.085 ;
        RECT 78.700 191.435 78.960 191.915 ;
        RECT 79.130 191.630 79.390 192.085 ;
        RECT 79.560 191.435 79.820 191.915 ;
        RECT 79.990 191.630 80.250 192.085 ;
        RECT 80.420 191.435 80.680 191.960 ;
        RECT 80.850 191.615 81.100 192.425 ;
        RECT 81.270 192.065 81.585 192.675 ;
        RECT 81.280 191.435 81.525 191.895 ;
        RECT 81.755 191.435 82.045 192.160 ;
        RECT 83.800 191.980 84.140 192.810 ;
        RECT 85.620 192.300 85.970 193.550 ;
        RECT 87.735 192.895 91.245 193.985 ;
        RECT 87.735 192.205 89.385 192.725 ;
        RECT 89.555 192.375 91.245 192.895 ;
        RECT 91.415 192.845 91.800 193.815 ;
        RECT 91.970 193.525 92.295 193.985 ;
        RECT 92.815 193.355 93.095 193.815 ;
        RECT 91.970 193.135 93.095 193.355 ;
        RECT 82.215 191.435 87.560 191.980 ;
        RECT 87.735 191.435 91.245 192.205 ;
        RECT 91.415 192.175 91.695 192.845 ;
        RECT 91.970 192.675 92.420 193.135 ;
        RECT 93.285 192.965 93.685 193.815 ;
        RECT 94.085 193.525 94.355 193.985 ;
        RECT 94.525 193.355 94.810 193.815 ;
        RECT 91.865 192.345 92.420 192.675 ;
        RECT 92.590 192.405 93.685 192.965 ;
        RECT 91.970 192.235 92.420 192.345 ;
        RECT 91.415 191.605 91.800 192.175 ;
        RECT 91.970 192.065 93.095 192.235 ;
        RECT 91.970 191.435 92.295 191.895 ;
        RECT 92.815 191.605 93.095 192.065 ;
        RECT 93.285 191.605 93.685 192.405 ;
        RECT 93.855 193.135 94.810 193.355 ;
        RECT 95.185 193.315 95.355 193.815 ;
        RECT 95.525 193.485 95.855 193.985 ;
        RECT 95.185 193.145 95.850 193.315 ;
        RECT 93.855 192.235 94.065 193.135 ;
        RECT 94.235 192.405 94.925 192.965 ;
        RECT 95.100 192.325 95.450 192.975 ;
        RECT 93.855 192.065 94.810 192.235 ;
        RECT 95.620 192.155 95.850 193.145 ;
        RECT 94.085 191.435 94.355 191.895 ;
        RECT 94.525 191.605 94.810 192.065 ;
        RECT 95.185 191.985 95.850 192.155 ;
        RECT 95.185 191.695 95.355 191.985 ;
        RECT 95.525 191.435 95.855 191.815 ;
        RECT 96.025 191.695 96.210 193.815 ;
        RECT 96.450 193.525 96.715 193.985 ;
        RECT 96.885 193.390 97.135 193.815 ;
        RECT 97.345 193.540 98.450 193.710 ;
        RECT 96.830 193.260 97.135 193.390 ;
        RECT 96.380 192.065 96.660 193.015 ;
        RECT 96.830 192.155 97.000 193.260 ;
        RECT 97.170 192.475 97.410 193.070 ;
        RECT 97.580 193.005 98.110 193.370 ;
        RECT 97.580 192.305 97.750 193.005 ;
        RECT 98.280 192.925 98.450 193.540 ;
        RECT 98.620 193.185 98.790 193.985 ;
        RECT 98.960 193.485 99.210 193.815 ;
        RECT 99.435 193.515 100.320 193.685 ;
        RECT 98.280 192.835 98.790 192.925 ;
        RECT 96.830 192.025 97.055 192.155 ;
        RECT 97.225 192.085 97.750 192.305 ;
        RECT 97.920 192.665 98.790 192.835 ;
        RECT 96.465 191.435 96.715 191.895 ;
        RECT 96.885 191.885 97.055 192.025 ;
        RECT 97.920 191.885 98.090 192.665 ;
        RECT 98.620 192.595 98.790 192.665 ;
        RECT 98.300 192.415 98.500 192.445 ;
        RECT 98.960 192.415 99.130 193.485 ;
        RECT 99.300 192.595 99.490 193.315 ;
        RECT 98.300 192.115 99.130 192.415 ;
        RECT 99.660 192.385 99.980 193.345 ;
        RECT 96.885 191.715 97.220 191.885 ;
        RECT 97.415 191.715 98.090 191.885 ;
        RECT 98.410 191.435 98.780 191.935 ;
        RECT 98.960 191.885 99.130 192.115 ;
        RECT 99.515 192.055 99.980 192.385 ;
        RECT 100.150 192.675 100.320 193.515 ;
        RECT 100.500 193.485 100.815 193.985 ;
        RECT 101.045 193.255 101.385 193.815 ;
        RECT 100.490 192.880 101.385 193.255 ;
        RECT 101.555 192.975 101.725 193.985 ;
        RECT 101.195 192.675 101.385 192.880 ;
        RECT 101.895 192.925 102.225 193.770 ;
        RECT 101.895 192.845 102.285 192.925 ;
        RECT 102.070 192.795 102.285 192.845 ;
        RECT 100.150 192.345 101.025 192.675 ;
        RECT 101.195 192.345 101.945 192.675 ;
        RECT 100.150 191.885 100.320 192.345 ;
        RECT 101.195 192.175 101.395 192.345 ;
        RECT 102.115 192.215 102.285 192.795 ;
        RECT 102.060 192.175 102.285 192.215 ;
        RECT 98.960 191.715 99.365 191.885 ;
        RECT 99.535 191.715 100.320 191.885 ;
        RECT 100.595 191.435 100.805 191.965 ;
        RECT 101.065 191.650 101.395 192.175 ;
        RECT 101.905 192.090 102.285 192.175 ;
        RECT 102.460 192.845 102.795 193.815 ;
        RECT 102.965 192.845 103.135 193.985 ;
        RECT 103.305 193.645 105.335 193.815 ;
        RECT 102.460 192.175 102.630 192.845 ;
        RECT 103.305 192.675 103.475 193.645 ;
        RECT 102.800 192.345 103.055 192.675 ;
        RECT 103.280 192.345 103.475 192.675 ;
        RECT 103.645 193.305 104.770 193.475 ;
        RECT 102.885 192.175 103.055 192.345 ;
        RECT 103.645 192.175 103.815 193.305 ;
        RECT 101.565 191.435 101.735 192.045 ;
        RECT 101.905 191.655 102.235 192.090 ;
        RECT 102.460 191.605 102.715 192.175 ;
        RECT 102.885 192.005 103.815 192.175 ;
        RECT 103.985 192.965 104.995 193.135 ;
        RECT 103.985 192.165 104.155 192.965 ;
        RECT 104.360 192.285 104.635 192.765 ;
        RECT 104.355 192.115 104.635 192.285 ;
        RECT 103.640 191.970 103.815 192.005 ;
        RECT 102.885 191.435 103.215 191.835 ;
        RECT 103.640 191.605 104.170 191.970 ;
        RECT 104.360 191.605 104.635 192.115 ;
        RECT 104.805 191.605 104.995 192.965 ;
        RECT 105.165 192.980 105.335 193.645 ;
        RECT 105.505 193.225 105.675 193.985 ;
        RECT 105.910 193.225 106.425 193.635 ;
        RECT 105.165 192.790 105.915 192.980 ;
        RECT 106.085 192.415 106.425 193.225 ;
        RECT 107.515 192.820 107.805 193.985 ;
        RECT 108.065 193.315 108.235 193.815 ;
        RECT 108.405 193.485 108.735 193.985 ;
        RECT 108.065 193.145 108.730 193.315 ;
        RECT 105.195 192.245 106.425 192.415 ;
        RECT 107.980 192.325 108.330 192.975 ;
        RECT 105.175 191.435 105.685 191.970 ;
        RECT 105.905 191.640 106.150 192.245 ;
        RECT 107.515 191.435 107.805 192.160 ;
        RECT 108.500 192.155 108.730 193.145 ;
        RECT 108.065 191.985 108.730 192.155 ;
        RECT 108.065 191.695 108.235 191.985 ;
        RECT 108.405 191.435 108.735 191.815 ;
        RECT 108.905 191.695 109.090 193.815 ;
        RECT 109.330 193.525 109.595 193.985 ;
        RECT 109.765 193.390 110.015 193.815 ;
        RECT 110.225 193.540 111.330 193.710 ;
        RECT 109.710 193.260 110.015 193.390 ;
        RECT 109.260 192.065 109.540 193.015 ;
        RECT 109.710 192.155 109.880 193.260 ;
        RECT 110.050 192.475 110.290 193.070 ;
        RECT 110.460 193.005 110.990 193.370 ;
        RECT 110.460 192.305 110.630 193.005 ;
        RECT 111.160 192.925 111.330 193.540 ;
        RECT 111.500 193.185 111.670 193.985 ;
        RECT 111.840 193.485 112.090 193.815 ;
        RECT 112.315 193.515 113.200 193.685 ;
        RECT 111.160 192.835 111.670 192.925 ;
        RECT 109.710 192.025 109.935 192.155 ;
        RECT 110.105 192.085 110.630 192.305 ;
        RECT 110.800 192.665 111.670 192.835 ;
        RECT 109.345 191.435 109.595 191.895 ;
        RECT 109.765 191.885 109.935 192.025 ;
        RECT 110.800 191.885 110.970 192.665 ;
        RECT 111.500 192.595 111.670 192.665 ;
        RECT 111.180 192.415 111.380 192.445 ;
        RECT 111.840 192.415 112.010 193.485 ;
        RECT 112.180 192.595 112.370 193.315 ;
        RECT 111.180 192.115 112.010 192.415 ;
        RECT 112.540 192.385 112.860 193.345 ;
        RECT 109.765 191.715 110.100 191.885 ;
        RECT 110.295 191.715 110.970 191.885 ;
        RECT 111.290 191.435 111.660 191.935 ;
        RECT 111.840 191.885 112.010 192.115 ;
        RECT 112.395 192.055 112.860 192.385 ;
        RECT 113.030 192.675 113.200 193.515 ;
        RECT 113.380 193.485 113.695 193.985 ;
        RECT 113.925 193.255 114.265 193.815 ;
        RECT 113.370 192.880 114.265 193.255 ;
        RECT 114.435 192.975 114.605 193.985 ;
        RECT 114.075 192.675 114.265 192.880 ;
        RECT 114.775 192.925 115.105 193.770 ;
        RECT 114.775 192.845 115.165 192.925 ;
        RECT 115.335 192.895 117.925 193.985 ;
        RECT 114.950 192.795 115.165 192.845 ;
        RECT 113.030 192.345 113.905 192.675 ;
        RECT 114.075 192.345 114.825 192.675 ;
        RECT 113.030 191.885 113.200 192.345 ;
        RECT 114.075 192.175 114.275 192.345 ;
        RECT 114.995 192.215 115.165 192.795 ;
        RECT 114.940 192.175 115.165 192.215 ;
        RECT 111.840 191.715 112.245 191.885 ;
        RECT 112.415 191.715 113.200 191.885 ;
        RECT 113.475 191.435 113.685 191.965 ;
        RECT 113.945 191.650 114.275 192.175 ;
        RECT 114.785 192.090 115.165 192.175 ;
        RECT 115.335 192.205 116.545 192.725 ;
        RECT 116.715 192.375 117.925 192.895 ;
        RECT 118.100 192.845 118.435 193.815 ;
        RECT 118.605 192.845 118.775 193.985 ;
        RECT 118.945 193.645 120.975 193.815 ;
        RECT 114.445 191.435 114.615 192.045 ;
        RECT 114.785 191.655 115.115 192.090 ;
        RECT 115.335 191.435 117.925 192.205 ;
        RECT 118.100 192.175 118.270 192.845 ;
        RECT 118.945 192.675 119.115 193.645 ;
        RECT 118.440 192.345 118.695 192.675 ;
        RECT 118.920 192.345 119.115 192.675 ;
        RECT 119.285 193.305 120.410 193.475 ;
        RECT 118.525 192.175 118.695 192.345 ;
        RECT 119.285 192.175 119.455 193.305 ;
        RECT 118.100 191.605 118.355 192.175 ;
        RECT 118.525 192.005 119.455 192.175 ;
        RECT 119.625 192.965 120.635 193.135 ;
        RECT 119.625 192.165 119.795 192.965 ;
        RECT 119.280 191.970 119.455 192.005 ;
        RECT 118.525 191.435 118.855 191.835 ;
        RECT 119.280 191.605 119.810 191.970 ;
        RECT 120.000 191.945 120.275 192.765 ;
        RECT 119.995 191.775 120.275 191.945 ;
        RECT 120.000 191.605 120.275 191.775 ;
        RECT 120.445 191.605 120.635 192.965 ;
        RECT 120.805 192.980 120.975 193.645 ;
        RECT 121.145 193.225 121.315 193.985 ;
        RECT 121.550 193.225 122.065 193.635 ;
        RECT 120.805 192.790 121.555 192.980 ;
        RECT 121.725 192.415 122.065 193.225 ;
        RECT 122.350 193.355 122.635 193.815 ;
        RECT 122.805 193.525 123.075 193.985 ;
        RECT 122.350 193.135 123.305 193.355 ;
        RECT 120.835 192.245 122.065 192.415 ;
        RECT 122.235 192.405 122.925 192.965 ;
        RECT 120.815 191.435 121.325 191.970 ;
        RECT 121.545 191.640 121.790 192.245 ;
        RECT 123.095 192.235 123.305 193.135 ;
        RECT 122.350 192.065 123.305 192.235 ;
        RECT 123.475 192.965 123.875 193.815 ;
        RECT 124.065 193.355 124.345 193.815 ;
        RECT 124.865 193.525 125.190 193.985 ;
        RECT 124.065 193.135 125.190 193.355 ;
        RECT 123.475 192.405 124.570 192.965 ;
        RECT 124.740 192.675 125.190 193.135 ;
        RECT 125.360 192.845 125.745 193.815 ;
        RECT 125.915 192.895 127.125 193.985 ;
        RECT 127.410 193.355 127.695 193.815 ;
        RECT 127.865 193.525 128.135 193.985 ;
        RECT 127.410 193.135 128.365 193.355 ;
        RECT 122.350 191.605 122.635 192.065 ;
        RECT 122.805 191.435 123.075 191.895 ;
        RECT 123.475 191.605 123.875 192.405 ;
        RECT 124.740 192.345 125.295 192.675 ;
        RECT 124.740 192.235 125.190 192.345 ;
        RECT 124.065 192.065 125.190 192.235 ;
        RECT 125.465 192.175 125.745 192.845 ;
        RECT 124.065 191.605 124.345 192.065 ;
        RECT 124.865 191.435 125.190 191.895 ;
        RECT 125.360 191.605 125.745 192.175 ;
        RECT 125.915 192.185 126.435 192.725 ;
        RECT 126.605 192.355 127.125 192.895 ;
        RECT 127.295 192.405 127.985 192.965 ;
        RECT 128.155 192.235 128.365 193.135 ;
        RECT 125.915 191.435 127.125 192.185 ;
        RECT 127.410 192.065 128.365 192.235 ;
        RECT 128.535 192.965 128.935 193.815 ;
        RECT 129.125 193.355 129.405 193.815 ;
        RECT 129.925 193.525 130.250 193.985 ;
        RECT 129.125 193.135 130.250 193.355 ;
        RECT 128.535 192.405 129.630 192.965 ;
        RECT 129.800 192.675 130.250 193.135 ;
        RECT 130.420 192.845 130.805 193.815 ;
        RECT 131.065 193.055 131.235 193.815 ;
        RECT 131.450 193.225 131.780 193.985 ;
        RECT 131.065 192.885 131.780 193.055 ;
        RECT 131.950 192.910 132.205 193.815 ;
        RECT 127.410 191.605 127.695 192.065 ;
        RECT 127.865 191.435 128.135 191.895 ;
        RECT 128.535 191.605 128.935 192.405 ;
        RECT 129.800 192.345 130.355 192.675 ;
        RECT 129.800 192.235 130.250 192.345 ;
        RECT 129.125 192.065 130.250 192.235 ;
        RECT 130.525 192.175 130.805 192.845 ;
        RECT 130.975 192.335 131.330 192.705 ;
        RECT 131.610 192.675 131.780 192.885 ;
        RECT 131.610 192.345 131.865 192.675 ;
        RECT 129.125 191.605 129.405 192.065 ;
        RECT 129.925 191.435 130.250 191.895 ;
        RECT 130.420 191.605 130.805 192.175 ;
        RECT 131.610 192.155 131.780 192.345 ;
        RECT 132.035 192.180 132.205 192.910 ;
        RECT 132.380 192.835 132.640 193.985 ;
        RECT 133.275 192.820 133.565 193.985 ;
        RECT 133.735 193.135 133.995 193.815 ;
        RECT 134.165 193.205 134.415 193.985 ;
        RECT 134.665 193.435 134.915 193.815 ;
        RECT 135.085 193.605 135.440 193.985 ;
        RECT 136.445 193.595 136.780 193.815 ;
        RECT 136.045 193.435 136.275 193.475 ;
        RECT 134.665 193.235 136.275 193.435 ;
        RECT 134.665 193.225 135.500 193.235 ;
        RECT 136.090 193.145 136.275 193.235 ;
        RECT 131.065 191.985 131.780 192.155 ;
        RECT 131.065 191.605 131.235 191.985 ;
        RECT 131.450 191.435 131.780 191.815 ;
        RECT 131.950 191.605 132.205 192.180 ;
        RECT 132.380 191.435 132.640 192.275 ;
        RECT 133.275 191.435 133.565 192.160 ;
        RECT 133.735 191.935 133.905 193.135 ;
        RECT 135.605 193.035 135.935 193.065 ;
        RECT 134.135 192.975 135.935 193.035 ;
        RECT 136.525 192.975 136.780 193.595 ;
        RECT 136.955 193.550 142.300 193.985 ;
        RECT 134.075 192.865 136.780 192.975 ;
        RECT 134.075 192.830 134.275 192.865 ;
        RECT 134.075 192.255 134.245 192.830 ;
        RECT 135.605 192.805 136.780 192.865 ;
        RECT 134.475 192.390 134.885 192.695 ;
        RECT 135.055 192.425 135.385 192.635 ;
        RECT 134.075 192.135 134.345 192.255 ;
        RECT 134.075 192.090 134.920 192.135 ;
        RECT 134.165 191.965 134.920 192.090 ;
        RECT 135.175 192.025 135.385 192.425 ;
        RECT 135.630 192.425 136.105 192.635 ;
        RECT 136.295 192.425 136.785 192.625 ;
        RECT 135.630 192.025 135.850 192.425 ;
        RECT 133.735 191.605 133.995 191.935 ;
        RECT 134.750 191.815 134.920 191.965 ;
        RECT 134.165 191.435 134.495 191.795 ;
        RECT 134.750 191.605 136.050 191.815 ;
        RECT 136.325 191.435 136.780 192.200 ;
        RECT 138.540 191.980 138.880 192.810 ;
        RECT 140.360 192.300 140.710 193.550 ;
        RECT 142.475 192.895 145.065 193.985 ;
        RECT 142.475 192.205 143.685 192.725 ;
        RECT 143.855 192.375 145.065 192.895 ;
        RECT 145.695 192.895 146.905 193.985 ;
        RECT 145.695 192.355 146.215 192.895 ;
        RECT 136.955 191.435 142.300 191.980 ;
        RECT 142.475 191.435 145.065 192.205 ;
        RECT 146.385 192.185 146.905 192.725 ;
        RECT 145.695 191.435 146.905 192.185 ;
        RECT 17.270 191.265 146.990 191.435 ;
        RECT 17.355 190.515 18.565 191.265 ;
        RECT 18.735 190.720 24.080 191.265 ;
        RECT 17.355 189.975 17.875 190.515 ;
        RECT 18.045 189.805 18.565 190.345 ;
        RECT 20.320 189.890 20.660 190.720 ;
        RECT 24.715 190.465 25.025 191.265 ;
        RECT 25.230 190.465 25.925 191.095 ;
        RECT 26.095 190.720 31.440 191.265 ;
        RECT 17.355 188.715 18.565 189.805 ;
        RECT 22.140 189.150 22.490 190.400 ;
        RECT 24.725 190.025 25.060 190.295 ;
        RECT 25.230 189.865 25.400 190.465 ;
        RECT 25.570 190.025 25.905 190.275 ;
        RECT 27.680 189.890 28.020 190.720 ;
        RECT 31.615 190.495 35.125 191.265 ;
        RECT 18.735 188.715 24.080 189.150 ;
        RECT 24.715 188.715 24.995 189.855 ;
        RECT 25.165 188.885 25.495 189.865 ;
        RECT 25.665 188.715 25.925 189.855 ;
        RECT 29.500 189.150 29.850 190.400 ;
        RECT 31.615 189.975 33.265 190.495 ;
        RECT 35.500 190.485 36.000 191.095 ;
        RECT 33.435 189.805 35.125 190.325 ;
        RECT 35.295 190.025 35.645 190.275 ;
        RECT 35.830 189.855 36.000 190.485 ;
        RECT 36.630 190.615 36.960 191.095 ;
        RECT 37.130 190.805 37.355 191.265 ;
        RECT 37.525 190.615 37.855 191.095 ;
        RECT 36.630 190.445 37.855 190.615 ;
        RECT 38.045 190.465 38.295 191.265 ;
        RECT 38.465 190.465 38.805 191.095 ;
        RECT 39.180 190.485 39.680 191.095 ;
        RECT 38.575 190.415 38.805 190.465 ;
        RECT 36.170 190.075 36.500 190.275 ;
        RECT 36.670 190.075 37.000 190.275 ;
        RECT 37.170 190.075 37.590 190.275 ;
        RECT 37.765 190.105 38.460 190.275 ;
        RECT 37.765 189.855 37.935 190.105 ;
        RECT 38.630 189.855 38.805 190.415 ;
        RECT 38.975 190.025 39.325 190.275 ;
        RECT 39.510 189.855 39.680 190.485 ;
        RECT 40.310 190.615 40.640 191.095 ;
        RECT 40.810 190.805 41.035 191.265 ;
        RECT 41.205 190.615 41.535 191.095 ;
        RECT 40.310 190.445 41.535 190.615 ;
        RECT 41.725 190.465 41.975 191.265 ;
        RECT 42.145 190.465 42.485 191.095 ;
        RECT 43.115 190.540 43.405 191.265 ;
        RECT 43.635 190.805 43.880 191.265 ;
        RECT 39.850 190.075 40.180 190.275 ;
        RECT 40.350 190.075 40.680 190.275 ;
        RECT 40.850 190.075 41.270 190.275 ;
        RECT 41.445 190.105 42.140 190.275 ;
        RECT 41.445 189.855 41.615 190.105 ;
        RECT 42.310 189.855 42.485 190.465 ;
        RECT 43.575 190.025 43.890 190.635 ;
        RECT 44.060 190.275 44.310 191.085 ;
        RECT 44.480 190.740 44.740 191.265 ;
        RECT 44.910 190.615 45.170 191.070 ;
        RECT 45.340 190.785 45.600 191.265 ;
        RECT 45.770 190.615 46.030 191.070 ;
        RECT 46.200 190.785 46.460 191.265 ;
        RECT 46.630 190.615 46.890 191.070 ;
        RECT 47.060 190.785 47.320 191.265 ;
        RECT 47.490 190.615 47.750 191.070 ;
        RECT 47.920 190.785 48.220 191.265 ;
        RECT 48.680 190.805 48.945 191.265 ;
        RECT 49.315 190.625 49.485 191.095 ;
        RECT 49.735 190.805 49.905 191.265 ;
        RECT 50.155 190.625 50.325 191.095 ;
        RECT 50.575 190.805 50.745 191.265 ;
        RECT 50.995 190.625 51.165 191.095 ;
        RECT 51.335 190.800 51.585 191.265 ;
        RECT 44.910 190.445 48.220 190.615 ;
        RECT 49.315 190.445 51.685 190.625 ;
        RECT 52.525 190.575 52.855 191.265 ;
        RECT 53.315 190.670 53.935 191.095 ;
        RECT 54.105 190.775 54.435 191.265 ;
        RECT 44.060 190.025 47.080 190.275 ;
        RECT 26.095 188.715 31.440 189.150 ;
        RECT 31.615 188.715 35.125 189.805 ;
        RECT 35.500 189.685 37.935 189.855 ;
        RECT 35.500 188.885 35.830 189.685 ;
        RECT 36.000 188.715 36.330 189.515 ;
        RECT 36.630 188.885 36.960 189.685 ;
        RECT 37.605 188.715 37.855 189.515 ;
        RECT 38.125 188.715 38.295 189.855 ;
        RECT 38.465 188.885 38.805 189.855 ;
        RECT 39.180 189.685 41.615 189.855 ;
        RECT 39.180 188.885 39.510 189.685 ;
        RECT 39.680 188.715 40.010 189.515 ;
        RECT 40.310 188.885 40.640 189.685 ;
        RECT 41.285 188.715 41.535 189.515 ;
        RECT 41.805 188.715 41.975 189.855 ;
        RECT 42.145 188.885 42.485 189.855 ;
        RECT 43.115 188.715 43.405 189.880 ;
        RECT 43.585 188.715 43.880 189.825 ;
        RECT 44.060 188.890 44.310 190.025 ;
        RECT 47.250 189.855 48.220 190.445 ;
        RECT 48.655 190.025 51.165 190.275 ;
        RECT 51.335 189.855 51.685 190.445 ;
        RECT 53.575 190.335 53.935 190.670 ;
        RECT 52.515 190.055 53.935 190.335 ;
        RECT 44.480 188.715 44.740 189.825 ;
        RECT 44.910 189.615 48.220 189.855 ;
        RECT 44.910 188.890 45.170 189.615 ;
        RECT 45.340 188.715 45.600 189.445 ;
        RECT 45.770 188.890 46.030 189.615 ;
        RECT 46.200 188.715 46.460 189.445 ;
        RECT 46.630 188.890 46.890 189.615 ;
        RECT 47.060 188.715 47.320 189.445 ;
        RECT 47.490 188.890 47.750 189.615 ;
        RECT 47.920 188.715 48.215 189.445 ;
        RECT 48.680 188.715 48.975 189.855 ;
        RECT 49.235 189.685 51.685 189.855 ;
        RECT 49.235 188.885 49.565 189.685 ;
        RECT 49.735 188.715 49.905 189.515 ;
        RECT 50.075 188.885 50.405 189.685 ;
        RECT 50.915 189.665 51.685 189.685 ;
        RECT 50.575 188.715 50.745 189.515 ;
        RECT 50.915 188.885 51.245 189.665 ;
        RECT 51.415 188.715 51.585 189.175 ;
        RECT 51.985 188.715 52.315 189.885 ;
        RECT 52.515 188.885 52.845 190.055 ;
        RECT 53.045 188.715 53.375 189.885 ;
        RECT 53.575 188.885 53.935 190.055 ;
        RECT 54.105 190.025 54.445 190.605 ;
        RECT 54.615 190.495 56.285 191.265 ;
        RECT 54.615 189.975 55.365 190.495 ;
        RECT 56.495 190.445 56.725 191.265 ;
        RECT 56.895 190.465 57.225 191.095 ;
        RECT 54.105 188.715 54.435 189.855 ;
        RECT 55.535 189.805 56.285 190.325 ;
        RECT 56.475 190.025 56.805 190.275 ;
        RECT 56.975 189.865 57.225 190.465 ;
        RECT 57.395 190.445 57.605 191.265 ;
        RECT 57.860 190.865 58.190 191.265 ;
        RECT 58.360 190.695 58.530 190.965 ;
        RECT 58.700 190.755 59.015 191.265 ;
        RECT 59.245 190.755 59.535 191.095 ;
        RECT 59.705 190.755 59.945 191.265 ;
        RECT 60.605 190.765 60.935 191.265 ;
        RECT 57.835 190.525 58.530 190.695 ;
        RECT 54.615 188.715 56.285 189.805 ;
        RECT 56.495 188.715 56.725 189.855 ;
        RECT 56.895 188.885 57.225 189.865 ;
        RECT 57.395 188.715 57.605 189.855 ;
        RECT 57.835 189.515 58.265 190.525 ;
        RECT 58.435 189.855 58.605 190.355 ;
        RECT 58.775 190.025 59.185 190.585 ;
        RECT 59.355 189.855 59.535 190.755 ;
        RECT 61.135 190.695 61.305 191.045 ;
        RECT 61.505 190.865 61.835 191.265 ;
        RECT 62.005 190.695 62.175 191.045 ;
        RECT 62.345 190.865 62.725 191.265 ;
        RECT 59.705 190.415 59.905 190.585 ;
        RECT 59.705 190.025 59.900 190.415 ;
        RECT 60.600 190.025 60.950 190.595 ;
        RECT 61.135 190.525 62.745 190.695 ;
        RECT 62.915 190.590 63.185 190.935 ;
        RECT 62.575 190.355 62.745 190.525 ;
        RECT 61.120 189.905 61.830 190.355 ;
        RECT 62.000 190.025 62.405 190.355 ;
        RECT 62.575 190.025 62.845 190.355 ;
        RECT 58.435 189.685 59.895 189.855 ;
        RECT 57.835 189.345 58.610 189.515 ;
        RECT 57.940 188.715 58.110 189.175 ;
        RECT 58.280 188.885 58.610 189.345 ;
        RECT 58.780 188.715 58.950 189.515 ;
        RECT 59.535 189.510 59.895 189.685 ;
        RECT 60.600 189.565 60.920 189.855 ;
        RECT 61.115 189.735 61.830 189.905 ;
        RECT 62.575 189.855 62.745 190.025 ;
        RECT 63.015 189.855 63.185 190.590 ;
        RECT 63.360 190.500 63.815 191.265 ;
        RECT 64.090 190.885 65.390 191.095 ;
        RECT 65.645 190.905 65.975 191.265 ;
        RECT 65.220 190.735 65.390 190.885 ;
        RECT 66.145 190.765 66.405 191.095 ;
        RECT 66.175 190.755 66.405 190.765 ;
        RECT 66.740 190.755 66.980 191.265 ;
        RECT 67.160 190.755 67.440 191.085 ;
        RECT 67.670 190.755 67.885 191.265 ;
        RECT 64.290 190.275 64.510 190.675 ;
        RECT 63.355 190.075 63.845 190.275 ;
        RECT 64.035 190.065 64.510 190.275 ;
        RECT 64.755 190.275 64.965 190.675 ;
        RECT 65.220 190.610 65.975 190.735 ;
        RECT 65.220 190.565 66.065 190.610 ;
        RECT 65.795 190.445 66.065 190.565 ;
        RECT 64.755 190.065 65.085 190.275 ;
        RECT 65.255 190.005 65.665 190.310 ;
        RECT 62.020 189.685 62.745 189.855 ;
        RECT 62.020 189.565 62.190 189.685 ;
        RECT 60.600 189.395 62.190 189.565 ;
        RECT 60.600 188.935 62.255 189.225 ;
        RECT 62.425 188.715 62.705 189.515 ;
        RECT 62.915 188.885 63.185 189.855 ;
        RECT 63.360 189.835 64.535 189.895 ;
        RECT 65.895 189.870 66.065 190.445 ;
        RECT 65.865 189.835 66.065 189.870 ;
        RECT 63.360 189.725 66.065 189.835 ;
        RECT 63.360 189.105 63.615 189.725 ;
        RECT 64.205 189.665 66.005 189.725 ;
        RECT 64.205 189.635 64.535 189.665 ;
        RECT 66.235 189.565 66.405 190.755 ;
        RECT 66.635 190.025 66.990 190.585 ;
        RECT 67.160 189.855 67.330 190.755 ;
        RECT 67.500 190.025 67.765 190.585 ;
        RECT 68.055 190.525 68.670 191.095 ;
        RECT 68.875 190.540 69.165 191.265 ;
        RECT 69.345 190.535 69.645 191.265 ;
        RECT 68.015 189.855 68.185 190.355 ;
        RECT 63.865 189.465 64.050 189.555 ;
        RECT 64.640 189.465 65.475 189.475 ;
        RECT 63.865 189.265 65.475 189.465 ;
        RECT 63.865 189.225 64.095 189.265 ;
        RECT 63.360 188.885 63.695 189.105 ;
        RECT 64.700 188.715 65.055 189.095 ;
        RECT 65.225 188.885 65.475 189.265 ;
        RECT 65.725 188.715 65.975 189.495 ;
        RECT 66.145 188.885 66.405 189.565 ;
        RECT 66.760 189.685 68.185 189.855 ;
        RECT 66.760 189.510 67.150 189.685 ;
        RECT 67.635 188.715 67.965 189.515 ;
        RECT 68.355 189.505 68.670 190.525 ;
        RECT 69.825 190.355 70.055 190.975 ;
        RECT 70.255 190.705 70.480 191.085 ;
        RECT 70.650 190.875 70.980 191.265 ;
        RECT 71.175 190.885 72.065 191.055 ;
        RECT 70.255 190.525 70.585 190.705 ;
        RECT 69.350 190.025 69.645 190.355 ;
        RECT 69.825 190.025 70.240 190.355 ;
        RECT 68.135 188.885 68.670 189.505 ;
        RECT 68.875 188.715 69.165 189.880 ;
        RECT 70.410 189.855 70.585 190.525 ;
        RECT 70.755 190.025 70.995 190.675 ;
        RECT 71.175 190.330 71.725 190.715 ;
        RECT 71.895 190.160 72.065 190.885 ;
        RECT 71.175 190.090 72.065 190.160 ;
        RECT 72.235 190.560 72.455 191.045 ;
        RECT 72.625 190.725 72.875 191.265 ;
        RECT 73.045 190.615 73.305 191.095 ;
        RECT 72.235 190.135 72.565 190.560 ;
        RECT 71.175 190.065 72.070 190.090 ;
        RECT 71.175 190.050 72.080 190.065 ;
        RECT 71.175 190.035 72.085 190.050 ;
        RECT 71.175 190.030 72.095 190.035 ;
        RECT 71.175 190.020 72.100 190.030 ;
        RECT 71.175 190.010 72.105 190.020 ;
        RECT 71.175 190.005 72.115 190.010 ;
        RECT 71.175 189.995 72.125 190.005 ;
        RECT 71.175 189.990 72.135 189.995 ;
        RECT 69.345 189.495 70.240 189.825 ;
        RECT 70.410 189.665 70.995 189.855 ;
        RECT 69.345 189.325 70.550 189.495 ;
        RECT 69.345 188.895 69.675 189.325 ;
        RECT 69.855 188.715 70.050 189.155 ;
        RECT 70.220 188.895 70.550 189.325 ;
        RECT 70.720 188.895 70.995 189.665 ;
        RECT 71.175 189.540 71.435 189.990 ;
        RECT 71.800 189.985 72.135 189.990 ;
        RECT 71.800 189.980 72.150 189.985 ;
        RECT 71.800 189.970 72.165 189.980 ;
        RECT 71.800 189.965 72.190 189.970 ;
        RECT 72.735 189.965 72.965 190.360 ;
        RECT 71.800 189.960 72.965 189.965 ;
        RECT 71.830 189.925 72.965 189.960 ;
        RECT 71.865 189.900 72.965 189.925 ;
        RECT 71.895 189.870 72.965 189.900 ;
        RECT 71.915 189.840 72.965 189.870 ;
        RECT 71.935 189.810 72.965 189.840 ;
        RECT 72.005 189.800 72.965 189.810 ;
        RECT 72.030 189.790 72.965 189.800 ;
        RECT 72.050 189.775 72.965 189.790 ;
        RECT 72.070 189.760 72.965 189.775 ;
        RECT 72.075 189.750 72.860 189.760 ;
        RECT 72.090 189.715 72.860 189.750 ;
        RECT 71.605 189.395 71.935 189.640 ;
        RECT 72.105 189.465 72.860 189.715 ;
        RECT 73.135 189.585 73.305 190.615 ;
        RECT 71.605 189.370 71.790 189.395 ;
        RECT 71.175 189.270 71.790 189.370 ;
        RECT 71.175 188.715 71.780 189.270 ;
        RECT 71.955 188.885 72.435 189.225 ;
        RECT 72.605 188.715 72.860 189.260 ;
        RECT 73.030 188.885 73.305 189.585 ;
        RECT 73.475 190.525 73.860 191.095 ;
        RECT 74.030 190.805 74.355 191.265 ;
        RECT 74.875 190.635 75.155 191.095 ;
        RECT 73.475 189.855 73.755 190.525 ;
        RECT 74.030 190.465 75.155 190.635 ;
        RECT 74.030 190.355 74.480 190.465 ;
        RECT 73.925 190.025 74.480 190.355 ;
        RECT 75.345 190.295 75.745 191.095 ;
        RECT 76.145 190.805 76.415 191.265 ;
        RECT 76.585 190.635 76.870 191.095 ;
        RECT 78.095 190.795 78.390 191.265 ;
        RECT 73.475 188.885 73.860 189.855 ;
        RECT 74.030 189.565 74.480 190.025 ;
        RECT 74.650 189.735 75.745 190.295 ;
        RECT 74.030 189.345 75.155 189.565 ;
        RECT 74.030 188.715 74.355 189.175 ;
        RECT 74.875 188.885 75.155 189.345 ;
        RECT 75.345 188.885 75.745 189.735 ;
        RECT 75.915 190.465 76.870 190.635 ;
        RECT 78.560 190.625 78.820 191.070 ;
        RECT 78.990 190.795 79.250 191.265 ;
        RECT 79.420 190.625 79.675 191.070 ;
        RECT 79.845 190.795 80.145 191.265 ;
        RECT 75.915 189.565 76.125 190.465 ;
        RECT 77.635 190.455 80.665 190.625 ;
        RECT 80.855 190.455 81.095 191.265 ;
        RECT 81.265 190.455 81.595 191.095 ;
        RECT 81.765 190.455 82.035 191.265 ;
        RECT 82.215 190.720 87.560 191.265 ;
        RECT 76.295 189.735 76.985 190.295 ;
        RECT 77.635 189.890 77.805 190.455 ;
        RECT 77.975 190.060 80.190 190.285 ;
        RECT 80.365 189.890 80.665 190.455 ;
        RECT 80.835 190.025 81.185 190.275 ;
        RECT 77.635 189.720 80.665 189.890 ;
        RECT 81.355 189.855 81.525 190.455 ;
        RECT 81.695 190.025 82.045 190.275 ;
        RECT 83.800 189.890 84.140 190.720 ;
        RECT 88.660 190.525 88.915 191.095 ;
        RECT 89.085 190.865 89.415 191.265 ;
        RECT 89.840 190.730 90.370 191.095 ;
        RECT 89.840 190.695 90.015 190.730 ;
        RECT 89.085 190.525 90.015 190.695 ;
        RECT 75.915 189.345 76.870 189.565 ;
        RECT 76.145 188.715 76.415 189.175 ;
        RECT 76.585 188.885 76.870 189.345 ;
        RECT 77.615 188.715 77.960 189.550 ;
        RECT 78.135 188.915 78.390 189.720 ;
        RECT 78.560 188.715 78.820 189.550 ;
        RECT 78.995 188.915 79.250 189.720 ;
        RECT 79.420 188.715 79.680 189.550 ;
        RECT 79.850 188.915 80.110 189.720 ;
        RECT 80.845 189.685 81.525 189.855 ;
        RECT 80.280 188.715 80.665 189.550 ;
        RECT 80.845 188.900 81.175 189.685 ;
        RECT 81.705 188.715 82.035 189.855 ;
        RECT 85.620 189.150 85.970 190.400 ;
        RECT 88.660 189.855 88.830 190.525 ;
        RECT 89.085 190.355 89.255 190.525 ;
        RECT 89.000 190.025 89.255 190.355 ;
        RECT 89.480 190.025 89.675 190.355 ;
        RECT 82.215 188.715 87.560 189.150 ;
        RECT 88.660 188.885 88.995 189.855 ;
        RECT 89.165 188.715 89.335 189.855 ;
        RECT 89.505 189.055 89.675 190.025 ;
        RECT 89.845 189.395 90.015 190.525 ;
        RECT 90.185 189.735 90.355 190.535 ;
        RECT 90.560 190.245 90.835 191.095 ;
        RECT 90.555 190.075 90.835 190.245 ;
        RECT 90.560 189.935 90.835 190.075 ;
        RECT 91.005 189.735 91.195 191.095 ;
        RECT 91.375 190.730 91.885 191.265 ;
        RECT 92.105 190.455 92.350 191.060 ;
        RECT 92.795 190.495 94.465 191.265 ;
        RECT 94.635 190.540 94.925 191.265 ;
        RECT 95.560 190.525 95.815 191.095 ;
        RECT 95.985 190.865 96.315 191.265 ;
        RECT 96.740 190.730 97.270 191.095 ;
        RECT 96.740 190.695 96.915 190.730 ;
        RECT 95.985 190.525 96.915 190.695 ;
        RECT 91.395 190.285 92.625 190.455 ;
        RECT 90.185 189.565 91.195 189.735 ;
        RECT 91.365 189.720 92.115 189.910 ;
        RECT 89.845 189.225 90.970 189.395 ;
        RECT 91.365 189.055 91.535 189.720 ;
        RECT 92.285 189.475 92.625 190.285 ;
        RECT 92.795 189.975 93.545 190.495 ;
        RECT 93.715 189.805 94.465 190.325 ;
        RECT 89.505 188.885 91.535 189.055 ;
        RECT 91.705 188.715 91.875 189.475 ;
        RECT 92.110 189.065 92.625 189.475 ;
        RECT 92.795 188.715 94.465 189.805 ;
        RECT 94.635 188.715 94.925 189.880 ;
        RECT 95.560 189.855 95.730 190.525 ;
        RECT 95.985 190.355 96.155 190.525 ;
        RECT 95.900 190.025 96.155 190.355 ;
        RECT 96.380 190.025 96.575 190.355 ;
        RECT 95.560 188.885 95.895 189.855 ;
        RECT 96.065 188.715 96.235 189.855 ;
        RECT 96.405 189.055 96.575 190.025 ;
        RECT 96.745 189.395 96.915 190.525 ;
        RECT 97.085 189.735 97.255 190.535 ;
        RECT 97.460 190.245 97.735 191.095 ;
        RECT 97.455 190.075 97.735 190.245 ;
        RECT 97.460 189.935 97.735 190.075 ;
        RECT 97.905 189.735 98.095 191.095 ;
        RECT 98.275 190.730 98.785 191.265 ;
        RECT 99.005 190.455 99.250 191.060 ;
        RECT 99.810 190.635 100.095 191.095 ;
        RECT 100.265 190.805 100.535 191.265 ;
        RECT 99.810 190.465 100.765 190.635 ;
        RECT 98.295 190.285 99.525 190.455 ;
        RECT 97.085 189.565 98.095 189.735 ;
        RECT 98.265 189.720 99.015 189.910 ;
        RECT 96.745 189.225 97.870 189.395 ;
        RECT 98.265 189.055 98.435 189.720 ;
        RECT 99.185 189.475 99.525 190.285 ;
        RECT 99.695 189.735 100.385 190.295 ;
        RECT 100.555 189.565 100.765 190.465 ;
        RECT 96.405 188.885 98.435 189.055 ;
        RECT 98.605 188.715 98.775 189.475 ;
        RECT 99.010 189.065 99.525 189.475 ;
        RECT 99.810 189.345 100.765 189.565 ;
        RECT 100.935 190.295 101.335 191.095 ;
        RECT 101.525 190.635 101.805 191.095 ;
        RECT 102.325 190.805 102.650 191.265 ;
        RECT 101.525 190.465 102.650 190.635 ;
        RECT 102.820 190.525 103.205 191.095 ;
        RECT 102.200 190.355 102.650 190.465 ;
        RECT 100.935 189.735 102.030 190.295 ;
        RECT 102.200 190.025 102.755 190.355 ;
        RECT 99.810 188.885 100.095 189.345 ;
        RECT 100.265 188.715 100.535 189.175 ;
        RECT 100.935 188.885 101.335 189.735 ;
        RECT 102.200 189.565 102.650 190.025 ;
        RECT 102.925 189.855 103.205 190.525 ;
        RECT 103.490 190.635 103.775 191.095 ;
        RECT 103.945 190.805 104.215 191.265 ;
        RECT 103.490 190.465 104.445 190.635 ;
        RECT 101.525 189.345 102.650 189.565 ;
        RECT 101.525 188.885 101.805 189.345 ;
        RECT 102.325 188.715 102.650 189.175 ;
        RECT 102.820 188.885 103.205 189.855 ;
        RECT 103.375 189.735 104.065 190.295 ;
        RECT 104.235 189.565 104.445 190.465 ;
        RECT 103.490 189.345 104.445 189.565 ;
        RECT 104.615 190.295 105.015 191.095 ;
        RECT 105.205 190.635 105.485 191.095 ;
        RECT 106.005 190.805 106.330 191.265 ;
        RECT 105.205 190.465 106.330 190.635 ;
        RECT 106.500 190.525 106.885 191.095 ;
        RECT 105.880 190.355 106.330 190.465 ;
        RECT 104.615 189.735 105.710 190.295 ;
        RECT 105.880 190.025 106.435 190.355 ;
        RECT 103.490 188.885 103.775 189.345 ;
        RECT 103.945 188.715 104.215 189.175 ;
        RECT 104.615 188.885 105.015 189.735 ;
        RECT 105.880 189.565 106.330 190.025 ;
        RECT 106.605 189.855 106.885 190.525 ;
        RECT 107.055 190.515 108.265 191.265 ;
        RECT 108.440 190.525 108.695 191.095 ;
        RECT 108.865 190.865 109.195 191.265 ;
        RECT 109.620 190.730 110.150 191.095 ;
        RECT 110.340 190.925 110.615 191.095 ;
        RECT 110.335 190.755 110.615 190.925 ;
        RECT 109.620 190.695 109.795 190.730 ;
        RECT 108.865 190.525 109.795 190.695 ;
        RECT 107.055 189.975 107.575 190.515 ;
        RECT 105.205 189.345 106.330 189.565 ;
        RECT 105.205 188.885 105.485 189.345 ;
        RECT 106.005 188.715 106.330 189.175 ;
        RECT 106.500 188.885 106.885 189.855 ;
        RECT 107.745 189.805 108.265 190.345 ;
        RECT 107.055 188.715 108.265 189.805 ;
        RECT 108.440 189.855 108.610 190.525 ;
        RECT 108.865 190.355 109.035 190.525 ;
        RECT 108.780 190.025 109.035 190.355 ;
        RECT 109.260 190.025 109.455 190.355 ;
        RECT 108.440 188.885 108.775 189.855 ;
        RECT 108.945 188.715 109.115 189.855 ;
        RECT 109.285 189.055 109.455 190.025 ;
        RECT 109.625 189.395 109.795 190.525 ;
        RECT 109.965 189.735 110.135 190.535 ;
        RECT 110.340 189.935 110.615 190.755 ;
        RECT 110.785 189.735 110.975 191.095 ;
        RECT 111.155 190.730 111.665 191.265 ;
        RECT 111.885 190.455 112.130 191.060 ;
        RECT 112.575 190.525 112.960 191.095 ;
        RECT 113.130 190.805 113.455 191.265 ;
        RECT 113.975 190.635 114.255 191.095 ;
        RECT 111.175 190.285 112.405 190.455 ;
        RECT 109.965 189.565 110.975 189.735 ;
        RECT 111.145 189.720 111.895 189.910 ;
        RECT 109.625 189.225 110.750 189.395 ;
        RECT 111.145 189.055 111.315 189.720 ;
        RECT 112.065 189.475 112.405 190.285 ;
        RECT 109.285 188.885 111.315 189.055 ;
        RECT 111.485 188.715 111.655 189.475 ;
        RECT 111.890 189.065 112.405 189.475 ;
        RECT 112.575 189.855 112.855 190.525 ;
        RECT 113.130 190.465 114.255 190.635 ;
        RECT 113.130 190.355 113.580 190.465 ;
        RECT 113.025 190.025 113.580 190.355 ;
        RECT 114.445 190.295 114.845 191.095 ;
        RECT 115.245 190.805 115.515 191.265 ;
        RECT 115.685 190.635 115.970 191.095 ;
        RECT 112.575 188.885 112.960 189.855 ;
        RECT 113.130 189.565 113.580 190.025 ;
        RECT 113.750 189.735 114.845 190.295 ;
        RECT 113.130 189.345 114.255 189.565 ;
        RECT 113.130 188.715 113.455 189.175 ;
        RECT 113.975 188.885 114.255 189.345 ;
        RECT 114.445 188.885 114.845 189.735 ;
        RECT 115.015 190.465 115.970 190.635 ;
        RECT 116.260 190.525 116.515 191.095 ;
        RECT 116.685 190.865 117.015 191.265 ;
        RECT 117.440 190.730 117.970 191.095 ;
        RECT 117.440 190.695 117.615 190.730 ;
        RECT 116.685 190.525 117.615 190.695 ;
        RECT 115.015 189.565 115.225 190.465 ;
        RECT 115.395 189.735 116.085 190.295 ;
        RECT 116.260 189.855 116.430 190.525 ;
        RECT 116.685 190.355 116.855 190.525 ;
        RECT 116.600 190.025 116.855 190.355 ;
        RECT 117.080 190.025 117.275 190.355 ;
        RECT 115.015 189.345 115.970 189.565 ;
        RECT 115.245 188.715 115.515 189.175 ;
        RECT 115.685 188.885 115.970 189.345 ;
        RECT 116.260 188.885 116.595 189.855 ;
        RECT 116.765 188.715 116.935 189.855 ;
        RECT 117.105 189.055 117.275 190.025 ;
        RECT 117.445 189.395 117.615 190.525 ;
        RECT 117.785 189.735 117.955 190.535 ;
        RECT 118.160 190.245 118.435 191.095 ;
        RECT 118.155 190.075 118.435 190.245 ;
        RECT 118.160 189.935 118.435 190.075 ;
        RECT 118.605 189.735 118.795 191.095 ;
        RECT 118.975 190.730 119.485 191.265 ;
        RECT 119.705 190.455 119.950 191.060 ;
        RECT 120.395 190.540 120.685 191.265 ;
        RECT 120.945 190.715 121.115 191.005 ;
        RECT 121.285 190.885 121.615 191.265 ;
        RECT 120.945 190.545 121.610 190.715 ;
        RECT 118.995 190.285 120.225 190.455 ;
        RECT 117.785 189.565 118.795 189.735 ;
        RECT 118.965 189.720 119.715 189.910 ;
        RECT 117.445 189.225 118.570 189.395 ;
        RECT 118.965 189.055 119.135 189.720 ;
        RECT 119.885 189.475 120.225 190.285 ;
        RECT 117.105 188.885 119.135 189.055 ;
        RECT 119.305 188.715 119.475 189.475 ;
        RECT 119.710 189.065 120.225 189.475 ;
        RECT 120.395 188.715 120.685 189.880 ;
        RECT 120.860 189.725 121.210 190.375 ;
        RECT 121.380 189.555 121.610 190.545 ;
        RECT 120.945 189.385 121.610 189.555 ;
        RECT 120.945 188.885 121.115 189.385 ;
        RECT 121.285 188.715 121.615 189.215 ;
        RECT 121.785 188.885 121.970 191.005 ;
        RECT 122.225 190.805 122.475 191.265 ;
        RECT 122.645 190.815 122.980 190.985 ;
        RECT 123.175 190.815 123.850 190.985 ;
        RECT 122.645 190.675 122.815 190.815 ;
        RECT 122.140 189.685 122.420 190.635 ;
        RECT 122.590 190.545 122.815 190.675 ;
        RECT 122.590 189.440 122.760 190.545 ;
        RECT 122.985 190.395 123.510 190.615 ;
        RECT 122.930 189.630 123.170 190.225 ;
        RECT 123.340 189.695 123.510 190.395 ;
        RECT 123.680 190.035 123.850 190.815 ;
        RECT 124.170 190.765 124.540 191.265 ;
        RECT 124.720 190.815 125.125 190.985 ;
        RECT 125.295 190.815 126.080 190.985 ;
        RECT 124.720 190.585 124.890 190.815 ;
        RECT 124.060 190.285 124.890 190.585 ;
        RECT 125.275 190.315 125.740 190.645 ;
        RECT 124.060 190.255 124.260 190.285 ;
        RECT 124.380 190.035 124.550 190.105 ;
        RECT 123.680 189.865 124.550 190.035 ;
        RECT 124.040 189.775 124.550 189.865 ;
        RECT 122.590 189.310 122.895 189.440 ;
        RECT 123.340 189.330 123.870 189.695 ;
        RECT 122.210 188.715 122.475 189.175 ;
        RECT 122.645 188.885 122.895 189.310 ;
        RECT 124.040 189.160 124.210 189.775 ;
        RECT 123.105 188.990 124.210 189.160 ;
        RECT 124.380 188.715 124.550 189.515 ;
        RECT 124.720 189.215 124.890 190.285 ;
        RECT 125.060 189.385 125.250 190.105 ;
        RECT 125.420 189.355 125.740 190.315 ;
        RECT 125.910 190.355 126.080 190.815 ;
        RECT 126.355 190.735 126.565 191.265 ;
        RECT 126.825 190.525 127.155 191.050 ;
        RECT 127.325 190.655 127.495 191.265 ;
        RECT 127.665 190.610 127.995 191.045 ;
        RECT 127.665 190.525 128.045 190.610 ;
        RECT 126.955 190.355 127.155 190.525 ;
        RECT 127.820 190.485 128.045 190.525 ;
        RECT 125.910 190.025 126.785 190.355 ;
        RECT 126.955 190.025 127.705 190.355 ;
        RECT 124.720 188.885 124.970 189.215 ;
        RECT 125.910 189.185 126.080 190.025 ;
        RECT 126.955 189.820 127.145 190.025 ;
        RECT 127.875 189.905 128.045 190.485 ;
        RECT 127.830 189.855 128.045 189.905 ;
        RECT 126.250 189.445 127.145 189.820 ;
        RECT 127.655 189.775 128.045 189.855 ;
        RECT 128.215 190.525 128.600 191.095 ;
        RECT 128.770 190.805 129.095 191.265 ;
        RECT 129.615 190.635 129.895 191.095 ;
        RECT 128.215 189.855 128.495 190.525 ;
        RECT 128.770 190.465 129.895 190.635 ;
        RECT 128.770 190.355 129.220 190.465 ;
        RECT 128.665 190.025 129.220 190.355 ;
        RECT 130.085 190.295 130.485 191.095 ;
        RECT 130.885 190.805 131.155 191.265 ;
        RECT 131.325 190.635 131.610 191.095 ;
        RECT 132.060 190.755 132.300 191.265 ;
        RECT 132.480 190.755 132.760 191.085 ;
        RECT 132.990 190.755 133.205 191.265 ;
        RECT 125.195 189.015 126.080 189.185 ;
        RECT 126.260 188.715 126.575 189.215 ;
        RECT 126.805 188.885 127.145 189.445 ;
        RECT 127.315 188.715 127.485 189.725 ;
        RECT 127.655 188.930 127.985 189.775 ;
        RECT 128.215 188.885 128.600 189.855 ;
        RECT 128.770 189.565 129.220 190.025 ;
        RECT 129.390 189.735 130.485 190.295 ;
        RECT 128.770 189.345 129.895 189.565 ;
        RECT 128.770 188.715 129.095 189.175 ;
        RECT 129.615 188.885 129.895 189.345 ;
        RECT 130.085 188.885 130.485 189.735 ;
        RECT 130.655 190.465 131.610 190.635 ;
        RECT 130.655 189.565 130.865 190.465 ;
        RECT 131.035 189.735 131.725 190.295 ;
        RECT 131.955 190.025 132.310 190.585 ;
        RECT 132.480 189.855 132.650 190.755 ;
        RECT 132.820 190.025 133.085 190.585 ;
        RECT 133.375 190.525 133.990 191.095 ;
        RECT 134.245 190.610 134.575 191.045 ;
        RECT 134.745 190.655 134.915 191.265 ;
        RECT 133.335 189.855 133.505 190.355 ;
        RECT 132.080 189.685 133.505 189.855 ;
        RECT 130.655 189.345 131.610 189.565 ;
        RECT 132.080 189.510 132.470 189.685 ;
        RECT 130.885 188.715 131.155 189.175 ;
        RECT 131.325 188.885 131.610 189.345 ;
        RECT 132.955 188.715 133.285 189.515 ;
        RECT 133.675 189.505 133.990 190.525 ;
        RECT 134.195 190.525 134.575 190.610 ;
        RECT 135.085 190.525 135.415 191.050 ;
        RECT 135.675 190.735 135.885 191.265 ;
        RECT 136.160 190.815 136.945 190.985 ;
        RECT 137.115 190.815 137.520 190.985 ;
        RECT 134.195 190.485 134.420 190.525 ;
        RECT 134.195 189.905 134.365 190.485 ;
        RECT 135.085 190.355 135.285 190.525 ;
        RECT 136.160 190.355 136.330 190.815 ;
        RECT 134.535 190.025 135.285 190.355 ;
        RECT 135.455 190.025 136.330 190.355 ;
        RECT 134.195 189.855 134.410 189.905 ;
        RECT 134.195 189.775 134.585 189.855 ;
        RECT 133.455 188.885 133.990 189.505 ;
        RECT 134.255 188.930 134.585 189.775 ;
        RECT 135.095 189.820 135.285 190.025 ;
        RECT 134.755 188.715 134.925 189.725 ;
        RECT 135.095 189.445 135.990 189.820 ;
        RECT 135.095 188.885 135.435 189.445 ;
        RECT 135.665 188.715 135.980 189.215 ;
        RECT 136.160 189.185 136.330 190.025 ;
        RECT 136.500 190.315 136.965 190.645 ;
        RECT 137.350 190.585 137.520 190.815 ;
        RECT 137.700 190.765 138.070 191.265 ;
        RECT 138.390 190.815 139.065 190.985 ;
        RECT 139.260 190.815 139.595 190.985 ;
        RECT 136.500 189.355 136.820 190.315 ;
        RECT 137.350 190.285 138.180 190.585 ;
        RECT 136.990 189.385 137.180 190.105 ;
        RECT 137.350 189.215 137.520 190.285 ;
        RECT 137.980 190.255 138.180 190.285 ;
        RECT 137.690 190.035 137.860 190.105 ;
        RECT 138.390 190.035 138.560 190.815 ;
        RECT 139.425 190.675 139.595 190.815 ;
        RECT 139.765 190.805 140.015 191.265 ;
        RECT 137.690 189.865 138.560 190.035 ;
        RECT 138.730 190.395 139.255 190.615 ;
        RECT 139.425 190.545 139.650 190.675 ;
        RECT 137.690 189.775 138.200 189.865 ;
        RECT 136.160 189.015 137.045 189.185 ;
        RECT 137.270 188.885 137.520 189.215 ;
        RECT 137.690 188.715 137.860 189.515 ;
        RECT 138.030 189.160 138.200 189.775 ;
        RECT 138.730 189.695 138.900 190.395 ;
        RECT 138.370 189.330 138.900 189.695 ;
        RECT 139.070 189.630 139.310 190.225 ;
        RECT 139.480 189.440 139.650 190.545 ;
        RECT 139.820 189.685 140.100 190.635 ;
        RECT 139.345 189.310 139.650 189.440 ;
        RECT 138.030 188.990 139.135 189.160 ;
        RECT 139.345 188.885 139.595 189.310 ;
        RECT 139.765 188.715 140.030 189.175 ;
        RECT 140.270 188.885 140.455 191.005 ;
        RECT 140.625 190.885 140.955 191.265 ;
        RECT 141.125 190.715 141.295 191.005 ;
        RECT 140.630 190.545 141.295 190.715 ;
        RECT 140.630 189.555 140.860 190.545 ;
        RECT 141.555 190.495 145.065 191.265 ;
        RECT 145.695 190.515 146.905 191.265 ;
        RECT 141.030 189.725 141.380 190.375 ;
        RECT 141.555 189.975 143.205 190.495 ;
        RECT 143.375 189.805 145.065 190.325 ;
        RECT 140.630 189.385 141.295 189.555 ;
        RECT 140.625 188.715 140.955 189.215 ;
        RECT 141.125 188.885 141.295 189.385 ;
        RECT 141.555 188.715 145.065 189.805 ;
        RECT 145.695 189.805 146.215 190.345 ;
        RECT 146.385 189.975 146.905 190.515 ;
        RECT 145.695 188.715 146.905 189.805 ;
        RECT 17.270 188.545 146.990 188.715 ;
        RECT 17.355 187.455 18.565 188.545 ;
        RECT 18.735 187.455 22.245 188.545 ;
        RECT 17.355 186.745 17.875 187.285 ;
        RECT 18.045 186.915 18.565 187.455 ;
        RECT 18.735 186.765 20.385 187.285 ;
        RECT 20.555 186.935 22.245 187.455 ;
        RECT 22.415 187.675 22.690 188.375 ;
        RECT 22.860 188.000 23.115 188.545 ;
        RECT 23.285 188.035 23.765 188.375 ;
        RECT 23.940 187.990 24.545 188.545 ;
        RECT 23.930 187.890 24.545 187.990 ;
        RECT 23.930 187.865 24.115 187.890 ;
        RECT 17.355 185.995 18.565 186.745 ;
        RECT 18.735 185.995 22.245 186.765 ;
        RECT 22.415 186.645 22.585 187.675 ;
        RECT 22.860 187.545 23.615 187.795 ;
        RECT 23.785 187.620 24.115 187.865 ;
        RECT 22.860 187.510 23.630 187.545 ;
        RECT 22.860 187.500 23.645 187.510 ;
        RECT 22.755 187.485 23.650 187.500 ;
        RECT 22.755 187.470 23.670 187.485 ;
        RECT 22.755 187.460 23.690 187.470 ;
        RECT 22.755 187.450 23.715 187.460 ;
        RECT 22.755 187.420 23.785 187.450 ;
        RECT 22.755 187.390 23.805 187.420 ;
        RECT 22.755 187.360 23.825 187.390 ;
        RECT 22.755 187.335 23.855 187.360 ;
        RECT 22.755 187.300 23.890 187.335 ;
        RECT 22.755 187.295 23.920 187.300 ;
        RECT 22.755 186.900 22.985 187.295 ;
        RECT 23.530 187.290 23.920 187.295 ;
        RECT 23.555 187.280 23.920 187.290 ;
        RECT 23.570 187.275 23.920 187.280 ;
        RECT 23.585 187.270 23.920 187.275 ;
        RECT 24.285 187.270 24.545 187.720 ;
        RECT 24.900 187.575 25.290 187.750 ;
        RECT 25.775 187.745 26.105 188.545 ;
        RECT 26.275 187.755 26.810 188.375 ;
        RECT 24.900 187.405 26.325 187.575 ;
        RECT 23.585 187.265 24.545 187.270 ;
        RECT 23.595 187.255 24.545 187.265 ;
        RECT 23.605 187.250 24.545 187.255 ;
        RECT 23.615 187.240 24.545 187.250 ;
        RECT 23.620 187.230 24.545 187.240 ;
        RECT 23.625 187.225 24.545 187.230 ;
        RECT 23.635 187.210 24.545 187.225 ;
        RECT 23.640 187.195 24.545 187.210 ;
        RECT 23.650 187.170 24.545 187.195 ;
        RECT 23.155 186.700 23.485 187.125 ;
        RECT 22.415 186.165 22.675 186.645 ;
        RECT 22.845 185.995 23.095 186.535 ;
        RECT 23.265 186.215 23.485 186.700 ;
        RECT 23.655 187.100 24.545 187.170 ;
        RECT 23.655 186.375 23.825 187.100 ;
        RECT 23.995 186.545 24.545 186.930 ;
        RECT 24.775 186.675 25.130 187.235 ;
        RECT 25.300 186.505 25.470 187.405 ;
        RECT 25.640 186.675 25.905 187.235 ;
        RECT 26.155 186.905 26.325 187.405 ;
        RECT 26.495 186.735 26.810 187.755 ;
        RECT 27.055 187.405 27.285 188.545 ;
        RECT 27.455 187.395 27.785 188.375 ;
        RECT 27.955 187.405 28.165 188.545 ;
        RECT 28.395 187.405 28.655 188.545 ;
        RECT 28.825 187.395 29.155 188.375 ;
        RECT 29.325 187.405 29.605 188.545 ;
        RECT 27.035 186.985 27.365 187.235 ;
        RECT 23.655 186.205 24.545 186.375 ;
        RECT 24.880 185.995 25.120 186.505 ;
        RECT 25.300 186.175 25.580 186.505 ;
        RECT 25.810 185.995 26.025 186.505 ;
        RECT 26.195 186.165 26.810 186.735 ;
        RECT 27.055 185.995 27.285 186.815 ;
        RECT 27.535 186.795 27.785 187.395 ;
        RECT 28.415 186.985 28.750 187.235 ;
        RECT 27.455 186.165 27.785 186.795 ;
        RECT 27.955 185.995 28.165 186.815 ;
        RECT 28.920 186.795 29.090 187.395 ;
        RECT 30.235 187.380 30.525 188.545 ;
        RECT 30.695 187.455 34.205 188.545 ;
        RECT 29.260 186.965 29.595 187.235 ;
        RECT 28.395 186.165 29.090 186.795 ;
        RECT 29.295 185.995 29.605 186.795 ;
        RECT 30.695 186.765 32.345 187.285 ;
        RECT 32.515 186.935 34.205 187.455 ;
        RECT 35.040 187.575 35.370 188.375 ;
        RECT 35.540 187.745 35.870 188.545 ;
        RECT 36.170 187.575 36.500 188.375 ;
        RECT 37.145 187.745 37.395 188.545 ;
        RECT 35.040 187.405 37.475 187.575 ;
        RECT 37.665 187.405 37.835 188.545 ;
        RECT 38.005 187.405 38.345 188.375 ;
        RECT 38.515 187.405 38.795 188.545 ;
        RECT 34.835 186.985 35.185 187.235 ;
        RECT 35.370 186.775 35.540 187.405 ;
        RECT 35.710 186.985 36.040 187.185 ;
        RECT 36.210 186.985 36.540 187.185 ;
        RECT 36.710 186.985 37.130 187.185 ;
        RECT 37.305 187.155 37.475 187.405 ;
        RECT 37.305 186.985 38.000 187.155 ;
        RECT 30.235 185.995 30.525 186.720 ;
        RECT 30.695 185.995 34.205 186.765 ;
        RECT 35.040 186.165 35.540 186.775 ;
        RECT 36.170 186.645 37.395 186.815 ;
        RECT 38.170 186.795 38.345 187.405 ;
        RECT 38.965 187.395 39.295 188.375 ;
        RECT 39.465 187.405 39.725 188.545 ;
        RECT 39.895 187.405 40.155 188.545 ;
        RECT 40.395 188.035 42.010 188.365 ;
        RECT 38.525 186.965 38.860 187.235 ;
        RECT 39.030 186.845 39.200 187.395 ;
        RECT 40.405 187.235 40.575 187.795 ;
        RECT 40.835 187.695 42.010 187.865 ;
        RECT 42.180 187.745 42.460 188.545 ;
        RECT 40.835 187.405 41.165 187.695 ;
        RECT 41.840 187.575 42.010 187.695 ;
        RECT 41.335 187.235 41.580 187.525 ;
        RECT 41.840 187.405 42.500 187.575 ;
        RECT 42.670 187.405 42.945 188.375 ;
        RECT 43.365 187.815 43.660 188.545 ;
        RECT 43.830 187.645 44.090 188.370 ;
        RECT 44.260 187.815 44.520 188.545 ;
        RECT 44.690 187.645 44.950 188.370 ;
        RECT 45.120 187.815 45.380 188.545 ;
        RECT 45.550 187.645 45.810 188.370 ;
        RECT 45.980 187.815 46.240 188.545 ;
        RECT 46.410 187.645 46.670 188.370 ;
        RECT 42.330 187.235 42.500 187.405 ;
        RECT 39.370 186.985 39.705 187.235 ;
        RECT 39.900 186.985 40.235 187.235 ;
        RECT 40.405 186.905 41.120 187.235 ;
        RECT 41.335 186.905 42.160 187.235 ;
        RECT 42.330 186.905 42.605 187.235 ;
        RECT 39.030 186.795 39.205 186.845 ;
        RECT 40.405 186.815 40.655 186.905 ;
        RECT 36.170 186.165 36.500 186.645 ;
        RECT 36.670 185.995 36.895 186.455 ;
        RECT 37.065 186.165 37.395 186.645 ;
        RECT 37.585 185.995 37.835 186.795 ;
        RECT 38.005 186.165 38.345 186.795 ;
        RECT 38.515 185.995 38.825 186.795 ;
        RECT 39.030 186.165 39.725 186.795 ;
        RECT 39.895 185.995 40.155 186.815 ;
        RECT 40.325 186.395 40.655 186.815 ;
        RECT 42.330 186.735 42.500 186.905 ;
        RECT 40.835 186.565 42.500 186.735 ;
        RECT 42.775 186.670 42.945 187.405 ;
        RECT 40.835 186.165 41.095 186.565 ;
        RECT 41.265 185.995 41.595 186.395 ;
        RECT 41.765 186.215 41.935 186.565 ;
        RECT 42.105 185.995 42.480 186.395 ;
        RECT 42.670 186.325 42.945 186.670 ;
        RECT 43.360 187.405 46.670 187.645 ;
        RECT 46.840 187.435 47.100 188.545 ;
        RECT 43.360 186.815 44.330 187.405 ;
        RECT 47.270 187.235 47.520 188.370 ;
        RECT 47.700 187.435 47.995 188.545 ;
        RECT 48.175 188.110 53.520 188.545 ;
        RECT 44.500 186.985 47.520 187.235 ;
        RECT 43.360 186.645 46.670 186.815 ;
        RECT 43.360 185.995 43.660 186.475 ;
        RECT 43.830 186.190 44.090 186.645 ;
        RECT 44.260 185.995 44.520 186.475 ;
        RECT 44.690 186.190 44.950 186.645 ;
        RECT 45.120 185.995 45.380 186.475 ;
        RECT 45.550 186.190 45.810 186.645 ;
        RECT 45.980 185.995 46.240 186.475 ;
        RECT 46.410 186.190 46.670 186.645 ;
        RECT 46.840 185.995 47.100 186.520 ;
        RECT 47.270 186.175 47.520 186.985 ;
        RECT 47.690 186.625 48.005 187.235 ;
        RECT 49.760 186.540 50.100 187.370 ;
        RECT 51.580 186.860 51.930 188.110 ;
        RECT 53.695 187.455 55.365 188.545 ;
        RECT 53.695 186.765 54.445 187.285 ;
        RECT 54.615 186.935 55.365 187.455 ;
        RECT 55.995 187.380 56.285 188.545 ;
        RECT 56.920 187.405 57.240 188.545 ;
        RECT 57.420 187.235 57.615 188.285 ;
        RECT 57.795 187.695 58.125 188.375 ;
        RECT 58.325 187.745 58.580 188.545 ;
        RECT 57.795 187.415 58.145 187.695 ;
        RECT 58.920 187.635 59.170 188.365 ;
        RECT 59.340 187.815 59.670 188.545 ;
        RECT 59.840 187.635 60.025 188.365 ;
        RECT 56.980 187.185 57.240 187.235 ;
        RECT 56.975 187.015 57.240 187.185 ;
        RECT 56.980 186.905 57.240 187.015 ;
        RECT 57.420 186.905 57.805 187.235 ;
        RECT 57.975 187.035 58.145 187.415 ;
        RECT 58.335 187.205 58.580 187.565 ;
        RECT 58.920 187.435 60.025 187.635 ;
        RECT 60.195 187.235 60.425 188.365 ;
        RECT 60.605 187.695 61.330 188.365 ;
        RECT 57.975 186.865 58.495 187.035 ;
        RECT 47.700 185.995 47.945 186.455 ;
        RECT 48.175 185.995 53.520 186.540 ;
        RECT 53.695 185.995 55.365 186.765 ;
        RECT 55.995 185.995 56.285 186.720 ;
        RECT 56.920 186.525 58.135 186.695 ;
        RECT 56.920 186.175 57.210 186.525 ;
        RECT 57.405 185.995 57.735 186.355 ;
        RECT 57.905 186.220 58.135 186.525 ;
        RECT 58.325 186.300 58.495 186.865 ;
        RECT 58.765 186.675 59.105 187.235 ;
        RECT 59.275 186.905 59.915 187.235 ;
        RECT 60.095 186.905 60.425 187.235 ;
        RECT 60.605 186.905 60.905 187.525 ;
        RECT 58.755 185.995 59.095 186.505 ;
        RECT 59.275 186.175 59.525 186.905 ;
        RECT 61.115 186.725 61.330 187.695 ;
        RECT 61.515 187.575 61.805 188.375 ;
        RECT 61.975 187.745 62.210 188.545 ;
        RECT 62.395 188.205 63.930 188.375 ;
        RECT 62.395 187.575 62.725 188.205 ;
        RECT 61.515 187.405 62.725 187.575 ;
        RECT 61.515 186.905 61.760 187.235 ;
        RECT 61.930 186.735 62.100 187.405 ;
        RECT 62.895 187.235 63.130 187.980 ;
        RECT 62.270 186.905 62.670 187.235 ;
        RECT 62.840 186.905 63.130 187.235 ;
        RECT 63.320 187.235 63.590 187.980 ;
        RECT 63.760 187.575 63.930 188.205 ;
        RECT 64.100 187.745 64.505 188.545 ;
        RECT 63.760 187.405 64.505 187.575 ;
        RECT 63.320 186.905 63.660 187.235 ;
        RECT 63.830 186.905 64.165 187.235 ;
        RECT 64.335 186.905 64.505 187.405 ;
        RECT 64.675 186.980 65.025 188.375 ;
        RECT 65.195 188.110 70.540 188.545 ;
        RECT 59.850 186.535 61.330 186.725 ;
        RECT 59.850 186.175 60.035 186.535 ;
        RECT 60.215 185.995 60.545 186.365 ;
        RECT 60.725 186.175 60.950 186.535 ;
        RECT 61.515 186.165 62.100 186.735 ;
        RECT 62.350 186.565 63.745 186.735 ;
        RECT 62.350 186.220 62.680 186.565 ;
        RECT 62.895 185.995 63.270 186.395 ;
        RECT 63.450 186.220 63.745 186.565 ;
        RECT 63.915 185.995 64.585 186.735 ;
        RECT 64.755 186.165 65.025 186.980 ;
        RECT 66.780 186.540 67.120 187.370 ;
        RECT 68.600 186.860 68.950 188.110 ;
        RECT 70.715 187.455 71.925 188.545 ;
        RECT 70.715 186.745 71.235 187.285 ;
        RECT 71.405 186.915 71.925 187.455 ;
        RECT 72.100 188.190 73.180 188.360 ;
        RECT 72.100 187.405 72.435 188.190 ;
        RECT 72.605 187.235 72.840 187.915 ;
        RECT 73.010 187.575 73.180 188.190 ;
        RECT 73.445 187.745 73.760 188.545 ;
        RECT 73.010 187.405 73.325 187.575 ;
        RECT 72.100 186.905 72.435 187.235 ;
        RECT 72.605 186.905 72.985 187.235 ;
        RECT 65.195 185.995 70.540 186.540 ;
        RECT 70.715 185.995 71.925 186.745 ;
        RECT 73.155 186.735 73.325 187.405 ;
        RECT 72.100 186.565 73.325 186.735 ;
        RECT 73.495 186.565 73.765 187.575 ;
        RECT 73.995 187.485 74.325 188.330 ;
        RECT 74.495 187.535 74.665 188.545 ;
        RECT 74.835 187.815 75.175 188.375 ;
        RECT 75.405 188.045 75.720 188.545 ;
        RECT 75.900 188.075 76.785 188.245 ;
        RECT 73.935 187.405 74.325 187.485 ;
        RECT 74.835 187.440 75.730 187.815 ;
        RECT 73.935 187.355 74.150 187.405 ;
        RECT 73.935 186.775 74.105 187.355 ;
        RECT 74.835 187.235 75.025 187.440 ;
        RECT 75.900 187.235 76.070 188.075 ;
        RECT 77.010 188.045 77.260 188.375 ;
        RECT 74.275 186.905 75.025 187.235 ;
        RECT 75.195 186.905 76.070 187.235 ;
        RECT 73.935 186.735 74.160 186.775 ;
        RECT 74.825 186.735 75.025 186.905 ;
        RECT 73.935 186.650 74.315 186.735 ;
        RECT 72.100 186.295 72.355 186.565 ;
        RECT 72.525 185.995 72.855 186.395 ;
        RECT 73.025 186.295 73.195 186.565 ;
        RECT 73.365 185.995 73.695 186.395 ;
        RECT 73.985 186.215 74.315 186.650 ;
        RECT 74.485 185.995 74.655 186.605 ;
        RECT 74.825 186.210 75.155 186.735 ;
        RECT 75.415 185.995 75.625 186.525 ;
        RECT 75.900 186.445 76.070 186.905 ;
        RECT 76.240 186.945 76.560 187.905 ;
        RECT 76.730 187.155 76.920 187.875 ;
        RECT 77.090 186.975 77.260 188.045 ;
        RECT 77.430 187.745 77.600 188.545 ;
        RECT 77.770 188.100 78.875 188.270 ;
        RECT 77.770 187.485 77.940 188.100 ;
        RECT 79.085 187.950 79.335 188.375 ;
        RECT 79.505 188.085 79.770 188.545 ;
        RECT 78.110 187.565 78.640 187.930 ;
        RECT 79.085 187.820 79.390 187.950 ;
        RECT 77.430 187.395 77.940 187.485 ;
        RECT 77.430 187.225 78.300 187.395 ;
        RECT 77.430 187.155 77.600 187.225 ;
        RECT 77.720 186.975 77.920 187.005 ;
        RECT 76.240 186.615 76.705 186.945 ;
        RECT 77.090 186.675 77.920 186.975 ;
        RECT 77.090 186.445 77.260 186.675 ;
        RECT 75.900 186.275 76.685 186.445 ;
        RECT 76.855 186.275 77.260 186.445 ;
        RECT 77.440 185.995 77.810 186.495 ;
        RECT 78.130 186.445 78.300 187.225 ;
        RECT 78.470 186.865 78.640 187.565 ;
        RECT 78.810 187.035 79.050 187.630 ;
        RECT 78.470 186.645 78.995 186.865 ;
        RECT 79.220 186.715 79.390 187.820 ;
        RECT 79.165 186.585 79.390 186.715 ;
        RECT 79.560 186.625 79.840 187.575 ;
        RECT 79.165 186.445 79.335 186.585 ;
        RECT 78.130 186.275 78.805 186.445 ;
        RECT 79.000 186.275 79.335 186.445 ;
        RECT 79.505 185.995 79.755 186.455 ;
        RECT 80.010 186.255 80.195 188.375 ;
        RECT 80.365 188.045 80.695 188.545 ;
        RECT 80.865 187.875 81.035 188.375 ;
        RECT 80.370 187.705 81.035 187.875 ;
        RECT 80.370 186.715 80.600 187.705 ;
        RECT 80.770 186.885 81.120 187.535 ;
        RECT 81.755 187.380 82.045 188.545 ;
        RECT 82.215 187.455 83.885 188.545 ;
        RECT 84.605 187.875 84.775 188.375 ;
        RECT 84.945 188.045 85.275 188.545 ;
        RECT 84.605 187.705 85.270 187.875 ;
        RECT 82.215 186.765 82.965 187.285 ;
        RECT 83.135 186.935 83.885 187.455 ;
        RECT 84.520 186.885 84.870 187.535 ;
        RECT 80.370 186.545 81.035 186.715 ;
        RECT 80.365 185.995 80.695 186.375 ;
        RECT 80.865 186.255 81.035 186.545 ;
        RECT 81.755 185.995 82.045 186.720 ;
        RECT 82.215 185.995 83.885 186.765 ;
        RECT 85.040 186.715 85.270 187.705 ;
        RECT 84.605 186.545 85.270 186.715 ;
        RECT 84.605 186.255 84.775 186.545 ;
        RECT 84.945 185.995 85.275 186.375 ;
        RECT 85.445 186.255 85.630 188.375 ;
        RECT 85.870 188.085 86.135 188.545 ;
        RECT 86.305 187.950 86.555 188.375 ;
        RECT 86.765 188.100 87.870 188.270 ;
        RECT 86.250 187.820 86.555 187.950 ;
        RECT 85.800 186.625 86.080 187.575 ;
        RECT 86.250 186.715 86.420 187.820 ;
        RECT 86.590 187.035 86.830 187.630 ;
        RECT 87.000 187.565 87.530 187.930 ;
        RECT 87.000 186.865 87.170 187.565 ;
        RECT 87.700 187.485 87.870 188.100 ;
        RECT 88.040 187.745 88.210 188.545 ;
        RECT 88.380 188.045 88.630 188.375 ;
        RECT 88.855 188.075 89.740 188.245 ;
        RECT 87.700 187.395 88.210 187.485 ;
        RECT 86.250 186.585 86.475 186.715 ;
        RECT 86.645 186.645 87.170 186.865 ;
        RECT 87.340 187.225 88.210 187.395 ;
        RECT 85.885 185.995 86.135 186.455 ;
        RECT 86.305 186.445 86.475 186.585 ;
        RECT 87.340 186.445 87.510 187.225 ;
        RECT 88.040 187.155 88.210 187.225 ;
        RECT 87.720 186.975 87.920 187.005 ;
        RECT 88.380 186.975 88.550 188.045 ;
        RECT 88.720 187.155 88.910 187.875 ;
        RECT 87.720 186.675 88.550 186.975 ;
        RECT 89.080 186.945 89.400 187.905 ;
        RECT 86.305 186.275 86.640 186.445 ;
        RECT 86.835 186.275 87.510 186.445 ;
        RECT 87.830 185.995 88.200 186.495 ;
        RECT 88.380 186.445 88.550 186.675 ;
        RECT 88.935 186.615 89.400 186.945 ;
        RECT 89.570 187.235 89.740 188.075 ;
        RECT 89.920 188.045 90.235 188.545 ;
        RECT 90.465 187.815 90.805 188.375 ;
        RECT 89.910 187.440 90.805 187.815 ;
        RECT 90.975 187.535 91.145 188.545 ;
        RECT 90.615 187.235 90.805 187.440 ;
        RECT 91.315 187.485 91.645 188.330 ;
        RECT 92.855 187.485 93.185 188.330 ;
        RECT 93.355 187.535 93.525 188.545 ;
        RECT 93.695 187.815 94.035 188.375 ;
        RECT 94.265 188.045 94.580 188.545 ;
        RECT 94.760 188.075 95.645 188.245 ;
        RECT 91.315 187.405 91.705 187.485 ;
        RECT 91.490 187.355 91.705 187.405 ;
        RECT 89.570 186.905 90.445 187.235 ;
        RECT 90.615 186.905 91.365 187.235 ;
        RECT 89.570 186.445 89.740 186.905 ;
        RECT 90.615 186.735 90.815 186.905 ;
        RECT 91.535 186.775 91.705 187.355 ;
        RECT 91.480 186.735 91.705 186.775 ;
        RECT 88.380 186.275 88.785 186.445 ;
        RECT 88.955 186.275 89.740 186.445 ;
        RECT 90.015 185.995 90.225 186.525 ;
        RECT 90.485 186.210 90.815 186.735 ;
        RECT 91.325 186.650 91.705 186.735 ;
        RECT 92.795 187.405 93.185 187.485 ;
        RECT 93.695 187.440 94.590 187.815 ;
        RECT 92.795 187.355 93.010 187.405 ;
        RECT 92.795 186.775 92.965 187.355 ;
        RECT 93.695 187.235 93.885 187.440 ;
        RECT 94.760 187.235 94.930 188.075 ;
        RECT 95.870 188.045 96.120 188.375 ;
        RECT 93.135 186.905 93.885 187.235 ;
        RECT 94.055 186.905 94.930 187.235 ;
        RECT 92.795 186.735 93.020 186.775 ;
        RECT 93.685 186.735 93.885 186.905 ;
        RECT 92.795 186.650 93.175 186.735 ;
        RECT 90.985 185.995 91.155 186.605 ;
        RECT 91.325 186.215 91.655 186.650 ;
        RECT 92.845 186.215 93.175 186.650 ;
        RECT 93.345 185.995 93.515 186.605 ;
        RECT 93.685 186.210 94.015 186.735 ;
        RECT 94.275 185.995 94.485 186.525 ;
        RECT 94.760 186.445 94.930 186.905 ;
        RECT 95.100 186.945 95.420 187.905 ;
        RECT 95.590 187.155 95.780 187.875 ;
        RECT 95.950 186.975 96.120 188.045 ;
        RECT 96.290 187.745 96.460 188.545 ;
        RECT 96.630 188.100 97.735 188.270 ;
        RECT 96.630 187.485 96.800 188.100 ;
        RECT 97.945 187.950 98.195 188.375 ;
        RECT 98.365 188.085 98.630 188.545 ;
        RECT 96.970 187.565 97.500 187.930 ;
        RECT 97.945 187.820 98.250 187.950 ;
        RECT 96.290 187.395 96.800 187.485 ;
        RECT 96.290 187.225 97.160 187.395 ;
        RECT 96.290 187.155 96.460 187.225 ;
        RECT 96.580 186.975 96.780 187.005 ;
        RECT 95.100 186.615 95.565 186.945 ;
        RECT 95.950 186.675 96.780 186.975 ;
        RECT 95.950 186.445 96.120 186.675 ;
        RECT 94.760 186.275 95.545 186.445 ;
        RECT 95.715 186.275 96.120 186.445 ;
        RECT 96.300 185.995 96.670 186.495 ;
        RECT 96.990 186.445 97.160 187.225 ;
        RECT 97.330 186.865 97.500 187.565 ;
        RECT 97.670 187.035 97.910 187.630 ;
        RECT 97.330 186.645 97.855 186.865 ;
        RECT 98.080 186.715 98.250 187.820 ;
        RECT 98.025 186.585 98.250 186.715 ;
        RECT 98.420 186.625 98.700 187.575 ;
        RECT 98.025 186.445 98.195 186.585 ;
        RECT 96.990 186.275 97.665 186.445 ;
        RECT 97.860 186.275 98.195 186.445 ;
        RECT 98.365 185.995 98.615 186.455 ;
        RECT 98.870 186.255 99.055 188.375 ;
        RECT 99.225 188.045 99.555 188.545 ;
        RECT 99.725 187.875 99.895 188.375 ;
        RECT 99.230 187.705 99.895 187.875 ;
        RECT 99.230 186.715 99.460 187.705 ;
        RECT 99.630 186.885 99.980 187.535 ;
        RECT 100.160 187.405 100.495 188.375 ;
        RECT 100.665 187.405 100.835 188.545 ;
        RECT 101.005 188.205 103.035 188.375 ;
        RECT 100.160 186.735 100.330 187.405 ;
        RECT 101.005 187.235 101.175 188.205 ;
        RECT 100.500 186.905 100.755 187.235 ;
        RECT 100.980 186.905 101.175 187.235 ;
        RECT 101.345 187.865 102.470 188.035 ;
        RECT 100.585 186.735 100.755 186.905 ;
        RECT 101.345 186.735 101.515 187.865 ;
        RECT 99.230 186.545 99.895 186.715 ;
        RECT 99.225 185.995 99.555 186.375 ;
        RECT 99.725 186.255 99.895 186.545 ;
        RECT 100.160 186.165 100.415 186.735 ;
        RECT 100.585 186.565 101.515 186.735 ;
        RECT 101.685 187.525 102.695 187.695 ;
        RECT 101.685 186.725 101.855 187.525 ;
        RECT 101.340 186.530 101.515 186.565 ;
        RECT 100.585 185.995 100.915 186.395 ;
        RECT 101.340 186.165 101.870 186.530 ;
        RECT 102.060 186.505 102.335 187.325 ;
        RECT 102.055 186.335 102.335 186.505 ;
        RECT 102.060 186.165 102.335 186.335 ;
        RECT 102.505 186.165 102.695 187.525 ;
        RECT 102.865 187.540 103.035 188.205 ;
        RECT 103.205 187.785 103.375 188.545 ;
        RECT 103.610 187.785 104.125 188.195 ;
        RECT 102.865 187.350 103.615 187.540 ;
        RECT 103.785 186.975 104.125 187.785 ;
        RECT 104.295 187.455 106.885 188.545 ;
        RECT 102.895 186.805 104.125 186.975 ;
        RECT 102.875 185.995 103.385 186.530 ;
        RECT 103.605 186.200 103.850 186.805 ;
        RECT 104.295 186.765 105.505 187.285 ;
        RECT 105.675 186.935 106.885 187.455 ;
        RECT 107.515 187.380 107.805 188.545 ;
        RECT 107.975 187.695 108.235 188.375 ;
        RECT 108.405 187.765 108.655 188.545 ;
        RECT 108.905 187.995 109.155 188.375 ;
        RECT 109.325 188.165 109.680 188.545 ;
        RECT 110.685 188.155 111.020 188.375 ;
        RECT 110.285 187.995 110.515 188.035 ;
        RECT 108.905 187.795 110.515 187.995 ;
        RECT 108.905 187.785 109.740 187.795 ;
        RECT 110.330 187.705 110.515 187.795 ;
        RECT 104.295 185.995 106.885 186.765 ;
        RECT 107.515 185.995 107.805 186.720 ;
        RECT 107.975 186.505 108.145 187.695 ;
        RECT 109.845 187.595 110.175 187.625 ;
        RECT 108.375 187.535 110.175 187.595 ;
        RECT 110.765 187.535 111.020 188.155 ;
        RECT 111.195 188.110 116.540 188.545 ;
        RECT 108.315 187.425 111.020 187.535 ;
        RECT 108.315 187.390 108.515 187.425 ;
        RECT 108.315 186.815 108.485 187.390 ;
        RECT 109.845 187.365 111.020 187.425 ;
        RECT 108.715 186.950 109.125 187.255 ;
        RECT 109.295 186.985 109.625 187.195 ;
        RECT 108.315 186.695 108.585 186.815 ;
        RECT 108.315 186.650 109.160 186.695 ;
        RECT 108.405 186.525 109.160 186.650 ;
        RECT 109.415 186.585 109.625 186.985 ;
        RECT 109.870 186.985 110.345 187.195 ;
        RECT 110.535 186.985 111.025 187.185 ;
        RECT 109.870 186.585 110.090 186.985 ;
        RECT 107.975 186.495 108.205 186.505 ;
        RECT 107.975 186.165 108.235 186.495 ;
        RECT 108.990 186.375 109.160 186.525 ;
        RECT 108.405 185.995 108.735 186.355 ;
        RECT 108.990 186.165 110.290 186.375 ;
        RECT 110.565 185.995 111.020 186.760 ;
        RECT 112.780 186.540 113.120 187.370 ;
        RECT 114.600 186.860 114.950 188.110 ;
        RECT 116.775 187.485 117.105 188.330 ;
        RECT 117.275 187.535 117.445 188.545 ;
        RECT 117.615 187.815 117.955 188.375 ;
        RECT 118.185 188.045 118.500 188.545 ;
        RECT 118.680 188.075 119.565 188.245 ;
        RECT 116.715 187.405 117.105 187.485 ;
        RECT 117.615 187.440 118.510 187.815 ;
        RECT 116.715 187.355 116.930 187.405 ;
        RECT 116.715 186.775 116.885 187.355 ;
        RECT 117.615 187.235 117.805 187.440 ;
        RECT 118.680 187.235 118.850 188.075 ;
        RECT 119.790 188.045 120.040 188.375 ;
        RECT 117.055 186.905 117.805 187.235 ;
        RECT 117.975 186.905 118.850 187.235 ;
        RECT 116.715 186.735 116.940 186.775 ;
        RECT 117.605 186.735 117.805 186.905 ;
        RECT 116.715 186.650 117.095 186.735 ;
        RECT 111.195 185.995 116.540 186.540 ;
        RECT 116.765 186.215 117.095 186.650 ;
        RECT 117.265 185.995 117.435 186.605 ;
        RECT 117.605 186.210 117.935 186.735 ;
        RECT 118.195 185.995 118.405 186.525 ;
        RECT 118.680 186.445 118.850 186.905 ;
        RECT 119.020 186.945 119.340 187.905 ;
        RECT 119.510 187.155 119.700 187.875 ;
        RECT 119.870 186.975 120.040 188.045 ;
        RECT 120.210 187.745 120.380 188.545 ;
        RECT 120.550 188.100 121.655 188.270 ;
        RECT 120.550 187.485 120.720 188.100 ;
        RECT 121.865 187.950 122.115 188.375 ;
        RECT 122.285 188.085 122.550 188.545 ;
        RECT 120.890 187.565 121.420 187.930 ;
        RECT 121.865 187.820 122.170 187.950 ;
        RECT 120.210 187.395 120.720 187.485 ;
        RECT 120.210 187.225 121.080 187.395 ;
        RECT 120.210 187.155 120.380 187.225 ;
        RECT 120.500 186.975 120.700 187.005 ;
        RECT 119.020 186.615 119.485 186.945 ;
        RECT 119.870 186.675 120.700 186.975 ;
        RECT 119.870 186.445 120.040 186.675 ;
        RECT 118.680 186.275 119.465 186.445 ;
        RECT 119.635 186.275 120.040 186.445 ;
        RECT 120.220 185.995 120.590 186.495 ;
        RECT 120.910 186.445 121.080 187.225 ;
        RECT 121.250 186.865 121.420 187.565 ;
        RECT 121.590 187.035 121.830 187.630 ;
        RECT 121.250 186.645 121.775 186.865 ;
        RECT 122.000 186.715 122.170 187.820 ;
        RECT 121.945 186.585 122.170 186.715 ;
        RECT 122.340 186.625 122.620 187.575 ;
        RECT 121.945 186.445 122.115 186.585 ;
        RECT 120.910 186.275 121.585 186.445 ;
        RECT 121.780 186.275 122.115 186.445 ;
        RECT 122.285 185.995 122.535 186.455 ;
        RECT 122.790 186.255 122.975 188.375 ;
        RECT 123.145 188.045 123.475 188.545 ;
        RECT 123.645 187.875 123.815 188.375 ;
        RECT 123.150 187.705 123.815 187.875 ;
        RECT 123.150 186.715 123.380 187.705 ;
        RECT 124.075 187.695 124.335 188.375 ;
        RECT 124.505 187.765 124.755 188.545 ;
        RECT 125.005 187.995 125.255 188.375 ;
        RECT 125.425 188.165 125.780 188.545 ;
        RECT 126.785 188.155 127.120 188.375 ;
        RECT 126.385 187.995 126.615 188.035 ;
        RECT 125.005 187.795 126.615 187.995 ;
        RECT 125.005 187.785 125.840 187.795 ;
        RECT 126.430 187.705 126.615 187.795 ;
        RECT 123.550 186.885 123.900 187.535 ;
        RECT 123.150 186.545 123.815 186.715 ;
        RECT 123.145 185.995 123.475 186.375 ;
        RECT 123.645 186.255 123.815 186.545 ;
        RECT 124.075 186.495 124.245 187.695 ;
        RECT 125.945 187.595 126.275 187.625 ;
        RECT 124.475 187.535 126.275 187.595 ;
        RECT 126.865 187.535 127.120 188.155 ;
        RECT 124.415 187.425 127.120 187.535 ;
        RECT 124.415 187.390 124.615 187.425 ;
        RECT 124.415 186.815 124.585 187.390 ;
        RECT 125.945 187.365 127.120 187.425 ;
        RECT 127.300 187.405 127.575 188.375 ;
        RECT 127.785 187.745 128.065 188.545 ;
        RECT 128.235 188.035 129.425 188.325 ;
        RECT 129.685 188.205 130.845 188.375 ;
        RECT 128.235 187.695 129.405 187.865 ;
        RECT 129.685 187.705 129.855 188.205 ;
        RECT 128.235 187.575 128.405 187.695 ;
        RECT 127.745 187.405 128.405 187.575 ;
        RECT 124.815 186.950 125.225 187.255 ;
        RECT 125.395 186.985 125.725 187.195 ;
        RECT 124.415 186.695 124.685 186.815 ;
        RECT 124.415 186.650 125.260 186.695 ;
        RECT 124.505 186.525 125.260 186.650 ;
        RECT 125.515 186.585 125.725 186.985 ;
        RECT 125.970 186.985 126.445 187.195 ;
        RECT 126.635 186.985 127.125 187.185 ;
        RECT 125.970 186.585 126.190 186.985 ;
        RECT 124.075 186.165 124.335 186.495 ;
        RECT 125.090 186.375 125.260 186.525 ;
        RECT 124.505 185.995 124.835 186.355 ;
        RECT 125.090 186.165 126.390 186.375 ;
        RECT 126.665 185.995 127.120 186.760 ;
        RECT 127.300 186.670 127.470 187.405 ;
        RECT 127.745 187.235 127.915 187.405 ;
        RECT 128.715 187.235 128.910 187.525 ;
        RECT 129.080 187.405 129.405 187.695 ;
        RECT 130.115 187.575 130.285 188.035 ;
        RECT 130.515 187.955 130.845 188.205 ;
        RECT 131.070 188.125 131.400 188.545 ;
        RECT 131.655 187.955 131.940 188.375 ;
        RECT 130.515 187.785 131.940 187.955 ;
        RECT 132.185 187.745 132.515 188.545 ;
        RECT 132.765 187.825 133.100 188.335 ;
        RECT 129.660 187.235 129.865 187.525 ;
        RECT 130.115 187.405 132.485 187.575 ;
        RECT 132.315 187.235 132.485 187.405 ;
        RECT 127.640 186.905 127.915 187.235 ;
        RECT 128.085 186.905 128.910 187.235 ;
        RECT 129.080 186.905 129.425 187.235 ;
        RECT 129.660 187.185 130.010 187.235 ;
        RECT 129.655 187.015 130.010 187.185 ;
        RECT 129.660 186.905 130.010 187.015 ;
        RECT 127.745 186.735 127.915 186.905 ;
        RECT 127.300 186.325 127.575 186.670 ;
        RECT 127.745 186.565 129.410 186.735 ;
        RECT 127.765 185.995 128.145 186.395 ;
        RECT 128.315 186.215 128.485 186.565 ;
        RECT 128.655 185.995 128.985 186.395 ;
        RECT 129.155 186.215 129.410 186.565 ;
        RECT 129.605 185.995 129.935 186.715 ;
        RECT 130.320 186.570 130.740 187.235 ;
        RECT 130.910 186.845 131.200 187.235 ;
        RECT 131.390 186.845 131.660 187.235 ;
        RECT 131.870 187.185 132.120 187.235 ;
        RECT 131.870 187.015 132.125 187.185 ;
        RECT 131.870 186.905 132.120 187.015 ;
        RECT 132.315 186.905 132.620 187.235 ;
        RECT 130.910 186.675 131.205 186.845 ;
        RECT 131.390 186.675 131.665 186.845 ;
        RECT 132.315 186.735 132.485 186.905 ;
        RECT 130.910 186.575 131.200 186.675 ;
        RECT 131.390 186.575 131.660 186.675 ;
        RECT 131.925 186.565 132.485 186.735 ;
        RECT 131.925 186.395 132.095 186.565 ;
        RECT 132.845 186.470 133.100 187.825 ;
        RECT 133.275 187.380 133.565 188.545 ;
        RECT 133.825 187.875 133.995 188.375 ;
        RECT 134.165 188.045 134.495 188.545 ;
        RECT 133.825 187.705 134.490 187.875 ;
        RECT 133.740 186.885 134.090 187.535 ;
        RECT 130.480 186.225 132.095 186.395 ;
        RECT 132.265 185.995 132.595 186.395 ;
        RECT 132.765 186.210 133.100 186.470 ;
        RECT 133.275 185.995 133.565 186.720 ;
        RECT 134.260 186.715 134.490 187.705 ;
        RECT 133.825 186.545 134.490 186.715 ;
        RECT 133.825 186.255 133.995 186.545 ;
        RECT 134.165 185.995 134.495 186.375 ;
        RECT 134.665 186.255 134.850 188.375 ;
        RECT 135.090 188.085 135.355 188.545 ;
        RECT 135.525 187.950 135.775 188.375 ;
        RECT 135.985 188.100 137.090 188.270 ;
        RECT 135.470 187.820 135.775 187.950 ;
        RECT 135.020 186.625 135.300 187.575 ;
        RECT 135.470 186.715 135.640 187.820 ;
        RECT 135.810 187.035 136.050 187.630 ;
        RECT 136.220 187.565 136.750 187.930 ;
        RECT 136.220 186.865 136.390 187.565 ;
        RECT 136.920 187.485 137.090 188.100 ;
        RECT 137.260 187.745 137.430 188.545 ;
        RECT 137.600 188.045 137.850 188.375 ;
        RECT 138.075 188.075 138.960 188.245 ;
        RECT 136.920 187.395 137.430 187.485 ;
        RECT 135.470 186.585 135.695 186.715 ;
        RECT 135.865 186.645 136.390 186.865 ;
        RECT 136.560 187.225 137.430 187.395 ;
        RECT 135.105 185.995 135.355 186.455 ;
        RECT 135.525 186.445 135.695 186.585 ;
        RECT 136.560 186.445 136.730 187.225 ;
        RECT 137.260 187.155 137.430 187.225 ;
        RECT 136.940 186.975 137.140 187.005 ;
        RECT 137.600 186.975 137.770 188.045 ;
        RECT 137.940 187.155 138.130 187.875 ;
        RECT 136.940 186.675 137.770 186.975 ;
        RECT 138.300 186.945 138.620 187.905 ;
        RECT 135.525 186.275 135.860 186.445 ;
        RECT 136.055 186.275 136.730 186.445 ;
        RECT 137.050 185.995 137.420 186.495 ;
        RECT 137.600 186.445 137.770 186.675 ;
        RECT 138.155 186.615 138.620 186.945 ;
        RECT 138.790 187.235 138.960 188.075 ;
        RECT 139.140 188.045 139.455 188.545 ;
        RECT 139.685 187.815 140.025 188.375 ;
        RECT 139.130 187.440 140.025 187.815 ;
        RECT 140.195 187.535 140.365 188.545 ;
        RECT 139.835 187.235 140.025 187.440 ;
        RECT 140.535 187.485 140.865 188.330 ;
        RECT 141.095 187.695 141.355 188.375 ;
        RECT 141.525 187.765 141.775 188.545 ;
        RECT 142.025 187.995 142.275 188.375 ;
        RECT 142.445 188.165 142.800 188.545 ;
        RECT 143.805 188.155 144.140 188.375 ;
        RECT 143.405 187.995 143.635 188.035 ;
        RECT 142.025 187.795 143.635 187.995 ;
        RECT 142.025 187.785 142.860 187.795 ;
        RECT 143.450 187.705 143.635 187.795 ;
        RECT 140.535 187.405 140.925 187.485 ;
        RECT 140.710 187.355 140.925 187.405 ;
        RECT 138.790 186.905 139.665 187.235 ;
        RECT 139.835 186.905 140.585 187.235 ;
        RECT 138.790 186.445 138.960 186.905 ;
        RECT 139.835 186.735 140.035 186.905 ;
        RECT 140.755 186.775 140.925 187.355 ;
        RECT 140.700 186.735 140.925 186.775 ;
        RECT 137.600 186.275 138.005 186.445 ;
        RECT 138.175 186.275 138.960 186.445 ;
        RECT 139.235 185.995 139.445 186.525 ;
        RECT 139.705 186.210 140.035 186.735 ;
        RECT 140.545 186.650 140.925 186.735 ;
        RECT 140.205 185.995 140.375 186.605 ;
        RECT 140.545 186.215 140.875 186.650 ;
        RECT 141.095 186.495 141.265 187.695 ;
        RECT 142.965 187.595 143.295 187.625 ;
        RECT 141.495 187.535 143.295 187.595 ;
        RECT 143.885 187.535 144.140 188.155 ;
        RECT 141.435 187.425 144.140 187.535 ;
        RECT 144.315 187.455 145.525 188.545 ;
        RECT 141.435 187.390 141.635 187.425 ;
        RECT 141.435 186.815 141.605 187.390 ;
        RECT 142.965 187.365 144.140 187.425 ;
        RECT 141.835 186.950 142.245 187.255 ;
        RECT 142.415 186.985 142.745 187.195 ;
        RECT 141.435 186.695 141.705 186.815 ;
        RECT 141.435 186.650 142.280 186.695 ;
        RECT 141.525 186.525 142.280 186.650 ;
        RECT 142.535 186.585 142.745 186.985 ;
        RECT 142.990 186.985 143.465 187.195 ;
        RECT 143.655 186.985 144.145 187.185 ;
        RECT 142.990 186.585 143.210 186.985 ;
        RECT 141.095 186.165 141.355 186.495 ;
        RECT 142.110 186.375 142.280 186.525 ;
        RECT 141.525 185.995 141.855 186.355 ;
        RECT 142.110 186.165 143.410 186.375 ;
        RECT 143.685 185.995 144.140 186.760 ;
        RECT 144.315 186.745 144.835 187.285 ;
        RECT 145.005 186.915 145.525 187.455 ;
        RECT 145.695 187.455 146.905 188.545 ;
        RECT 145.695 186.915 146.215 187.455 ;
        RECT 146.385 186.745 146.905 187.285 ;
        RECT 144.315 185.995 145.525 186.745 ;
        RECT 145.695 185.995 146.905 186.745 ;
        RECT 17.270 185.825 146.990 185.995 ;
        RECT 17.355 185.075 18.565 185.825 ;
        RECT 19.745 185.275 19.915 185.565 ;
        RECT 20.085 185.445 20.415 185.825 ;
        RECT 19.745 185.105 20.410 185.275 ;
        RECT 17.355 184.535 17.875 185.075 ;
        RECT 18.045 184.365 18.565 184.905 ;
        RECT 17.355 183.275 18.565 184.365 ;
        RECT 19.660 184.285 20.010 184.935 ;
        RECT 20.180 184.115 20.410 185.105 ;
        RECT 19.745 183.945 20.410 184.115 ;
        RECT 19.745 183.445 19.915 183.945 ;
        RECT 20.085 183.275 20.415 183.775 ;
        RECT 20.585 183.445 20.770 185.565 ;
        RECT 21.025 185.365 21.275 185.825 ;
        RECT 21.445 185.375 21.780 185.545 ;
        RECT 21.975 185.375 22.650 185.545 ;
        RECT 21.445 185.235 21.615 185.375 ;
        RECT 20.940 184.245 21.220 185.195 ;
        RECT 21.390 185.105 21.615 185.235 ;
        RECT 21.390 184.000 21.560 185.105 ;
        RECT 21.785 184.955 22.310 185.175 ;
        RECT 21.730 184.190 21.970 184.785 ;
        RECT 22.140 184.255 22.310 184.955 ;
        RECT 22.480 184.595 22.650 185.375 ;
        RECT 22.970 185.325 23.340 185.825 ;
        RECT 23.520 185.375 23.925 185.545 ;
        RECT 24.095 185.375 24.880 185.545 ;
        RECT 23.520 185.145 23.690 185.375 ;
        RECT 22.860 184.845 23.690 185.145 ;
        RECT 24.075 184.875 24.540 185.205 ;
        RECT 22.860 184.815 23.060 184.845 ;
        RECT 23.180 184.595 23.350 184.665 ;
        RECT 22.480 184.425 23.350 184.595 ;
        RECT 22.840 184.335 23.350 184.425 ;
        RECT 21.390 183.870 21.695 184.000 ;
        RECT 22.140 183.890 22.670 184.255 ;
        RECT 21.010 183.275 21.275 183.735 ;
        RECT 21.445 183.445 21.695 183.870 ;
        RECT 22.840 183.720 23.010 184.335 ;
        RECT 21.905 183.550 23.010 183.720 ;
        RECT 23.180 183.275 23.350 184.075 ;
        RECT 23.520 183.775 23.690 184.845 ;
        RECT 23.860 183.945 24.050 184.665 ;
        RECT 24.220 183.915 24.540 184.875 ;
        RECT 24.710 184.915 24.880 185.375 ;
        RECT 25.155 185.295 25.365 185.825 ;
        RECT 25.625 185.085 25.955 185.610 ;
        RECT 26.125 185.215 26.295 185.825 ;
        RECT 26.465 185.170 26.795 185.605 ;
        RECT 27.015 185.445 27.905 185.615 ;
        RECT 26.465 185.085 26.845 185.170 ;
        RECT 25.755 184.915 25.955 185.085 ;
        RECT 26.620 185.045 26.845 185.085 ;
        RECT 24.710 184.585 25.585 184.915 ;
        RECT 25.755 184.585 26.505 184.915 ;
        RECT 23.520 183.445 23.770 183.775 ;
        RECT 24.710 183.745 24.880 184.585 ;
        RECT 25.755 184.380 25.945 184.585 ;
        RECT 26.675 184.465 26.845 185.045 ;
        RECT 27.015 184.890 27.565 185.275 ;
        RECT 27.735 184.720 27.905 185.445 ;
        RECT 26.630 184.415 26.845 184.465 ;
        RECT 25.050 184.005 25.945 184.380 ;
        RECT 26.455 184.335 26.845 184.415 ;
        RECT 27.015 184.650 27.905 184.720 ;
        RECT 28.075 185.120 28.295 185.605 ;
        RECT 28.465 185.285 28.715 185.825 ;
        RECT 28.885 185.175 29.145 185.655 ;
        RECT 28.075 184.695 28.405 185.120 ;
        RECT 27.015 184.625 27.910 184.650 ;
        RECT 27.015 184.610 27.920 184.625 ;
        RECT 27.015 184.595 27.925 184.610 ;
        RECT 27.015 184.590 27.935 184.595 ;
        RECT 27.015 184.580 27.940 184.590 ;
        RECT 27.015 184.570 27.945 184.580 ;
        RECT 27.015 184.565 27.955 184.570 ;
        RECT 27.015 184.555 27.965 184.565 ;
        RECT 27.015 184.550 27.975 184.555 ;
        RECT 23.995 183.575 24.880 183.745 ;
        RECT 25.060 183.275 25.375 183.775 ;
        RECT 25.605 183.445 25.945 184.005 ;
        RECT 26.115 183.275 26.285 184.285 ;
        RECT 26.455 183.490 26.785 184.335 ;
        RECT 27.015 184.100 27.275 184.550 ;
        RECT 27.640 184.545 27.975 184.550 ;
        RECT 27.640 184.540 27.990 184.545 ;
        RECT 27.640 184.530 28.005 184.540 ;
        RECT 27.640 184.525 28.030 184.530 ;
        RECT 28.575 184.525 28.805 184.920 ;
        RECT 27.640 184.520 28.805 184.525 ;
        RECT 27.670 184.485 28.805 184.520 ;
        RECT 27.705 184.460 28.805 184.485 ;
        RECT 27.735 184.430 28.805 184.460 ;
        RECT 27.755 184.400 28.805 184.430 ;
        RECT 27.775 184.370 28.805 184.400 ;
        RECT 27.845 184.360 28.805 184.370 ;
        RECT 27.870 184.350 28.805 184.360 ;
        RECT 27.890 184.335 28.805 184.350 ;
        RECT 27.910 184.320 28.805 184.335 ;
        RECT 27.915 184.310 28.700 184.320 ;
        RECT 27.930 184.275 28.700 184.310 ;
        RECT 27.445 183.955 27.775 184.200 ;
        RECT 27.945 184.025 28.700 184.275 ;
        RECT 28.975 184.145 29.145 185.175 ;
        RECT 27.445 183.930 27.630 183.955 ;
        RECT 27.015 183.830 27.630 183.930 ;
        RECT 27.015 183.275 27.620 183.830 ;
        RECT 27.795 183.445 28.275 183.785 ;
        RECT 28.445 183.275 28.700 183.820 ;
        RECT 28.870 183.445 29.145 184.145 ;
        RECT 29.315 185.175 29.575 185.655 ;
        RECT 29.745 185.285 29.995 185.825 ;
        RECT 29.315 184.145 29.485 185.175 ;
        RECT 30.165 185.120 30.385 185.605 ;
        RECT 29.655 184.525 29.885 184.920 ;
        RECT 30.055 184.695 30.385 185.120 ;
        RECT 30.555 185.445 31.445 185.615 ;
        RECT 30.555 184.720 30.725 185.445 ;
        RECT 30.895 184.890 31.445 185.275 ;
        RECT 31.655 185.005 31.885 185.825 ;
        RECT 32.055 185.025 32.385 185.655 ;
        RECT 30.555 184.650 31.445 184.720 ;
        RECT 30.550 184.625 31.445 184.650 ;
        RECT 30.540 184.610 31.445 184.625 ;
        RECT 30.535 184.595 31.445 184.610 ;
        RECT 30.525 184.590 31.445 184.595 ;
        RECT 30.520 184.580 31.445 184.590 ;
        RECT 31.635 184.585 31.965 184.835 ;
        RECT 30.515 184.570 31.445 184.580 ;
        RECT 30.505 184.565 31.445 184.570 ;
        RECT 30.495 184.555 31.445 184.565 ;
        RECT 30.485 184.550 31.445 184.555 ;
        RECT 30.485 184.545 30.820 184.550 ;
        RECT 30.470 184.540 30.820 184.545 ;
        RECT 30.455 184.530 30.820 184.540 ;
        RECT 30.430 184.525 30.820 184.530 ;
        RECT 29.655 184.520 30.820 184.525 ;
        RECT 29.655 184.485 30.790 184.520 ;
        RECT 29.655 184.460 30.755 184.485 ;
        RECT 29.655 184.430 30.725 184.460 ;
        RECT 29.655 184.400 30.705 184.430 ;
        RECT 29.655 184.370 30.685 184.400 ;
        RECT 29.655 184.360 30.615 184.370 ;
        RECT 29.655 184.350 30.590 184.360 ;
        RECT 29.655 184.335 30.570 184.350 ;
        RECT 29.655 184.320 30.550 184.335 ;
        RECT 29.760 184.310 30.545 184.320 ;
        RECT 29.760 184.275 30.530 184.310 ;
        RECT 29.315 183.445 29.590 184.145 ;
        RECT 29.760 184.025 30.515 184.275 ;
        RECT 30.685 183.955 31.015 184.200 ;
        RECT 31.185 184.100 31.445 184.550 ;
        RECT 32.135 184.425 32.385 185.025 ;
        RECT 32.555 185.005 32.765 185.825 ;
        RECT 32.995 185.055 36.505 185.825 ;
        RECT 37.295 185.265 37.625 185.655 ;
        RECT 37.795 185.435 38.980 185.605 ;
        RECT 39.240 185.355 39.410 185.825 ;
        RECT 37.295 185.085 37.805 185.265 ;
        RECT 32.995 184.535 34.645 185.055 ;
        RECT 30.830 183.930 31.015 183.955 ;
        RECT 30.830 183.830 31.445 183.930 ;
        RECT 29.760 183.275 30.015 183.820 ;
        RECT 30.185 183.445 30.665 183.785 ;
        RECT 30.840 183.275 31.445 183.830 ;
        RECT 31.655 183.275 31.885 184.415 ;
        RECT 32.055 183.445 32.385 184.425 ;
        RECT 32.555 183.275 32.765 184.415 ;
        RECT 34.815 184.365 36.505 184.885 ;
        RECT 37.135 184.625 37.465 184.915 ;
        RECT 37.635 184.455 37.805 185.085 ;
        RECT 38.210 185.175 38.595 185.265 ;
        RECT 39.580 185.175 39.910 185.640 ;
        RECT 38.210 185.005 39.910 185.175 ;
        RECT 40.080 185.005 40.250 185.825 ;
        RECT 40.420 185.005 41.105 185.645 ;
        RECT 41.295 185.015 41.535 185.825 ;
        RECT 41.705 185.015 42.035 185.655 ;
        RECT 42.205 185.015 42.475 185.825 ;
        RECT 43.115 185.100 43.405 185.825 ;
        RECT 43.575 185.085 44.015 185.645 ;
        RECT 44.185 185.085 44.635 185.825 ;
        RECT 44.805 185.255 44.975 185.655 ;
        RECT 45.145 185.425 45.565 185.825 ;
        RECT 45.735 185.255 45.965 185.655 ;
        RECT 44.805 185.085 45.965 185.255 ;
        RECT 46.135 185.085 46.625 185.655 ;
        RECT 46.795 185.280 52.140 185.825 ;
        RECT 52.315 185.280 57.660 185.825 ;
        RECT 37.975 184.625 38.305 184.835 ;
        RECT 38.485 184.585 38.865 184.835 ;
        RECT 39.055 184.805 39.540 184.835 ;
        RECT 39.035 184.635 39.540 184.805 ;
        RECT 32.995 183.275 36.505 184.365 ;
        RECT 37.290 184.285 38.375 184.455 ;
        RECT 37.290 183.445 37.590 184.285 ;
        RECT 37.785 183.275 38.035 184.115 ;
        RECT 38.205 184.035 38.375 184.285 ;
        RECT 38.545 184.205 38.865 184.585 ;
        RECT 39.055 184.625 39.540 184.635 ;
        RECT 39.730 184.625 40.180 184.835 ;
        RECT 40.350 184.625 40.685 184.835 ;
        RECT 39.055 184.205 39.430 184.625 ;
        RECT 40.350 184.455 40.520 184.625 ;
        RECT 39.600 184.285 40.520 184.455 ;
        RECT 39.600 184.035 39.770 184.285 ;
        RECT 38.205 183.865 39.770 184.035 ;
        RECT 38.625 183.445 39.430 183.865 ;
        RECT 39.940 183.275 40.270 184.115 ;
        RECT 40.855 184.035 41.105 185.005 ;
        RECT 41.275 184.585 41.625 184.835 ;
        RECT 41.795 184.415 41.965 185.015 ;
        RECT 42.135 184.585 42.485 184.835 ;
        RECT 40.440 183.445 41.105 184.035 ;
        RECT 41.285 184.245 41.965 184.415 ;
        RECT 41.285 183.460 41.615 184.245 ;
        RECT 42.145 183.275 42.475 184.415 ;
        RECT 43.115 183.275 43.405 184.440 ;
        RECT 43.575 184.075 43.885 185.085 ;
        RECT 44.055 184.465 44.225 184.915 ;
        RECT 44.395 184.635 44.785 184.915 ;
        RECT 44.970 184.585 45.215 184.915 ;
        RECT 44.055 184.295 44.845 184.465 ;
        RECT 43.575 183.445 44.015 184.075 ;
        RECT 44.190 183.275 44.505 184.125 ;
        RECT 44.675 183.615 44.845 184.295 ;
        RECT 45.015 183.785 45.215 184.585 ;
        RECT 45.415 183.785 45.665 184.915 ;
        RECT 45.880 184.585 46.285 184.915 ;
        RECT 46.455 184.415 46.625 185.085 ;
        RECT 48.380 184.450 48.720 185.280 ;
        RECT 45.855 184.245 46.625 184.415 ;
        RECT 45.855 183.615 46.105 184.245 ;
        RECT 44.675 183.445 46.105 183.615 ;
        RECT 46.285 183.275 46.615 184.075 ;
        RECT 50.200 183.710 50.550 184.960 ;
        RECT 53.900 184.450 54.240 185.280 ;
        RECT 57.835 185.055 60.425 185.825 ;
        RECT 55.720 183.710 56.070 184.960 ;
        RECT 57.835 184.535 59.045 185.055 ;
        RECT 61.075 185.015 61.315 185.825 ;
        RECT 61.485 185.015 61.815 185.655 ;
        RECT 61.985 185.015 62.255 185.825 ;
        RECT 59.215 184.365 60.425 184.885 ;
        RECT 61.055 184.585 61.405 184.835 ;
        RECT 61.575 184.415 61.745 185.015 ;
        RECT 61.915 184.585 62.265 184.835 ;
        RECT 46.795 183.275 52.140 183.710 ;
        RECT 52.315 183.275 57.660 183.710 ;
        RECT 57.835 183.275 60.425 184.365 ;
        RECT 61.065 184.245 61.745 184.415 ;
        RECT 61.065 183.460 61.395 184.245 ;
        RECT 61.925 183.275 62.255 184.415 ;
        RECT 62.900 184.225 63.235 185.645 ;
        RECT 63.415 185.455 64.160 185.825 ;
        RECT 64.725 185.285 64.980 185.645 ;
        RECT 65.160 185.455 65.490 185.825 ;
        RECT 65.670 185.285 65.895 185.645 ;
        RECT 63.410 185.095 65.895 185.285 ;
        RECT 63.410 184.405 63.635 185.095 ;
        RECT 66.115 185.055 68.705 185.825 ;
        RECT 68.875 185.100 69.165 185.825 ;
        RECT 69.335 185.055 72.845 185.825 ;
        RECT 73.015 185.075 74.225 185.825 ;
        RECT 74.510 185.195 74.795 185.655 ;
        RECT 74.965 185.365 75.235 185.825 ;
        RECT 63.835 184.585 64.115 184.915 ;
        RECT 64.295 184.585 64.870 184.915 ;
        RECT 65.050 184.585 65.485 184.915 ;
        RECT 65.665 184.585 65.935 184.915 ;
        RECT 66.115 184.535 67.325 185.055 ;
        RECT 63.410 184.225 65.905 184.405 ;
        RECT 67.495 184.365 68.705 184.885 ;
        RECT 69.335 184.535 70.985 185.055 ;
        RECT 62.900 183.455 63.165 184.225 ;
        RECT 63.335 183.275 63.665 183.995 ;
        RECT 63.855 183.815 65.045 184.045 ;
        RECT 63.855 183.455 64.115 183.815 ;
        RECT 64.285 183.275 64.615 183.645 ;
        RECT 64.785 183.455 65.045 183.815 ;
        RECT 65.615 183.455 65.905 184.225 ;
        RECT 66.115 183.275 68.705 184.365 ;
        RECT 68.875 183.275 69.165 184.440 ;
        RECT 71.155 184.365 72.845 184.885 ;
        RECT 73.015 184.535 73.535 185.075 ;
        RECT 74.510 185.025 75.465 185.195 ;
        RECT 73.705 184.365 74.225 184.905 ;
        RECT 69.335 183.275 72.845 184.365 ;
        RECT 73.015 183.275 74.225 184.365 ;
        RECT 74.395 184.295 75.085 184.855 ;
        RECT 75.255 184.125 75.465 185.025 ;
        RECT 74.510 183.905 75.465 184.125 ;
        RECT 75.635 184.855 76.035 185.655 ;
        RECT 76.225 185.195 76.505 185.655 ;
        RECT 77.025 185.365 77.350 185.825 ;
        RECT 76.225 185.025 77.350 185.195 ;
        RECT 77.520 185.085 77.905 185.655 ;
        RECT 76.900 184.915 77.350 185.025 ;
        RECT 75.635 184.295 76.730 184.855 ;
        RECT 76.900 184.585 77.455 184.915 ;
        RECT 74.510 183.445 74.795 183.905 ;
        RECT 74.965 183.275 75.235 183.735 ;
        RECT 75.635 183.445 76.035 184.295 ;
        RECT 76.900 184.125 77.350 184.585 ;
        RECT 77.625 184.415 77.905 185.085 ;
        RECT 78.095 185.015 78.335 185.825 ;
        RECT 78.505 185.015 78.835 185.655 ;
        RECT 79.005 185.015 79.275 185.825 ;
        RECT 79.455 185.280 84.800 185.825 ;
        RECT 78.075 184.585 78.425 184.835 ;
        RECT 78.595 184.415 78.765 185.015 ;
        RECT 78.935 184.585 79.285 184.835 ;
        RECT 81.040 184.450 81.380 185.280 ;
        RECT 84.975 185.055 86.645 185.825 ;
        RECT 87.365 185.275 87.535 185.565 ;
        RECT 87.705 185.445 88.035 185.825 ;
        RECT 87.365 185.105 88.030 185.275 ;
        RECT 76.225 183.905 77.350 184.125 ;
        RECT 76.225 183.445 76.505 183.905 ;
        RECT 77.025 183.275 77.350 183.735 ;
        RECT 77.520 183.445 77.905 184.415 ;
        RECT 78.085 184.245 78.765 184.415 ;
        RECT 78.085 183.460 78.415 184.245 ;
        RECT 78.945 183.275 79.275 184.415 ;
        RECT 82.860 183.710 83.210 184.960 ;
        RECT 84.975 184.535 85.725 185.055 ;
        RECT 85.895 184.365 86.645 184.885 ;
        RECT 79.455 183.275 84.800 183.710 ;
        RECT 84.975 183.275 86.645 184.365 ;
        RECT 87.280 184.285 87.630 184.935 ;
        RECT 87.800 184.115 88.030 185.105 ;
        RECT 87.365 183.945 88.030 184.115 ;
        RECT 87.365 183.445 87.535 183.945 ;
        RECT 87.705 183.275 88.035 183.775 ;
        RECT 88.205 183.445 88.390 185.565 ;
        RECT 88.645 185.365 88.895 185.825 ;
        RECT 89.065 185.375 89.400 185.545 ;
        RECT 89.595 185.375 90.270 185.545 ;
        RECT 89.065 185.235 89.235 185.375 ;
        RECT 88.560 184.245 88.840 185.195 ;
        RECT 89.010 185.105 89.235 185.235 ;
        RECT 89.010 184.000 89.180 185.105 ;
        RECT 89.405 184.955 89.930 185.175 ;
        RECT 89.350 184.190 89.590 184.785 ;
        RECT 89.760 184.255 89.930 184.955 ;
        RECT 90.100 184.595 90.270 185.375 ;
        RECT 90.590 185.325 90.960 185.825 ;
        RECT 91.140 185.375 91.545 185.545 ;
        RECT 91.715 185.375 92.500 185.545 ;
        RECT 91.140 185.145 91.310 185.375 ;
        RECT 90.480 184.845 91.310 185.145 ;
        RECT 91.695 184.875 92.160 185.205 ;
        RECT 90.480 184.815 90.680 184.845 ;
        RECT 90.800 184.595 90.970 184.665 ;
        RECT 90.100 184.425 90.970 184.595 ;
        RECT 90.460 184.335 90.970 184.425 ;
        RECT 89.010 183.870 89.315 184.000 ;
        RECT 89.760 183.890 90.290 184.255 ;
        RECT 88.630 183.275 88.895 183.735 ;
        RECT 89.065 183.445 89.315 183.870 ;
        RECT 90.460 183.720 90.630 184.335 ;
        RECT 89.525 183.550 90.630 183.720 ;
        RECT 90.800 183.275 90.970 184.075 ;
        RECT 91.140 183.775 91.310 184.845 ;
        RECT 91.480 183.945 91.670 184.665 ;
        RECT 91.840 183.915 92.160 184.875 ;
        RECT 92.330 184.915 92.500 185.375 ;
        RECT 92.775 185.295 92.985 185.825 ;
        RECT 93.245 185.085 93.575 185.610 ;
        RECT 93.745 185.215 93.915 185.825 ;
        RECT 94.085 185.170 94.415 185.605 ;
        RECT 94.085 185.085 94.465 185.170 ;
        RECT 94.635 185.100 94.925 185.825 ;
        RECT 93.375 184.915 93.575 185.085 ;
        RECT 94.240 185.045 94.465 185.085 ;
        RECT 92.330 184.585 93.205 184.915 ;
        RECT 93.375 184.585 94.125 184.915 ;
        RECT 91.140 183.445 91.390 183.775 ;
        RECT 92.330 183.745 92.500 184.585 ;
        RECT 93.375 184.380 93.565 184.585 ;
        RECT 94.295 184.465 94.465 185.045 ;
        RECT 94.250 184.415 94.465 184.465 ;
        RECT 95.095 185.085 95.480 185.655 ;
        RECT 95.650 185.365 95.975 185.825 ;
        RECT 96.495 185.195 96.775 185.655 ;
        RECT 92.670 184.005 93.565 184.380 ;
        RECT 94.075 184.335 94.465 184.415 ;
        RECT 91.615 183.575 92.500 183.745 ;
        RECT 92.680 183.275 92.995 183.775 ;
        RECT 93.225 183.445 93.565 184.005 ;
        RECT 93.735 183.275 93.905 184.285 ;
        RECT 94.075 183.490 94.405 184.335 ;
        RECT 94.635 183.275 94.925 184.440 ;
        RECT 95.095 184.415 95.375 185.085 ;
        RECT 95.650 185.025 96.775 185.195 ;
        RECT 95.650 184.915 96.100 185.025 ;
        RECT 95.545 184.585 96.100 184.915 ;
        RECT 96.965 184.855 97.365 185.655 ;
        RECT 97.765 185.365 98.035 185.825 ;
        RECT 98.205 185.195 98.490 185.655 ;
        RECT 95.095 183.445 95.480 184.415 ;
        RECT 95.650 184.125 96.100 184.585 ;
        RECT 96.270 184.295 97.365 184.855 ;
        RECT 95.650 183.905 96.775 184.125 ;
        RECT 95.650 183.275 95.975 183.735 ;
        RECT 96.495 183.445 96.775 183.905 ;
        RECT 96.965 183.445 97.365 184.295 ;
        RECT 97.535 185.025 98.490 185.195 ;
        RECT 98.775 185.085 99.160 185.655 ;
        RECT 99.330 185.365 99.655 185.825 ;
        RECT 100.175 185.195 100.455 185.655 ;
        RECT 97.535 184.125 97.745 185.025 ;
        RECT 97.915 184.295 98.605 184.855 ;
        RECT 98.775 184.415 99.055 185.085 ;
        RECT 99.330 185.025 100.455 185.195 ;
        RECT 99.330 184.915 99.780 185.025 ;
        RECT 99.225 184.585 99.780 184.915 ;
        RECT 100.645 184.855 101.045 185.655 ;
        RECT 101.445 185.365 101.715 185.825 ;
        RECT 101.885 185.195 102.170 185.655 ;
        RECT 97.535 183.905 98.490 184.125 ;
        RECT 97.765 183.275 98.035 183.735 ;
        RECT 98.205 183.445 98.490 183.905 ;
        RECT 98.775 183.445 99.160 184.415 ;
        RECT 99.330 184.125 99.780 184.585 ;
        RECT 99.950 184.295 101.045 184.855 ;
        RECT 99.330 183.905 100.455 184.125 ;
        RECT 99.330 183.275 99.655 183.735 ;
        RECT 100.175 183.445 100.455 183.905 ;
        RECT 100.645 183.445 101.045 184.295 ;
        RECT 101.215 185.025 102.170 185.195 ;
        RECT 102.455 185.085 102.840 185.655 ;
        RECT 103.010 185.365 103.335 185.825 ;
        RECT 103.855 185.195 104.135 185.655 ;
        RECT 101.215 184.125 101.425 185.025 ;
        RECT 101.595 184.295 102.285 184.855 ;
        RECT 102.455 184.415 102.735 185.085 ;
        RECT 103.010 185.025 104.135 185.195 ;
        RECT 103.010 184.915 103.460 185.025 ;
        RECT 102.905 184.585 103.460 184.915 ;
        RECT 104.325 184.855 104.725 185.655 ;
        RECT 105.125 185.365 105.395 185.825 ;
        RECT 105.565 185.195 105.850 185.655 ;
        RECT 106.615 185.355 106.910 185.825 ;
        RECT 101.215 183.905 102.170 184.125 ;
        RECT 101.445 183.275 101.715 183.735 ;
        RECT 101.885 183.445 102.170 183.905 ;
        RECT 102.455 183.445 102.840 184.415 ;
        RECT 103.010 184.125 103.460 184.585 ;
        RECT 103.630 184.295 104.725 184.855 ;
        RECT 103.010 183.905 104.135 184.125 ;
        RECT 103.010 183.275 103.335 183.735 ;
        RECT 103.855 183.445 104.135 183.905 ;
        RECT 104.325 183.445 104.725 184.295 ;
        RECT 104.895 185.025 105.850 185.195 ;
        RECT 107.080 185.185 107.340 185.630 ;
        RECT 107.510 185.355 107.770 185.825 ;
        RECT 107.940 185.185 108.195 185.630 ;
        RECT 108.365 185.355 108.665 185.825 ;
        RECT 104.895 184.125 105.105 185.025 ;
        RECT 106.155 185.015 109.185 185.185 ;
        RECT 105.275 184.295 105.965 184.855 ;
        RECT 106.155 184.450 106.325 185.015 ;
        RECT 106.495 184.620 108.710 184.845 ;
        RECT 108.885 184.450 109.185 185.015 ;
        RECT 106.155 184.280 109.185 184.450 ;
        RECT 109.355 185.105 109.695 185.615 ;
        RECT 104.895 183.905 105.850 184.125 ;
        RECT 105.125 183.275 105.395 183.735 ;
        RECT 105.565 183.445 105.850 183.905 ;
        RECT 106.135 183.275 106.480 184.110 ;
        RECT 106.655 183.475 106.910 184.280 ;
        RECT 107.080 183.275 107.340 184.110 ;
        RECT 107.515 183.475 107.770 184.280 ;
        RECT 107.940 183.275 108.200 184.110 ;
        RECT 108.370 183.475 108.630 184.280 ;
        RECT 108.800 183.275 109.185 184.110 ;
        RECT 109.355 183.705 109.615 185.105 ;
        RECT 109.865 185.025 110.135 185.825 ;
        RECT 109.790 184.585 110.120 184.835 ;
        RECT 110.315 184.585 110.595 185.555 ;
        RECT 110.775 184.585 111.075 185.555 ;
        RECT 111.255 184.585 111.605 185.550 ;
        RECT 111.825 185.325 112.320 185.655 ;
        RECT 109.805 184.415 110.120 184.585 ;
        RECT 111.825 184.415 111.995 185.325 ;
        RECT 112.575 185.280 117.920 185.825 ;
        RECT 109.805 184.245 111.995 184.415 ;
        RECT 109.355 183.445 109.695 183.705 ;
        RECT 109.865 183.275 110.195 184.075 ;
        RECT 110.660 183.445 110.910 184.245 ;
        RECT 111.095 183.275 111.425 183.995 ;
        RECT 111.645 183.445 111.895 184.245 ;
        RECT 112.165 183.835 112.405 185.145 ;
        RECT 114.160 184.450 114.500 185.280 ;
        RECT 118.095 185.055 119.765 185.825 ;
        RECT 120.395 185.100 120.685 185.825 ;
        RECT 120.855 185.055 123.445 185.825 ;
        RECT 124.110 185.085 124.725 185.655 ;
        RECT 124.895 185.315 125.110 185.825 ;
        RECT 125.340 185.315 125.620 185.645 ;
        RECT 125.800 185.315 126.040 185.825 ;
        RECT 126.375 185.445 127.265 185.615 ;
        RECT 115.980 183.710 116.330 184.960 ;
        RECT 118.095 184.535 118.845 185.055 ;
        RECT 119.015 184.365 119.765 184.885 ;
        RECT 120.855 184.535 122.065 185.055 ;
        RECT 112.065 183.275 112.400 183.655 ;
        RECT 112.575 183.275 117.920 183.710 ;
        RECT 118.095 183.275 119.765 184.365 ;
        RECT 120.395 183.275 120.685 184.440 ;
        RECT 122.235 184.365 123.445 184.885 ;
        RECT 120.855 183.275 123.445 184.365 ;
        RECT 124.110 184.065 124.425 185.085 ;
        RECT 124.595 184.415 124.765 184.915 ;
        RECT 125.015 184.585 125.280 185.145 ;
        RECT 125.450 184.415 125.620 185.315 ;
        RECT 125.790 184.585 126.145 185.145 ;
        RECT 126.375 184.890 126.925 185.275 ;
        RECT 127.095 184.720 127.265 185.445 ;
        RECT 126.375 184.650 127.265 184.720 ;
        RECT 127.435 185.145 127.655 185.605 ;
        RECT 127.825 185.285 128.075 185.825 ;
        RECT 128.245 185.175 128.505 185.655 ;
        RECT 127.435 185.120 127.685 185.145 ;
        RECT 127.435 184.695 127.765 185.120 ;
        RECT 126.375 184.625 127.270 184.650 ;
        RECT 126.375 184.610 127.280 184.625 ;
        RECT 126.375 184.595 127.285 184.610 ;
        RECT 126.375 184.590 127.295 184.595 ;
        RECT 126.375 184.580 127.300 184.590 ;
        RECT 126.375 184.570 127.305 184.580 ;
        RECT 126.375 184.565 127.315 184.570 ;
        RECT 126.375 184.555 127.325 184.565 ;
        RECT 126.375 184.550 127.335 184.555 ;
        RECT 124.595 184.245 126.020 184.415 ;
        RECT 124.110 183.445 124.645 184.065 ;
        RECT 124.815 183.275 125.145 184.075 ;
        RECT 125.630 184.070 126.020 184.245 ;
        RECT 126.375 184.100 126.635 184.550 ;
        RECT 127.000 184.545 127.335 184.550 ;
        RECT 127.000 184.540 127.350 184.545 ;
        RECT 127.000 184.530 127.365 184.540 ;
        RECT 127.000 184.525 127.390 184.530 ;
        RECT 127.935 184.525 128.165 184.920 ;
        RECT 127.000 184.520 128.165 184.525 ;
        RECT 127.030 184.485 128.165 184.520 ;
        RECT 127.065 184.460 128.165 184.485 ;
        RECT 127.095 184.430 128.165 184.460 ;
        RECT 127.115 184.400 128.165 184.430 ;
        RECT 127.135 184.370 128.165 184.400 ;
        RECT 127.205 184.360 128.165 184.370 ;
        RECT 127.230 184.350 128.165 184.360 ;
        RECT 127.250 184.335 128.165 184.350 ;
        RECT 127.270 184.320 128.165 184.335 ;
        RECT 127.275 184.310 128.060 184.320 ;
        RECT 127.290 184.275 128.060 184.310 ;
        RECT 126.805 183.955 127.135 184.200 ;
        RECT 127.305 184.025 128.060 184.275 ;
        RECT 128.335 184.145 128.505 185.175 ;
        RECT 128.685 185.015 128.955 185.825 ;
        RECT 129.125 185.015 129.455 185.655 ;
        RECT 129.625 185.015 129.865 185.825 ;
        RECT 130.975 185.025 131.285 185.825 ;
        RECT 131.490 185.025 132.185 185.655 ;
        RECT 132.685 185.425 133.015 185.825 ;
        RECT 133.185 185.255 133.515 185.595 ;
        RECT 134.565 185.425 134.895 185.825 ;
        RECT 132.530 185.085 134.895 185.255 ;
        RECT 135.065 185.100 135.395 185.610 ;
        RECT 135.580 185.425 135.915 185.825 ;
        RECT 136.085 185.255 136.290 185.655 ;
        RECT 136.500 185.345 136.775 185.825 ;
        RECT 136.985 185.325 137.245 185.655 ;
        RECT 128.675 184.585 129.025 184.835 ;
        RECT 129.195 184.415 129.365 185.015 ;
        RECT 129.535 184.585 129.885 184.835 ;
        RECT 130.985 184.585 131.320 184.855 ;
        RECT 131.490 184.425 131.660 185.025 ;
        RECT 131.830 184.585 132.165 184.835 ;
        RECT 126.805 183.930 126.990 183.955 ;
        RECT 126.375 183.830 126.990 183.930 ;
        RECT 126.375 183.275 126.980 183.830 ;
        RECT 127.155 183.445 127.635 183.785 ;
        RECT 127.805 183.275 128.060 183.820 ;
        RECT 128.230 183.445 128.505 184.145 ;
        RECT 128.685 183.275 129.015 184.415 ;
        RECT 129.195 184.245 129.875 184.415 ;
        RECT 129.545 183.460 129.875 184.245 ;
        RECT 130.975 183.275 131.255 184.415 ;
        RECT 131.425 183.445 131.755 184.425 ;
        RECT 131.925 183.275 132.185 184.415 ;
        RECT 132.530 184.085 132.700 185.085 ;
        RECT 134.725 184.915 134.895 185.085 ;
        RECT 132.870 184.255 133.115 184.915 ;
        RECT 133.330 184.255 133.595 184.915 ;
        RECT 133.790 184.255 134.075 184.915 ;
        RECT 134.250 184.585 134.555 184.915 ;
        RECT 134.725 184.585 135.035 184.915 ;
        RECT 134.250 184.255 134.465 184.585 ;
        RECT 132.530 183.915 132.985 184.085 ;
        RECT 132.655 183.485 132.985 183.915 ;
        RECT 133.165 183.915 134.455 184.085 ;
        RECT 133.165 183.495 133.415 183.915 ;
        RECT 133.645 183.275 133.975 183.745 ;
        RECT 134.205 183.495 134.455 183.915 ;
        RECT 134.645 183.275 134.895 184.415 ;
        RECT 135.205 184.335 135.395 185.100 ;
        RECT 135.065 183.485 135.395 184.335 ;
        RECT 135.605 185.085 136.290 185.255 ;
        RECT 135.605 184.055 135.945 185.085 ;
        RECT 136.115 184.415 136.365 184.915 ;
        RECT 136.545 184.585 136.905 185.165 ;
        RECT 137.075 184.415 137.245 185.325 ;
        RECT 137.505 185.275 137.675 185.565 ;
        RECT 137.845 185.445 138.175 185.825 ;
        RECT 137.505 185.105 138.170 185.275 ;
        RECT 136.115 184.245 137.245 184.415 ;
        RECT 137.420 184.285 137.770 184.935 ;
        RECT 135.605 183.880 136.270 184.055 ;
        RECT 135.580 183.275 135.915 183.700 ;
        RECT 136.085 183.475 136.270 183.880 ;
        RECT 136.475 183.275 136.805 184.055 ;
        RECT 136.975 183.475 137.245 184.245 ;
        RECT 137.940 184.115 138.170 185.105 ;
        RECT 137.505 183.945 138.170 184.115 ;
        RECT 137.505 183.445 137.675 183.945 ;
        RECT 137.845 183.275 138.175 183.775 ;
        RECT 138.345 183.445 138.530 185.565 ;
        RECT 138.785 185.365 139.035 185.825 ;
        RECT 139.205 185.375 139.540 185.545 ;
        RECT 139.735 185.375 140.410 185.545 ;
        RECT 139.205 185.235 139.375 185.375 ;
        RECT 138.700 184.245 138.980 185.195 ;
        RECT 139.150 185.105 139.375 185.235 ;
        RECT 139.150 184.000 139.320 185.105 ;
        RECT 139.545 184.955 140.070 185.175 ;
        RECT 139.490 184.190 139.730 184.785 ;
        RECT 139.900 184.255 140.070 184.955 ;
        RECT 140.240 184.595 140.410 185.375 ;
        RECT 140.730 185.325 141.100 185.825 ;
        RECT 141.280 185.375 141.685 185.545 ;
        RECT 141.855 185.375 142.640 185.545 ;
        RECT 141.280 185.145 141.450 185.375 ;
        RECT 140.620 184.845 141.450 185.145 ;
        RECT 141.835 184.875 142.300 185.205 ;
        RECT 140.620 184.815 140.820 184.845 ;
        RECT 140.940 184.595 141.110 184.665 ;
        RECT 140.240 184.425 141.110 184.595 ;
        RECT 140.600 184.335 141.110 184.425 ;
        RECT 139.150 183.870 139.455 184.000 ;
        RECT 139.900 183.890 140.430 184.255 ;
        RECT 138.770 183.275 139.035 183.735 ;
        RECT 139.205 183.445 139.455 183.870 ;
        RECT 140.600 183.720 140.770 184.335 ;
        RECT 139.665 183.550 140.770 183.720 ;
        RECT 140.940 183.275 141.110 184.075 ;
        RECT 141.280 183.775 141.450 184.845 ;
        RECT 141.620 183.945 141.810 184.665 ;
        RECT 141.980 183.915 142.300 184.875 ;
        RECT 142.470 184.915 142.640 185.375 ;
        RECT 142.915 185.295 143.125 185.825 ;
        RECT 143.385 185.085 143.715 185.610 ;
        RECT 143.885 185.215 144.055 185.825 ;
        RECT 144.225 185.170 144.555 185.605 ;
        RECT 144.225 185.085 144.605 185.170 ;
        RECT 143.515 184.915 143.715 185.085 ;
        RECT 144.380 185.045 144.605 185.085 ;
        RECT 145.695 185.075 146.905 185.825 ;
        RECT 142.470 184.585 143.345 184.915 ;
        RECT 143.515 184.585 144.265 184.915 ;
        RECT 141.280 183.445 141.530 183.775 ;
        RECT 142.470 183.745 142.640 184.585 ;
        RECT 143.515 184.380 143.705 184.585 ;
        RECT 144.435 184.465 144.605 185.045 ;
        RECT 144.390 184.415 144.605 184.465 ;
        RECT 142.810 184.005 143.705 184.380 ;
        RECT 144.215 184.335 144.605 184.415 ;
        RECT 145.695 184.365 146.215 184.905 ;
        RECT 146.385 184.535 146.905 185.075 ;
        RECT 141.755 183.575 142.640 183.745 ;
        RECT 142.820 183.275 143.135 183.775 ;
        RECT 143.365 183.445 143.705 184.005 ;
        RECT 143.875 183.275 144.045 184.285 ;
        RECT 144.215 183.490 144.545 184.335 ;
        RECT 145.695 183.275 146.905 184.365 ;
        RECT 17.270 183.105 146.990 183.275 ;
        RECT 17.355 182.015 18.565 183.105 ;
        RECT 18.735 182.015 21.325 183.105 ;
        RECT 22.015 182.045 22.345 182.890 ;
        RECT 22.515 182.095 22.685 183.105 ;
        RECT 22.855 182.375 23.195 182.935 ;
        RECT 23.425 182.605 23.740 183.105 ;
        RECT 23.920 182.635 24.805 182.805 ;
        RECT 17.355 181.305 17.875 181.845 ;
        RECT 18.045 181.475 18.565 182.015 ;
        RECT 18.735 181.325 19.945 181.845 ;
        RECT 20.115 181.495 21.325 182.015 ;
        RECT 21.955 181.965 22.345 182.045 ;
        RECT 22.855 182.000 23.750 182.375 ;
        RECT 21.955 181.915 22.170 181.965 ;
        RECT 21.955 181.335 22.125 181.915 ;
        RECT 22.855 181.795 23.045 182.000 ;
        RECT 23.920 181.795 24.090 182.635 ;
        RECT 25.030 182.605 25.280 182.935 ;
        RECT 22.295 181.465 23.045 181.795 ;
        RECT 23.215 181.465 24.090 181.795 ;
        RECT 17.355 180.555 18.565 181.305 ;
        RECT 18.735 180.555 21.325 181.325 ;
        RECT 21.955 181.295 22.180 181.335 ;
        RECT 22.845 181.295 23.045 181.465 ;
        RECT 21.955 181.210 22.335 181.295 ;
        RECT 22.005 180.775 22.335 181.210 ;
        RECT 22.505 180.555 22.675 181.165 ;
        RECT 22.845 180.770 23.175 181.295 ;
        RECT 23.435 180.555 23.645 181.085 ;
        RECT 23.920 181.005 24.090 181.465 ;
        RECT 24.260 181.505 24.580 182.465 ;
        RECT 24.750 181.715 24.940 182.435 ;
        RECT 25.110 181.535 25.280 182.605 ;
        RECT 25.450 182.305 25.620 183.105 ;
        RECT 25.790 182.660 26.895 182.830 ;
        RECT 25.790 182.045 25.960 182.660 ;
        RECT 27.105 182.510 27.355 182.935 ;
        RECT 27.525 182.645 27.790 183.105 ;
        RECT 26.130 182.125 26.660 182.490 ;
        RECT 27.105 182.380 27.410 182.510 ;
        RECT 25.450 181.955 25.960 182.045 ;
        RECT 25.450 181.785 26.320 181.955 ;
        RECT 25.450 181.715 25.620 181.785 ;
        RECT 25.740 181.535 25.940 181.565 ;
        RECT 24.260 181.175 24.725 181.505 ;
        RECT 25.110 181.235 25.940 181.535 ;
        RECT 25.110 181.005 25.280 181.235 ;
        RECT 23.920 180.835 24.705 181.005 ;
        RECT 24.875 180.835 25.280 181.005 ;
        RECT 25.460 180.555 25.830 181.055 ;
        RECT 26.150 181.005 26.320 181.785 ;
        RECT 26.490 181.425 26.660 182.125 ;
        RECT 26.830 181.595 27.070 182.190 ;
        RECT 26.490 181.205 27.015 181.425 ;
        RECT 27.240 181.275 27.410 182.380 ;
        RECT 27.185 181.145 27.410 181.275 ;
        RECT 27.580 181.185 27.860 182.135 ;
        RECT 27.185 181.005 27.355 181.145 ;
        RECT 26.150 180.835 26.825 181.005 ;
        RECT 27.020 180.835 27.355 181.005 ;
        RECT 27.525 180.555 27.775 181.015 ;
        RECT 28.030 180.815 28.215 182.935 ;
        RECT 28.385 182.605 28.715 183.105 ;
        RECT 28.885 182.435 29.055 182.935 ;
        RECT 28.390 182.265 29.055 182.435 ;
        RECT 28.390 181.275 28.620 182.265 ;
        RECT 28.790 181.445 29.140 182.095 ;
        RECT 30.235 181.940 30.525 183.105 ;
        RECT 30.695 182.670 36.040 183.105 ;
        RECT 28.390 181.105 29.055 181.275 ;
        RECT 28.385 180.555 28.715 180.935 ;
        RECT 28.885 180.815 29.055 181.105 ;
        RECT 30.235 180.555 30.525 181.280 ;
        RECT 32.280 181.100 32.620 181.930 ;
        RECT 34.100 181.420 34.450 182.670 ;
        RECT 36.215 182.015 37.425 183.105 ;
        RECT 37.605 182.305 37.935 183.105 ;
        RECT 38.115 182.765 39.545 182.935 ;
        RECT 38.115 182.135 38.365 182.765 ;
        RECT 36.215 181.305 36.735 181.845 ;
        RECT 36.905 181.475 37.425 182.015 ;
        RECT 37.595 181.965 38.365 182.135 ;
        RECT 30.695 180.555 36.040 181.100 ;
        RECT 36.215 180.555 37.425 181.305 ;
        RECT 37.595 181.295 37.765 181.965 ;
        RECT 37.935 181.465 38.340 181.795 ;
        RECT 38.555 181.465 38.805 182.595 ;
        RECT 39.005 181.795 39.205 182.595 ;
        RECT 39.375 182.085 39.545 182.765 ;
        RECT 39.715 182.255 40.030 183.105 ;
        RECT 40.205 182.305 40.645 182.935 ;
        RECT 39.375 181.915 40.165 182.085 ;
        RECT 39.005 181.465 39.250 181.795 ;
        RECT 39.435 181.465 39.825 181.745 ;
        RECT 39.995 181.465 40.165 181.915 ;
        RECT 40.335 181.295 40.645 182.305 ;
        RECT 37.595 180.725 38.085 181.295 ;
        RECT 38.255 181.125 39.415 181.295 ;
        RECT 38.255 180.725 38.485 181.125 ;
        RECT 38.655 180.555 39.075 180.955 ;
        RECT 39.245 180.725 39.415 181.125 ;
        RECT 39.585 180.555 40.035 181.295 ;
        RECT 40.205 180.735 40.645 181.295 ;
        RECT 40.815 181.995 41.075 182.935 ;
        RECT 41.245 182.705 41.575 183.105 ;
        RECT 42.720 182.840 42.975 182.935 ;
        RECT 41.835 182.670 42.975 182.840 ;
        RECT 43.145 182.725 43.475 182.895 ;
        RECT 41.835 182.445 42.005 182.670 ;
        RECT 41.245 182.275 42.005 182.445 ;
        RECT 42.720 182.535 42.975 182.670 ;
        RECT 40.815 181.280 40.990 181.995 ;
        RECT 41.245 181.795 41.415 182.275 ;
        RECT 42.270 182.185 42.440 182.375 ;
        RECT 42.720 182.365 43.130 182.535 ;
        RECT 41.160 181.465 41.415 181.795 ;
        RECT 41.640 181.465 41.970 182.085 ;
        RECT 42.270 182.015 42.790 182.185 ;
        RECT 42.140 181.465 42.430 181.845 ;
        RECT 42.620 181.295 42.790 182.015 ;
        RECT 40.815 180.725 41.075 181.280 ;
        RECT 41.910 181.125 42.790 181.295 ;
        RECT 42.960 181.340 43.130 182.365 ;
        RECT 43.305 182.475 43.475 182.725 ;
        RECT 43.645 182.645 43.895 183.105 ;
        RECT 44.065 182.475 44.245 182.935 ;
        RECT 43.305 182.305 44.245 182.475 ;
        RECT 43.330 181.825 43.810 182.125 ;
        RECT 42.960 181.170 43.310 181.340 ;
        RECT 43.550 181.235 43.810 181.825 ;
        RECT 44.010 181.235 44.270 182.125 ;
        RECT 44.495 181.965 44.775 183.105 ;
        RECT 44.945 181.955 45.275 182.935 ;
        RECT 45.445 181.965 45.705 183.105 ;
        RECT 46.395 182.045 46.725 182.890 ;
        RECT 46.895 182.095 47.065 183.105 ;
        RECT 47.235 182.375 47.575 182.935 ;
        RECT 47.805 182.605 48.120 183.105 ;
        RECT 48.300 182.635 49.185 182.805 ;
        RECT 46.335 181.965 46.725 182.045 ;
        RECT 47.235 182.000 48.130 182.375 ;
        RECT 44.505 181.525 44.840 181.795 ;
        RECT 45.010 181.355 45.180 181.955 ;
        RECT 46.335 181.915 46.550 181.965 ;
        RECT 45.350 181.545 45.685 181.795 ;
        RECT 41.245 180.555 41.675 181.000 ;
        RECT 41.910 180.725 42.080 181.125 ;
        RECT 42.250 180.555 42.970 180.955 ;
        RECT 43.140 180.725 43.310 181.170 ;
        RECT 43.885 180.555 44.285 181.065 ;
        RECT 44.495 180.555 44.805 181.355 ;
        RECT 45.010 180.725 45.705 181.355 ;
        RECT 46.335 181.335 46.505 181.915 ;
        RECT 47.235 181.795 47.425 182.000 ;
        RECT 48.300 181.795 48.470 182.635 ;
        RECT 49.410 182.605 49.660 182.935 ;
        RECT 46.675 181.465 47.425 181.795 ;
        RECT 47.595 181.465 48.470 181.795 ;
        RECT 46.335 181.295 46.560 181.335 ;
        RECT 47.225 181.295 47.425 181.465 ;
        RECT 46.335 181.210 46.715 181.295 ;
        RECT 46.385 180.775 46.715 181.210 ;
        RECT 46.885 180.555 47.055 181.165 ;
        RECT 47.225 180.770 47.555 181.295 ;
        RECT 47.815 180.555 48.025 181.085 ;
        RECT 48.300 181.005 48.470 181.465 ;
        RECT 48.640 181.505 48.960 182.465 ;
        RECT 49.130 181.715 49.320 182.435 ;
        RECT 49.490 181.535 49.660 182.605 ;
        RECT 49.830 182.305 50.000 183.105 ;
        RECT 50.170 182.660 51.275 182.830 ;
        RECT 50.170 182.045 50.340 182.660 ;
        RECT 51.485 182.510 51.735 182.935 ;
        RECT 51.905 182.645 52.170 183.105 ;
        RECT 50.510 182.125 51.040 182.490 ;
        RECT 51.485 182.380 51.790 182.510 ;
        RECT 49.830 181.955 50.340 182.045 ;
        RECT 49.830 181.785 50.700 181.955 ;
        RECT 49.830 181.715 50.000 181.785 ;
        RECT 50.120 181.535 50.320 181.565 ;
        RECT 48.640 181.175 49.105 181.505 ;
        RECT 49.490 181.235 50.320 181.535 ;
        RECT 49.490 181.005 49.660 181.235 ;
        RECT 48.300 180.835 49.085 181.005 ;
        RECT 49.255 180.835 49.660 181.005 ;
        RECT 49.840 180.555 50.210 181.055 ;
        RECT 50.530 181.005 50.700 181.785 ;
        RECT 50.870 181.425 51.040 182.125 ;
        RECT 51.210 181.595 51.450 182.190 ;
        RECT 50.870 181.205 51.395 181.425 ;
        RECT 51.620 181.275 51.790 182.380 ;
        RECT 51.565 181.145 51.790 181.275 ;
        RECT 51.960 181.185 52.240 182.135 ;
        RECT 51.565 181.005 51.735 181.145 ;
        RECT 50.530 180.835 51.205 181.005 ;
        RECT 51.400 180.835 51.735 181.005 ;
        RECT 51.905 180.555 52.155 181.015 ;
        RECT 52.410 180.815 52.595 182.935 ;
        RECT 52.765 182.605 53.095 183.105 ;
        RECT 53.265 182.435 53.435 182.935 ;
        RECT 52.770 182.265 53.435 182.435 ;
        RECT 52.770 181.275 53.000 182.265 ;
        RECT 53.170 181.445 53.520 182.095 ;
        RECT 53.695 182.015 55.365 183.105 ;
        RECT 53.695 181.325 54.445 181.845 ;
        RECT 54.615 181.495 55.365 182.015 ;
        RECT 55.995 181.940 56.285 183.105 ;
        RECT 56.455 182.670 61.800 183.105 ;
        RECT 52.770 181.105 53.435 181.275 ;
        RECT 52.765 180.555 53.095 180.935 ;
        RECT 53.265 180.815 53.435 181.105 ;
        RECT 53.695 180.555 55.365 181.325 ;
        RECT 55.995 180.555 56.285 181.280 ;
        RECT 58.040 181.100 58.380 181.930 ;
        RECT 59.860 181.420 60.210 182.670 ;
        RECT 61.975 182.015 63.645 183.105 ;
        RECT 61.975 181.325 62.725 181.845 ;
        RECT 62.895 181.495 63.645 182.015 ;
        RECT 64.275 182.235 64.550 182.935 ;
        RECT 64.720 182.560 64.975 183.105 ;
        RECT 65.145 182.595 65.625 182.935 ;
        RECT 65.800 182.550 66.405 183.105 ;
        RECT 65.790 182.450 66.405 182.550 ;
        RECT 66.585 182.495 66.915 182.925 ;
        RECT 67.095 182.665 67.290 183.105 ;
        RECT 67.460 182.495 67.790 182.925 ;
        RECT 65.790 182.425 65.975 182.450 ;
        RECT 56.455 180.555 61.800 181.100 ;
        RECT 61.975 180.555 63.645 181.325 ;
        RECT 64.275 181.205 64.445 182.235 ;
        RECT 64.720 182.105 65.475 182.355 ;
        RECT 65.645 182.180 65.975 182.425 ;
        RECT 66.585 182.325 67.790 182.495 ;
        RECT 64.720 182.070 65.490 182.105 ;
        RECT 64.720 182.060 65.505 182.070 ;
        RECT 64.615 182.045 65.510 182.060 ;
        RECT 64.615 182.030 65.530 182.045 ;
        RECT 64.615 182.020 65.550 182.030 ;
        RECT 64.615 182.010 65.575 182.020 ;
        RECT 64.615 181.980 65.645 182.010 ;
        RECT 64.615 181.950 65.665 181.980 ;
        RECT 64.615 181.920 65.685 181.950 ;
        RECT 64.615 181.895 65.715 181.920 ;
        RECT 64.615 181.860 65.750 181.895 ;
        RECT 64.615 181.855 65.780 181.860 ;
        RECT 64.615 181.460 64.845 181.855 ;
        RECT 65.390 181.850 65.780 181.855 ;
        RECT 65.415 181.840 65.780 181.850 ;
        RECT 65.430 181.835 65.780 181.840 ;
        RECT 65.445 181.830 65.780 181.835 ;
        RECT 66.145 181.830 66.405 182.280 ;
        RECT 66.585 181.995 67.480 182.325 ;
        RECT 67.960 182.155 68.235 182.925 ;
        RECT 65.445 181.825 66.405 181.830 ;
        RECT 65.455 181.815 66.405 181.825 ;
        RECT 65.465 181.810 66.405 181.815 ;
        RECT 65.475 181.800 66.405 181.810 ;
        RECT 65.480 181.790 66.405 181.800 ;
        RECT 67.650 181.965 68.235 182.155 ;
        RECT 68.425 182.135 68.755 182.920 ;
        RECT 68.425 181.965 69.105 182.135 ;
        RECT 69.285 181.965 69.615 183.105 ;
        RECT 70.915 182.435 71.195 183.105 ;
        RECT 71.365 182.215 71.665 182.765 ;
        RECT 71.865 182.385 72.195 183.105 ;
        RECT 72.385 182.385 72.845 182.935 ;
        RECT 65.485 181.785 66.405 181.790 ;
        RECT 65.495 181.770 66.405 181.785 ;
        RECT 65.500 181.755 66.405 181.770 ;
        RECT 65.510 181.730 66.405 181.755 ;
        RECT 65.015 181.260 65.345 181.685 ;
        RECT 65.095 181.235 65.345 181.260 ;
        RECT 64.275 180.725 64.535 181.205 ;
        RECT 64.705 180.555 64.955 181.095 ;
        RECT 65.125 180.775 65.345 181.235 ;
        RECT 65.515 181.660 66.405 181.730 ;
        RECT 65.515 180.935 65.685 181.660 ;
        RECT 65.855 181.105 66.405 181.490 ;
        RECT 66.590 181.465 66.885 181.795 ;
        RECT 67.065 181.465 67.480 181.795 ;
        RECT 65.515 180.765 66.405 180.935 ;
        RECT 66.585 180.555 66.885 181.285 ;
        RECT 67.065 180.845 67.295 181.465 ;
        RECT 67.650 181.295 67.825 181.965 ;
        RECT 67.495 181.115 67.825 181.295 ;
        RECT 67.995 181.145 68.235 181.795 ;
        RECT 68.415 181.545 68.765 181.795 ;
        RECT 68.935 181.365 69.105 181.965 ;
        RECT 70.730 181.795 70.995 182.155 ;
        RECT 71.365 182.045 72.305 182.215 ;
        RECT 72.135 181.795 72.305 182.045 ;
        RECT 69.275 181.545 69.625 181.795 ;
        RECT 70.730 181.545 71.405 181.795 ;
        RECT 71.625 181.545 71.965 181.795 ;
        RECT 72.135 181.465 72.425 181.795 ;
        RECT 72.135 181.375 72.305 181.465 ;
        RECT 67.495 180.735 67.720 181.115 ;
        RECT 67.890 180.555 68.220 180.945 ;
        RECT 68.435 180.555 68.675 181.365 ;
        RECT 68.845 180.725 69.175 181.365 ;
        RECT 69.345 180.555 69.615 181.365 ;
        RECT 70.915 181.185 72.305 181.375 ;
        RECT 70.915 180.825 71.245 181.185 ;
        RECT 72.595 181.015 72.845 182.385 ;
        RECT 73.075 182.045 73.405 182.890 ;
        RECT 73.575 182.095 73.745 183.105 ;
        RECT 73.915 182.375 74.255 182.935 ;
        RECT 74.485 182.605 74.800 183.105 ;
        RECT 74.980 182.635 75.865 182.805 ;
        RECT 73.015 181.965 73.405 182.045 ;
        RECT 73.915 182.000 74.810 182.375 ;
        RECT 73.015 181.915 73.230 181.965 ;
        RECT 73.015 181.335 73.185 181.915 ;
        RECT 73.915 181.795 74.105 182.000 ;
        RECT 74.980 181.795 75.150 182.635 ;
        RECT 76.090 182.605 76.340 182.935 ;
        RECT 73.355 181.465 74.105 181.795 ;
        RECT 74.275 181.465 75.150 181.795 ;
        RECT 73.015 181.295 73.240 181.335 ;
        RECT 73.905 181.295 74.105 181.465 ;
        RECT 73.015 181.210 73.395 181.295 ;
        RECT 71.865 180.555 72.115 181.015 ;
        RECT 72.285 180.725 72.845 181.015 ;
        RECT 73.065 180.775 73.395 181.210 ;
        RECT 73.565 180.555 73.735 181.165 ;
        RECT 73.905 180.770 74.235 181.295 ;
        RECT 74.495 180.555 74.705 181.085 ;
        RECT 74.980 181.005 75.150 181.465 ;
        RECT 75.320 181.505 75.640 182.465 ;
        RECT 75.810 181.715 76.000 182.435 ;
        RECT 76.170 181.535 76.340 182.605 ;
        RECT 76.510 182.305 76.680 183.105 ;
        RECT 76.850 182.660 77.955 182.830 ;
        RECT 76.850 182.045 77.020 182.660 ;
        RECT 78.165 182.510 78.415 182.935 ;
        RECT 78.585 182.645 78.850 183.105 ;
        RECT 77.190 182.125 77.720 182.490 ;
        RECT 78.165 182.380 78.470 182.510 ;
        RECT 76.510 181.955 77.020 182.045 ;
        RECT 76.510 181.785 77.380 181.955 ;
        RECT 76.510 181.715 76.680 181.785 ;
        RECT 76.800 181.535 77.000 181.565 ;
        RECT 75.320 181.175 75.785 181.505 ;
        RECT 76.170 181.235 77.000 181.535 ;
        RECT 76.170 181.005 76.340 181.235 ;
        RECT 74.980 180.835 75.765 181.005 ;
        RECT 75.935 180.835 76.340 181.005 ;
        RECT 76.520 180.555 76.890 181.055 ;
        RECT 77.210 181.005 77.380 181.785 ;
        RECT 77.550 181.425 77.720 182.125 ;
        RECT 77.890 181.595 78.130 182.190 ;
        RECT 77.550 181.205 78.075 181.425 ;
        RECT 78.300 181.275 78.470 182.380 ;
        RECT 78.245 181.145 78.470 181.275 ;
        RECT 78.640 181.185 78.920 182.135 ;
        RECT 78.245 181.005 78.415 181.145 ;
        RECT 77.210 180.835 77.885 181.005 ;
        RECT 78.080 180.835 78.415 181.005 ;
        RECT 78.585 180.555 78.835 181.015 ;
        RECT 79.090 180.815 79.275 182.935 ;
        RECT 79.445 182.605 79.775 183.105 ;
        RECT 79.945 182.435 80.115 182.935 ;
        RECT 79.450 182.265 80.115 182.435 ;
        RECT 79.450 181.275 79.680 182.265 ;
        RECT 79.850 181.445 80.200 182.095 ;
        RECT 80.375 182.015 81.585 183.105 ;
        RECT 80.375 181.305 80.895 181.845 ;
        RECT 81.065 181.475 81.585 182.015 ;
        RECT 81.755 181.940 82.045 183.105 ;
        RECT 82.215 182.015 85.725 183.105 ;
        RECT 86.445 182.435 86.615 182.935 ;
        RECT 86.785 182.605 87.115 183.105 ;
        RECT 86.445 182.265 87.110 182.435 ;
        RECT 82.215 181.325 83.865 181.845 ;
        RECT 84.035 181.495 85.725 182.015 ;
        RECT 86.360 181.445 86.710 182.095 ;
        RECT 79.450 181.105 80.115 181.275 ;
        RECT 79.445 180.555 79.775 180.935 ;
        RECT 79.945 180.815 80.115 181.105 ;
        RECT 80.375 180.555 81.585 181.305 ;
        RECT 81.755 180.555 82.045 181.280 ;
        RECT 82.215 180.555 85.725 181.325 ;
        RECT 86.880 181.275 87.110 182.265 ;
        RECT 86.445 181.105 87.110 181.275 ;
        RECT 86.445 180.815 86.615 181.105 ;
        RECT 86.785 180.555 87.115 180.935 ;
        RECT 87.285 180.815 87.470 182.935 ;
        RECT 87.710 182.645 87.975 183.105 ;
        RECT 88.145 182.510 88.395 182.935 ;
        RECT 88.605 182.660 89.710 182.830 ;
        RECT 88.090 182.380 88.395 182.510 ;
        RECT 87.640 181.185 87.920 182.135 ;
        RECT 88.090 181.275 88.260 182.380 ;
        RECT 88.430 181.595 88.670 182.190 ;
        RECT 88.840 182.125 89.370 182.490 ;
        RECT 88.840 181.425 89.010 182.125 ;
        RECT 89.540 182.045 89.710 182.660 ;
        RECT 89.880 182.305 90.050 183.105 ;
        RECT 90.220 182.605 90.470 182.935 ;
        RECT 90.695 182.635 91.580 182.805 ;
        RECT 89.540 181.955 90.050 182.045 ;
        RECT 88.090 181.145 88.315 181.275 ;
        RECT 88.485 181.205 89.010 181.425 ;
        RECT 89.180 181.785 90.050 181.955 ;
        RECT 87.725 180.555 87.975 181.015 ;
        RECT 88.145 181.005 88.315 181.145 ;
        RECT 89.180 181.005 89.350 181.785 ;
        RECT 89.880 181.715 90.050 181.785 ;
        RECT 89.560 181.535 89.760 181.565 ;
        RECT 90.220 181.535 90.390 182.605 ;
        RECT 90.560 181.715 90.750 182.435 ;
        RECT 89.560 181.235 90.390 181.535 ;
        RECT 90.920 181.505 91.240 182.465 ;
        RECT 88.145 180.835 88.480 181.005 ;
        RECT 88.675 180.835 89.350 181.005 ;
        RECT 89.670 180.555 90.040 181.055 ;
        RECT 90.220 181.005 90.390 181.235 ;
        RECT 90.775 181.175 91.240 181.505 ;
        RECT 91.410 181.795 91.580 182.635 ;
        RECT 91.760 182.605 92.075 183.105 ;
        RECT 92.305 182.375 92.645 182.935 ;
        RECT 91.750 182.000 92.645 182.375 ;
        RECT 92.815 182.095 92.985 183.105 ;
        RECT 92.455 181.795 92.645 182.000 ;
        RECT 93.155 182.045 93.485 182.890 ;
        RECT 93.155 181.965 93.545 182.045 ;
        RECT 93.330 181.915 93.545 181.965 ;
        RECT 91.410 181.465 92.285 181.795 ;
        RECT 92.455 181.465 93.205 181.795 ;
        RECT 91.410 181.005 91.580 181.465 ;
        RECT 92.455 181.295 92.655 181.465 ;
        RECT 93.375 181.335 93.545 181.915 ;
        RECT 93.320 181.295 93.545 181.335 ;
        RECT 90.220 180.835 90.625 181.005 ;
        RECT 90.795 180.835 91.580 181.005 ;
        RECT 91.855 180.555 92.065 181.085 ;
        RECT 92.325 180.770 92.655 181.295 ;
        RECT 93.165 181.210 93.545 181.295 ;
        RECT 93.720 181.965 94.055 182.935 ;
        RECT 94.225 181.965 94.395 183.105 ;
        RECT 94.565 182.765 96.595 182.935 ;
        RECT 93.720 181.295 93.890 181.965 ;
        RECT 94.565 181.795 94.735 182.765 ;
        RECT 94.060 181.465 94.315 181.795 ;
        RECT 94.540 181.465 94.735 181.795 ;
        RECT 94.905 182.425 96.030 182.595 ;
        RECT 94.145 181.295 94.315 181.465 ;
        RECT 94.905 181.295 95.075 182.425 ;
        RECT 92.825 180.555 92.995 181.165 ;
        RECT 93.165 180.775 93.495 181.210 ;
        RECT 93.720 180.725 93.975 181.295 ;
        RECT 94.145 181.125 95.075 181.295 ;
        RECT 95.245 182.085 96.255 182.255 ;
        RECT 95.245 181.285 95.415 182.085 ;
        RECT 94.900 181.090 95.075 181.125 ;
        RECT 94.145 180.555 94.475 180.955 ;
        RECT 94.900 180.725 95.430 181.090 ;
        RECT 95.620 181.065 95.895 181.885 ;
        RECT 95.615 180.895 95.895 181.065 ;
        RECT 95.620 180.725 95.895 180.895 ;
        RECT 96.065 180.725 96.255 182.085 ;
        RECT 96.425 182.100 96.595 182.765 ;
        RECT 96.765 182.345 96.935 183.105 ;
        RECT 97.170 182.345 97.685 182.755 ;
        RECT 96.425 181.910 97.175 182.100 ;
        RECT 97.345 181.535 97.685 182.345 ;
        RECT 97.855 182.015 100.445 183.105 ;
        RECT 96.455 181.365 97.685 181.535 ;
        RECT 96.435 180.555 96.945 181.090 ;
        RECT 97.165 180.760 97.410 181.365 ;
        RECT 97.855 181.325 99.065 181.845 ;
        RECT 99.235 181.495 100.445 182.015 ;
        RECT 100.620 181.965 100.955 182.935 ;
        RECT 101.125 181.965 101.295 183.105 ;
        RECT 101.465 182.765 103.495 182.935 ;
        RECT 97.855 180.555 100.445 181.325 ;
        RECT 100.620 181.295 100.790 181.965 ;
        RECT 101.465 181.795 101.635 182.765 ;
        RECT 100.960 181.465 101.215 181.795 ;
        RECT 101.440 181.465 101.635 181.795 ;
        RECT 101.805 182.425 102.930 182.595 ;
        RECT 101.045 181.295 101.215 181.465 ;
        RECT 101.805 181.295 101.975 182.425 ;
        RECT 100.620 180.725 100.875 181.295 ;
        RECT 101.045 181.125 101.975 181.295 ;
        RECT 102.145 182.085 103.155 182.255 ;
        RECT 102.145 181.285 102.315 182.085 ;
        RECT 101.800 181.090 101.975 181.125 ;
        RECT 101.045 180.555 101.375 180.955 ;
        RECT 101.800 180.725 102.330 181.090 ;
        RECT 102.520 181.065 102.795 181.885 ;
        RECT 102.515 180.895 102.795 181.065 ;
        RECT 102.520 180.725 102.795 180.895 ;
        RECT 102.965 180.725 103.155 182.085 ;
        RECT 103.325 182.100 103.495 182.765 ;
        RECT 103.665 182.345 103.835 183.105 ;
        RECT 104.070 182.345 104.585 182.755 ;
        RECT 103.325 181.910 104.075 182.100 ;
        RECT 104.245 181.535 104.585 182.345 ;
        RECT 105.685 181.965 106.015 183.105 ;
        RECT 106.545 182.135 106.875 182.920 ;
        RECT 106.195 181.965 106.875 182.135 ;
        RECT 105.675 181.545 106.025 181.795 ;
        RECT 103.355 181.365 104.585 181.535 ;
        RECT 106.195 181.365 106.365 181.965 ;
        RECT 107.515 181.940 107.805 183.105 ;
        RECT 108.065 182.435 108.235 182.935 ;
        RECT 108.405 182.605 108.735 183.105 ;
        RECT 108.065 182.265 108.730 182.435 ;
        RECT 106.535 181.545 106.885 181.795 ;
        RECT 107.980 181.445 108.330 182.095 ;
        RECT 103.335 180.555 103.845 181.090 ;
        RECT 104.065 180.760 104.310 181.365 ;
        RECT 105.685 180.555 105.955 181.365 ;
        RECT 106.125 180.725 106.455 181.365 ;
        RECT 106.625 180.555 106.865 181.365 ;
        RECT 107.515 180.555 107.805 181.280 ;
        RECT 108.500 181.275 108.730 182.265 ;
        RECT 108.065 181.105 108.730 181.275 ;
        RECT 108.065 180.815 108.235 181.105 ;
        RECT 108.405 180.555 108.735 180.935 ;
        RECT 108.905 180.815 109.090 182.935 ;
        RECT 109.330 182.645 109.595 183.105 ;
        RECT 109.765 182.510 110.015 182.935 ;
        RECT 110.225 182.660 111.330 182.830 ;
        RECT 109.710 182.380 110.015 182.510 ;
        RECT 109.260 181.185 109.540 182.135 ;
        RECT 109.710 181.275 109.880 182.380 ;
        RECT 110.050 181.595 110.290 182.190 ;
        RECT 110.460 182.125 110.990 182.490 ;
        RECT 110.460 181.425 110.630 182.125 ;
        RECT 111.160 182.045 111.330 182.660 ;
        RECT 111.500 182.305 111.670 183.105 ;
        RECT 111.840 182.605 112.090 182.935 ;
        RECT 112.315 182.635 113.200 182.805 ;
        RECT 111.160 181.955 111.670 182.045 ;
        RECT 109.710 181.145 109.935 181.275 ;
        RECT 110.105 181.205 110.630 181.425 ;
        RECT 110.800 181.785 111.670 181.955 ;
        RECT 109.345 180.555 109.595 181.015 ;
        RECT 109.765 181.005 109.935 181.145 ;
        RECT 110.800 181.005 110.970 181.785 ;
        RECT 111.500 181.715 111.670 181.785 ;
        RECT 111.180 181.535 111.380 181.565 ;
        RECT 111.840 181.535 112.010 182.605 ;
        RECT 112.180 181.715 112.370 182.435 ;
        RECT 111.180 181.235 112.010 181.535 ;
        RECT 112.540 181.505 112.860 182.465 ;
        RECT 109.765 180.835 110.100 181.005 ;
        RECT 110.295 180.835 110.970 181.005 ;
        RECT 111.290 180.555 111.660 181.055 ;
        RECT 111.840 181.005 112.010 181.235 ;
        RECT 112.395 181.175 112.860 181.505 ;
        RECT 113.030 181.795 113.200 182.635 ;
        RECT 113.380 182.605 113.695 183.105 ;
        RECT 113.925 182.375 114.265 182.935 ;
        RECT 113.370 182.000 114.265 182.375 ;
        RECT 114.435 182.095 114.605 183.105 ;
        RECT 114.075 181.795 114.265 182.000 ;
        RECT 114.775 182.045 115.105 182.890 ;
        RECT 115.335 182.670 120.680 183.105 ;
        RECT 114.775 181.965 115.165 182.045 ;
        RECT 114.950 181.915 115.165 181.965 ;
        RECT 113.030 181.465 113.905 181.795 ;
        RECT 114.075 181.465 114.825 181.795 ;
        RECT 113.030 181.005 113.200 181.465 ;
        RECT 114.075 181.295 114.275 181.465 ;
        RECT 114.995 181.335 115.165 181.915 ;
        RECT 114.940 181.295 115.165 181.335 ;
        RECT 111.840 180.835 112.245 181.005 ;
        RECT 112.415 180.835 113.200 181.005 ;
        RECT 113.475 180.555 113.685 181.085 ;
        RECT 113.945 180.770 114.275 181.295 ;
        RECT 114.785 181.210 115.165 181.295 ;
        RECT 114.445 180.555 114.615 181.165 ;
        RECT 114.785 180.775 115.115 181.210 ;
        RECT 116.920 181.100 117.260 181.930 ;
        RECT 118.740 181.420 119.090 182.670 ;
        RECT 120.855 182.015 122.525 183.105 ;
        RECT 120.855 181.325 121.605 181.845 ;
        RECT 121.775 181.495 122.525 182.015 ;
        RECT 123.155 181.965 123.435 183.105 ;
        RECT 123.605 181.955 123.935 182.935 ;
        RECT 124.105 181.965 124.365 183.105 ;
        RECT 124.535 182.670 129.880 183.105 ;
        RECT 123.165 181.525 123.500 181.795 ;
        RECT 123.670 181.355 123.840 181.955 ;
        RECT 124.010 181.545 124.345 181.795 ;
        RECT 115.335 180.555 120.680 181.100 ;
        RECT 120.855 180.555 122.525 181.325 ;
        RECT 123.155 180.555 123.465 181.355 ;
        RECT 123.670 180.725 124.365 181.355 ;
        RECT 126.120 181.100 126.460 181.930 ;
        RECT 127.940 181.420 128.290 182.670 ;
        RECT 130.525 181.965 130.855 183.105 ;
        RECT 131.385 182.135 131.715 182.920 ;
        RECT 131.035 181.965 131.715 182.135 ;
        RECT 131.905 181.965 132.235 183.105 ;
        RECT 132.765 182.135 133.095 182.920 ;
        RECT 132.415 181.965 133.095 182.135 ;
        RECT 130.515 181.545 130.865 181.795 ;
        RECT 131.035 181.365 131.205 181.965 ;
        RECT 131.375 181.545 131.725 181.795 ;
        RECT 131.895 181.545 132.245 181.795 ;
        RECT 132.415 181.365 132.585 181.965 ;
        RECT 133.275 181.940 133.565 183.105 ;
        RECT 133.745 182.135 134.075 182.920 ;
        RECT 133.745 181.965 134.425 182.135 ;
        RECT 134.605 181.965 134.935 183.105 ;
        RECT 136.040 182.715 136.375 182.935 ;
        RECT 137.380 182.725 137.735 183.105 ;
        RECT 136.040 182.095 136.295 182.715 ;
        RECT 136.545 182.555 136.775 182.595 ;
        RECT 137.905 182.555 138.155 182.935 ;
        RECT 136.545 182.355 138.155 182.555 ;
        RECT 136.545 182.265 136.730 182.355 ;
        RECT 137.320 182.345 138.155 182.355 ;
        RECT 138.405 182.325 138.655 183.105 ;
        RECT 138.825 182.255 139.085 182.935 ;
        RECT 136.885 182.155 137.215 182.185 ;
        RECT 136.885 182.095 138.685 182.155 ;
        RECT 136.040 181.985 138.745 182.095 ;
        RECT 132.755 181.545 133.105 181.795 ;
        RECT 133.735 181.545 134.085 181.795 ;
        RECT 134.255 181.365 134.425 181.965 ;
        RECT 136.040 181.925 137.215 181.985 ;
        RECT 138.545 181.950 138.745 181.985 ;
        RECT 134.595 181.545 134.945 181.795 ;
        RECT 136.035 181.545 136.525 181.745 ;
        RECT 136.715 181.545 137.190 181.755 ;
        RECT 124.535 180.555 129.880 181.100 ;
        RECT 130.525 180.555 130.795 181.365 ;
        RECT 130.965 180.725 131.295 181.365 ;
        RECT 131.465 180.555 131.705 181.365 ;
        RECT 131.905 180.555 132.175 181.365 ;
        RECT 132.345 180.725 132.675 181.365 ;
        RECT 132.845 180.555 133.085 181.365 ;
        RECT 133.275 180.555 133.565 181.280 ;
        RECT 133.755 180.555 133.995 181.365 ;
        RECT 134.165 180.725 134.495 181.365 ;
        RECT 134.665 180.555 134.935 181.365 ;
        RECT 136.040 180.555 136.495 181.320 ;
        RECT 136.970 181.145 137.190 181.545 ;
        RECT 137.435 181.545 137.765 181.755 ;
        RECT 137.435 181.145 137.645 181.545 ;
        RECT 137.935 181.510 138.345 181.815 ;
        RECT 138.575 181.375 138.745 181.950 ;
        RECT 138.475 181.255 138.745 181.375 ;
        RECT 137.900 181.210 138.745 181.255 ;
        RECT 137.900 181.085 138.655 181.210 ;
        RECT 137.900 180.935 138.070 181.085 ;
        RECT 138.915 181.055 139.085 182.255 ;
        RECT 139.315 181.965 139.525 183.105 ;
        RECT 139.695 181.955 140.025 182.935 ;
        RECT 140.195 181.965 140.425 183.105 ;
        RECT 140.635 181.965 140.895 183.105 ;
        RECT 141.065 181.955 141.395 182.935 ;
        RECT 141.565 181.965 141.845 183.105 ;
        RECT 142.015 182.015 145.525 183.105 ;
        RECT 136.770 180.725 138.070 180.935 ;
        RECT 138.325 180.555 138.655 180.915 ;
        RECT 138.825 180.725 139.085 181.055 ;
        RECT 139.315 180.555 139.525 181.375 ;
        RECT 139.695 181.355 139.945 181.955 ;
        RECT 141.155 181.915 141.330 181.955 ;
        RECT 140.115 181.545 140.445 181.795 ;
        RECT 140.655 181.545 140.990 181.795 ;
        RECT 139.695 180.725 140.025 181.355 ;
        RECT 140.195 180.555 140.425 181.375 ;
        RECT 141.160 181.355 141.330 181.915 ;
        RECT 141.500 181.525 141.835 181.795 ;
        RECT 140.635 180.725 141.330 181.355 ;
        RECT 141.535 180.555 141.845 181.355 ;
        RECT 142.015 181.325 143.665 181.845 ;
        RECT 143.835 181.495 145.525 182.015 ;
        RECT 145.695 182.015 146.905 183.105 ;
        RECT 145.695 181.475 146.215 182.015 ;
        RECT 142.015 180.555 145.525 181.325 ;
        RECT 146.385 181.305 146.905 181.845 ;
        RECT 145.695 180.555 146.905 181.305 ;
        RECT 17.270 180.385 146.990 180.555 ;
        RECT 17.355 179.635 18.565 180.385 ;
        RECT 18.735 179.840 24.080 180.385 ;
        RECT 24.255 179.840 29.600 180.385 ;
        RECT 17.355 179.095 17.875 179.635 ;
        RECT 18.045 178.925 18.565 179.465 ;
        RECT 20.320 179.010 20.660 179.840 ;
        RECT 17.355 177.835 18.565 178.925 ;
        RECT 22.140 178.270 22.490 179.520 ;
        RECT 25.840 179.010 26.180 179.840 ;
        RECT 29.775 179.615 33.285 180.385 ;
        RECT 33.455 179.635 34.665 180.385 ;
        RECT 34.835 179.745 35.175 180.150 ;
        RECT 35.345 179.915 35.515 180.385 ;
        RECT 35.685 179.745 35.935 180.150 ;
        RECT 27.660 178.270 28.010 179.520 ;
        RECT 29.775 179.095 31.425 179.615 ;
        RECT 31.595 178.925 33.285 179.445 ;
        RECT 33.455 179.095 33.975 179.635 ;
        RECT 34.835 179.565 35.935 179.745 ;
        RECT 36.105 179.780 36.355 180.150 ;
        RECT 36.525 179.905 36.970 180.075 ;
        RECT 37.140 180.045 37.360 180.090 ;
        RECT 34.145 178.925 34.665 179.465 ;
        RECT 36.105 179.395 36.275 179.780 ;
        RECT 18.735 177.835 24.080 178.270 ;
        RECT 24.255 177.835 29.600 178.270 ;
        RECT 29.775 177.835 33.285 178.925 ;
        RECT 33.455 177.835 34.665 178.925 ;
        RECT 34.835 178.825 35.180 179.395 ;
        RECT 35.350 179.145 35.910 179.395 ;
        RECT 36.080 179.225 36.275 179.395 ;
        RECT 34.835 177.835 35.180 178.655 ;
        RECT 35.350 178.045 35.525 179.145 ;
        RECT 36.080 178.975 36.250 179.225 ;
        RECT 36.525 179.115 36.695 179.905 ;
        RECT 37.140 179.875 37.365 180.045 ;
        RECT 37.140 179.735 37.360 179.875 ;
        RECT 36.865 179.565 37.360 179.735 ;
        RECT 37.640 179.720 37.810 180.385 ;
        RECT 38.005 179.645 38.345 180.215 ;
        RECT 38.680 179.875 38.920 180.385 ;
        RECT 39.100 179.875 39.380 180.205 ;
        RECT 39.610 179.875 39.825 180.385 ;
        RECT 36.865 179.370 37.040 179.565 ;
        RECT 37.210 179.195 37.660 179.395 ;
        RECT 35.695 178.585 36.250 178.975 ;
        RECT 36.420 178.975 36.695 179.115 ;
        RECT 37.830 179.025 38.000 179.475 ;
        RECT 36.420 178.755 37.435 178.975 ;
        RECT 37.605 178.855 38.000 179.025 ;
        RECT 37.605 178.585 37.775 178.855 ;
        RECT 38.170 178.675 38.345 179.645 ;
        RECT 38.575 179.145 38.930 179.705 ;
        RECT 39.100 178.975 39.270 179.875 ;
        RECT 39.440 179.145 39.705 179.705 ;
        RECT 39.995 179.645 40.610 180.215 ;
        RECT 39.955 178.975 40.125 179.475 ;
        RECT 35.695 178.415 37.775 178.585 ;
        RECT 35.695 178.180 36.025 178.415 ;
        RECT 36.315 177.835 36.715 178.235 ;
        RECT 37.585 177.835 37.915 178.235 ;
        RECT 38.085 178.005 38.345 178.675 ;
        RECT 38.700 178.805 40.125 178.975 ;
        RECT 38.700 178.630 39.090 178.805 ;
        RECT 39.575 177.835 39.905 178.635 ;
        RECT 40.295 178.625 40.610 179.645 ;
        RECT 40.815 179.615 42.485 180.385 ;
        RECT 43.115 179.660 43.405 180.385 ;
        RECT 43.575 179.660 43.835 180.215 ;
        RECT 44.005 179.940 44.435 180.385 ;
        RECT 44.670 179.815 44.840 180.215 ;
        RECT 45.010 179.985 45.730 180.385 ;
        RECT 40.815 179.095 41.565 179.615 ;
        RECT 41.735 178.925 42.485 179.445 ;
        RECT 40.075 178.005 40.610 178.625 ;
        RECT 40.815 177.835 42.485 178.925 ;
        RECT 43.115 177.835 43.405 179.000 ;
        RECT 43.575 178.945 43.750 179.660 ;
        RECT 44.670 179.645 45.550 179.815 ;
        RECT 45.900 179.770 46.070 180.215 ;
        RECT 46.645 179.875 47.045 180.385 ;
        RECT 47.305 179.995 47.635 180.385 ;
        RECT 47.805 179.815 47.975 180.135 ;
        RECT 48.145 179.995 48.475 180.385 ;
        RECT 48.890 179.985 49.845 180.155 ;
        RECT 43.920 179.145 44.175 179.475 ;
        RECT 43.575 178.005 43.835 178.945 ;
        RECT 44.005 178.665 44.175 179.145 ;
        RECT 44.400 178.855 44.730 179.475 ;
        RECT 44.900 179.095 45.190 179.475 ;
        RECT 45.380 178.925 45.550 179.645 ;
        RECT 45.030 178.755 45.550 178.925 ;
        RECT 45.720 179.600 46.070 179.770 ;
        RECT 44.005 178.495 44.765 178.665 ;
        RECT 45.030 178.565 45.200 178.755 ;
        RECT 45.720 178.575 45.890 179.600 ;
        RECT 46.310 179.115 46.570 179.705 ;
        RECT 46.090 178.815 46.570 179.115 ;
        RECT 46.770 178.815 47.030 179.705 ;
        RECT 47.255 179.645 49.505 179.815 ;
        RECT 47.255 178.685 47.425 179.645 ;
        RECT 47.595 179.025 47.840 179.475 ;
        RECT 48.010 179.195 48.560 179.395 ;
        RECT 48.730 179.225 49.105 179.395 ;
        RECT 48.730 179.025 48.900 179.225 ;
        RECT 49.275 179.145 49.505 179.645 ;
        RECT 47.595 178.855 48.900 179.025 ;
        RECT 49.675 179.105 49.845 179.985 ;
        RECT 50.015 179.550 50.305 180.385 ;
        RECT 50.675 179.755 51.005 180.115 ;
        RECT 51.625 179.925 51.875 180.385 ;
        RECT 52.045 179.925 52.605 180.215 ;
        RECT 50.675 179.565 52.065 179.755 ;
        RECT 51.895 179.475 52.065 179.565 ;
        RECT 50.490 179.145 51.165 179.395 ;
        RECT 51.385 179.145 51.725 179.395 ;
        RECT 51.895 179.145 52.185 179.475 ;
        RECT 49.675 178.935 50.305 179.105 ;
        RECT 44.595 178.270 44.765 178.495 ;
        RECT 45.480 178.405 45.890 178.575 ;
        RECT 46.065 178.465 47.005 178.635 ;
        RECT 45.480 178.270 45.735 178.405 ;
        RECT 44.005 177.835 44.335 178.235 ;
        RECT 44.595 178.100 45.735 178.270 ;
        RECT 46.065 178.215 46.235 178.465 ;
        RECT 45.480 178.005 45.735 178.100 ;
        RECT 45.905 178.045 46.235 178.215 ;
        RECT 46.405 177.835 46.655 178.295 ;
        RECT 46.825 178.005 47.005 178.465 ;
        RECT 47.255 178.005 47.635 178.685 ;
        RECT 48.225 177.835 48.395 178.685 ;
        RECT 48.565 178.515 49.805 178.685 ;
        RECT 48.565 178.005 48.895 178.515 ;
        RECT 49.065 177.835 49.235 178.345 ;
        RECT 49.405 178.005 49.805 178.515 ;
        RECT 49.985 178.005 50.305 178.935 ;
        RECT 50.490 178.785 50.755 179.145 ;
        RECT 51.895 178.895 52.065 179.145 ;
        RECT 51.125 178.725 52.065 178.895 ;
        RECT 50.675 177.835 50.955 178.505 ;
        RECT 51.125 178.175 51.425 178.725 ;
        RECT 52.355 178.555 52.605 179.925 ;
        RECT 52.775 179.615 56.285 180.385 ;
        RECT 56.985 179.985 57.315 180.385 ;
        RECT 57.485 179.815 57.655 180.085 ;
        RECT 57.825 179.985 58.155 180.385 ;
        RECT 58.325 179.815 58.580 180.085 ;
        RECT 52.775 179.095 54.425 179.615 ;
        RECT 54.595 178.925 56.285 179.445 ;
        RECT 51.625 177.835 51.955 178.555 ;
        RECT 52.145 178.005 52.605 178.555 ;
        RECT 52.775 177.835 56.285 178.925 ;
        RECT 56.915 178.805 57.185 179.815 ;
        RECT 57.355 179.645 58.580 179.815 ;
        RECT 58.755 179.645 59.075 180.125 ;
        RECT 59.245 179.815 59.475 180.215 ;
        RECT 59.645 179.995 59.995 180.385 ;
        RECT 59.245 179.735 59.755 179.815 ;
        RECT 60.165 179.735 60.495 180.215 ;
        RECT 59.245 179.645 60.495 179.735 ;
        RECT 57.355 178.975 57.525 179.645 ;
        RECT 57.695 179.145 58.075 179.475 ;
        RECT 58.245 179.145 58.580 179.475 ;
        RECT 57.355 178.805 57.670 178.975 ;
        RECT 56.920 177.835 57.235 178.635 ;
        RECT 57.500 178.190 57.670 178.805 ;
        RECT 57.840 178.465 58.075 179.145 ;
        RECT 58.245 178.190 58.580 178.975 ;
        RECT 58.755 178.715 58.925 179.645 ;
        RECT 59.585 179.565 60.495 179.645 ;
        RECT 60.665 179.565 60.835 180.385 ;
        RECT 61.340 179.645 61.805 180.190 ;
        RECT 59.095 179.055 59.265 179.475 ;
        RECT 59.495 179.225 60.095 179.395 ;
        RECT 59.095 178.885 59.755 179.055 ;
        RECT 58.755 178.515 59.415 178.715 ;
        RECT 59.585 178.685 59.755 178.885 ;
        RECT 59.925 179.025 60.095 179.225 ;
        RECT 60.265 179.195 60.960 179.395 ;
        RECT 61.220 179.025 61.465 179.475 ;
        RECT 59.925 178.855 61.465 179.025 ;
        RECT 61.635 178.685 61.805 179.645 ;
        RECT 59.585 178.515 61.805 178.685 ;
        RECT 61.975 179.645 62.440 180.190 ;
        RECT 61.975 178.685 62.145 179.645 ;
        RECT 62.945 179.565 63.115 180.385 ;
        RECT 63.285 179.735 63.615 180.215 ;
        RECT 63.785 179.995 64.135 180.385 ;
        RECT 64.305 179.815 64.535 180.215 ;
        RECT 64.025 179.735 64.535 179.815 ;
        RECT 63.285 179.645 64.535 179.735 ;
        RECT 64.705 179.645 65.025 180.125 ;
        RECT 63.285 179.565 64.195 179.645 ;
        RECT 62.315 179.025 62.560 179.475 ;
        RECT 62.820 179.195 63.515 179.395 ;
        RECT 63.685 179.225 64.285 179.395 ;
        RECT 63.685 179.025 63.855 179.225 ;
        RECT 64.515 179.055 64.685 179.475 ;
        RECT 62.315 178.855 63.855 179.025 ;
        RECT 64.025 178.885 64.685 179.055 ;
        RECT 64.025 178.685 64.195 178.885 ;
        RECT 64.855 178.715 65.025 179.645 ;
        RECT 61.975 178.515 64.195 178.685 ;
        RECT 64.365 178.515 65.025 178.715 ;
        RECT 65.195 179.645 65.580 180.215 ;
        RECT 65.750 179.925 66.075 180.385 ;
        RECT 66.595 179.755 66.875 180.215 ;
        RECT 65.195 178.975 65.475 179.645 ;
        RECT 65.750 179.585 66.875 179.755 ;
        RECT 65.750 179.475 66.200 179.585 ;
        RECT 65.645 179.145 66.200 179.475 ;
        RECT 67.065 179.415 67.465 180.215 ;
        RECT 67.865 179.925 68.135 180.385 ;
        RECT 68.305 179.755 68.590 180.215 ;
        RECT 59.245 178.345 59.415 178.515 ;
        RECT 57.500 178.020 58.580 178.190 ;
        RECT 58.775 177.835 59.075 178.345 ;
        RECT 59.245 178.175 59.625 178.345 ;
        RECT 60.205 177.835 60.835 178.345 ;
        RECT 61.005 178.005 61.335 178.515 ;
        RECT 61.505 177.835 61.805 178.345 ;
        RECT 61.975 177.835 62.275 178.345 ;
        RECT 62.445 178.005 62.775 178.515 ;
        RECT 64.365 178.345 64.535 178.515 ;
        RECT 62.945 177.835 63.575 178.345 ;
        RECT 64.155 178.175 64.535 178.345 ;
        RECT 64.705 177.835 65.005 178.345 ;
        RECT 65.195 178.005 65.580 178.975 ;
        RECT 65.750 178.685 66.200 179.145 ;
        RECT 66.370 178.855 67.465 179.415 ;
        RECT 65.750 178.465 66.875 178.685 ;
        RECT 65.750 177.835 66.075 178.295 ;
        RECT 66.595 178.005 66.875 178.465 ;
        RECT 67.065 178.005 67.465 178.855 ;
        RECT 67.635 179.585 68.590 179.755 ;
        RECT 68.875 179.660 69.165 180.385 ;
        RECT 69.335 179.645 69.720 180.215 ;
        RECT 69.890 179.925 70.215 180.385 ;
        RECT 70.735 179.755 71.015 180.215 ;
        RECT 67.635 178.685 67.845 179.585 ;
        RECT 68.015 178.855 68.705 179.415 ;
        RECT 67.635 178.465 68.590 178.685 ;
        RECT 67.865 177.835 68.135 178.295 ;
        RECT 68.305 178.005 68.590 178.465 ;
        RECT 68.875 177.835 69.165 179.000 ;
        RECT 69.335 178.975 69.615 179.645 ;
        RECT 69.890 179.585 71.015 179.755 ;
        RECT 69.890 179.475 70.340 179.585 ;
        RECT 69.785 179.145 70.340 179.475 ;
        RECT 71.205 179.415 71.605 180.215 ;
        RECT 72.005 179.925 72.275 180.385 ;
        RECT 72.445 179.755 72.730 180.215 ;
        RECT 73.085 179.985 73.415 180.385 ;
        RECT 73.585 179.815 73.755 180.085 ;
        RECT 73.925 179.985 74.255 180.385 ;
        RECT 74.425 179.815 74.680 180.085 ;
        RECT 69.335 178.005 69.720 178.975 ;
        RECT 69.890 178.685 70.340 179.145 ;
        RECT 70.510 178.855 71.605 179.415 ;
        RECT 69.890 178.465 71.015 178.685 ;
        RECT 69.890 177.835 70.215 178.295 ;
        RECT 70.735 178.005 71.015 178.465 ;
        RECT 71.205 178.005 71.605 178.855 ;
        RECT 71.775 179.585 72.730 179.755 ;
        RECT 71.775 178.685 71.985 179.585 ;
        RECT 72.155 178.855 72.845 179.415 ;
        RECT 73.015 178.805 73.285 179.815 ;
        RECT 73.455 179.645 74.680 179.815 ;
        RECT 73.455 178.975 73.625 179.645 ;
        RECT 74.855 179.615 77.445 180.385 ;
        RECT 77.705 179.835 77.875 180.125 ;
        RECT 78.045 180.005 78.375 180.385 ;
        RECT 77.705 179.665 78.370 179.835 ;
        RECT 73.795 179.145 74.175 179.475 ;
        RECT 74.345 179.145 74.680 179.475 ;
        RECT 73.455 178.805 73.770 178.975 ;
        RECT 71.775 178.465 72.730 178.685 ;
        RECT 72.005 177.835 72.275 178.295 ;
        RECT 72.445 178.005 72.730 178.465 ;
        RECT 73.020 177.835 73.335 178.635 ;
        RECT 73.600 178.190 73.770 178.805 ;
        RECT 73.940 178.465 74.175 179.145 ;
        RECT 74.855 179.095 76.065 179.615 ;
        RECT 74.345 178.190 74.680 178.975 ;
        RECT 76.235 178.925 77.445 179.445 ;
        RECT 73.600 178.020 74.680 178.190 ;
        RECT 74.855 177.835 77.445 178.925 ;
        RECT 77.620 178.845 77.970 179.495 ;
        RECT 78.140 178.675 78.370 179.665 ;
        RECT 77.705 178.505 78.370 178.675 ;
        RECT 77.705 178.005 77.875 178.505 ;
        RECT 78.045 177.835 78.375 178.335 ;
        RECT 78.545 178.005 78.730 180.125 ;
        RECT 78.985 179.925 79.235 180.385 ;
        RECT 79.405 179.935 79.740 180.105 ;
        RECT 79.935 179.935 80.610 180.105 ;
        RECT 79.405 179.795 79.575 179.935 ;
        RECT 78.900 178.805 79.180 179.755 ;
        RECT 79.350 179.665 79.575 179.795 ;
        RECT 79.350 178.560 79.520 179.665 ;
        RECT 79.745 179.515 80.270 179.735 ;
        RECT 79.690 178.750 79.930 179.345 ;
        RECT 80.100 178.815 80.270 179.515 ;
        RECT 80.440 179.155 80.610 179.935 ;
        RECT 80.930 179.885 81.300 180.385 ;
        RECT 81.480 179.935 81.885 180.105 ;
        RECT 82.055 179.935 82.840 180.105 ;
        RECT 81.480 179.705 81.650 179.935 ;
        RECT 80.820 179.405 81.650 179.705 ;
        RECT 82.035 179.435 82.500 179.765 ;
        RECT 80.820 179.375 81.020 179.405 ;
        RECT 81.140 179.155 81.310 179.225 ;
        RECT 80.440 178.985 81.310 179.155 ;
        RECT 80.800 178.895 81.310 178.985 ;
        RECT 79.350 178.430 79.655 178.560 ;
        RECT 80.100 178.450 80.630 178.815 ;
        RECT 78.970 177.835 79.235 178.295 ;
        RECT 79.405 178.005 79.655 178.430 ;
        RECT 80.800 178.280 80.970 178.895 ;
        RECT 79.865 178.110 80.970 178.280 ;
        RECT 81.140 177.835 81.310 178.635 ;
        RECT 81.480 178.335 81.650 179.405 ;
        RECT 81.820 178.505 82.010 179.225 ;
        RECT 82.180 178.475 82.500 179.435 ;
        RECT 82.670 179.475 82.840 179.935 ;
        RECT 83.115 179.855 83.325 180.385 ;
        RECT 83.585 179.645 83.915 180.170 ;
        RECT 84.085 179.775 84.255 180.385 ;
        RECT 84.425 179.730 84.755 180.165 ;
        RECT 84.975 179.840 90.320 180.385 ;
        RECT 84.425 179.645 84.805 179.730 ;
        RECT 83.715 179.475 83.915 179.645 ;
        RECT 84.580 179.605 84.805 179.645 ;
        RECT 82.670 179.145 83.545 179.475 ;
        RECT 83.715 179.145 84.465 179.475 ;
        RECT 81.480 178.005 81.730 178.335 ;
        RECT 82.670 178.305 82.840 179.145 ;
        RECT 83.715 178.940 83.905 179.145 ;
        RECT 84.635 179.025 84.805 179.605 ;
        RECT 84.590 178.975 84.805 179.025 ;
        RECT 86.560 179.010 86.900 179.840 ;
        RECT 90.495 179.615 94.005 180.385 ;
        RECT 94.635 179.660 94.925 180.385 ;
        RECT 95.100 179.645 95.355 180.215 ;
        RECT 95.525 179.985 95.855 180.385 ;
        RECT 96.280 179.850 96.810 180.215 ;
        RECT 96.280 179.815 96.455 179.850 ;
        RECT 95.525 179.645 96.455 179.815 ;
        RECT 83.010 178.565 83.905 178.940 ;
        RECT 84.415 178.895 84.805 178.975 ;
        RECT 81.955 178.135 82.840 178.305 ;
        RECT 83.020 177.835 83.335 178.335 ;
        RECT 83.565 178.005 83.905 178.565 ;
        RECT 84.075 177.835 84.245 178.845 ;
        RECT 84.415 178.050 84.745 178.895 ;
        RECT 88.380 178.270 88.730 179.520 ;
        RECT 90.495 179.095 92.145 179.615 ;
        RECT 92.315 178.925 94.005 179.445 ;
        RECT 84.975 177.835 90.320 178.270 ;
        RECT 90.495 177.835 94.005 178.925 ;
        RECT 94.635 177.835 94.925 179.000 ;
        RECT 95.100 178.975 95.270 179.645 ;
        RECT 95.525 179.475 95.695 179.645 ;
        RECT 95.440 179.145 95.695 179.475 ;
        RECT 95.920 179.145 96.115 179.475 ;
        RECT 95.100 178.005 95.435 178.975 ;
        RECT 95.605 177.835 95.775 178.975 ;
        RECT 95.945 178.175 96.115 179.145 ;
        RECT 96.285 178.515 96.455 179.645 ;
        RECT 96.625 178.855 96.795 179.655 ;
        RECT 97.000 179.365 97.275 180.215 ;
        RECT 96.995 179.195 97.275 179.365 ;
        RECT 97.000 179.055 97.275 179.195 ;
        RECT 97.445 178.855 97.635 180.215 ;
        RECT 97.815 179.850 98.325 180.385 ;
        RECT 98.545 179.575 98.790 180.180 ;
        RECT 99.235 179.615 100.905 180.385 ;
        RECT 101.135 179.925 101.380 180.385 ;
        RECT 97.835 179.405 99.065 179.575 ;
        RECT 96.625 178.685 97.635 178.855 ;
        RECT 97.805 178.840 98.555 179.030 ;
        RECT 96.285 178.345 97.410 178.515 ;
        RECT 97.805 178.175 97.975 178.840 ;
        RECT 98.725 178.595 99.065 179.405 ;
        RECT 99.235 179.095 99.985 179.615 ;
        RECT 100.155 178.925 100.905 179.445 ;
        RECT 101.075 179.145 101.390 179.755 ;
        RECT 101.560 179.395 101.810 180.205 ;
        RECT 101.980 179.860 102.240 180.385 ;
        RECT 102.410 179.735 102.670 180.190 ;
        RECT 102.840 179.905 103.100 180.385 ;
        RECT 103.270 179.735 103.530 180.190 ;
        RECT 103.700 179.905 103.960 180.385 ;
        RECT 104.130 179.735 104.390 180.190 ;
        RECT 104.560 179.905 104.820 180.385 ;
        RECT 104.990 179.735 105.250 180.190 ;
        RECT 105.420 179.905 105.720 180.385 ;
        RECT 102.410 179.565 105.720 179.735 ;
        RECT 101.560 179.145 104.580 179.395 ;
        RECT 95.945 178.005 97.975 178.175 ;
        RECT 98.145 177.835 98.315 178.595 ;
        RECT 98.550 178.185 99.065 178.595 ;
        RECT 99.235 177.835 100.905 178.925 ;
        RECT 101.085 177.835 101.380 178.945 ;
        RECT 101.560 178.010 101.810 179.145 ;
        RECT 104.750 178.975 105.720 179.565 ;
        RECT 106.135 179.615 107.805 180.385 ;
        RECT 108.065 179.835 108.235 180.125 ;
        RECT 108.405 180.005 108.735 180.385 ;
        RECT 108.065 179.665 108.730 179.835 ;
        RECT 106.135 179.095 106.885 179.615 ;
        RECT 101.980 177.835 102.240 178.945 ;
        RECT 102.410 178.735 105.720 178.975 ;
        RECT 107.055 178.925 107.805 179.445 ;
        RECT 102.410 178.010 102.670 178.735 ;
        RECT 102.840 177.835 103.100 178.565 ;
        RECT 103.270 178.010 103.530 178.735 ;
        RECT 103.700 177.835 103.960 178.565 ;
        RECT 104.130 178.010 104.390 178.735 ;
        RECT 104.560 177.835 104.820 178.565 ;
        RECT 104.990 178.010 105.250 178.735 ;
        RECT 105.420 177.835 105.715 178.565 ;
        RECT 106.135 177.835 107.805 178.925 ;
        RECT 107.980 178.845 108.330 179.495 ;
        RECT 108.500 178.675 108.730 179.665 ;
        RECT 108.065 178.505 108.730 178.675 ;
        RECT 108.065 178.005 108.235 178.505 ;
        RECT 108.405 177.835 108.735 178.335 ;
        RECT 108.905 178.005 109.090 180.125 ;
        RECT 109.345 179.925 109.595 180.385 ;
        RECT 109.765 179.935 110.100 180.105 ;
        RECT 110.295 179.935 110.970 180.105 ;
        RECT 109.765 179.795 109.935 179.935 ;
        RECT 109.260 178.805 109.540 179.755 ;
        RECT 109.710 179.665 109.935 179.795 ;
        RECT 109.710 178.560 109.880 179.665 ;
        RECT 110.105 179.515 110.630 179.735 ;
        RECT 110.050 178.750 110.290 179.345 ;
        RECT 110.460 178.815 110.630 179.515 ;
        RECT 110.800 179.155 110.970 179.935 ;
        RECT 111.290 179.885 111.660 180.385 ;
        RECT 111.840 179.935 112.245 180.105 ;
        RECT 112.415 179.935 113.200 180.105 ;
        RECT 111.840 179.705 112.010 179.935 ;
        RECT 111.180 179.405 112.010 179.705 ;
        RECT 112.395 179.435 112.860 179.765 ;
        RECT 111.180 179.375 111.380 179.405 ;
        RECT 111.500 179.155 111.670 179.225 ;
        RECT 110.800 178.985 111.670 179.155 ;
        RECT 111.160 178.895 111.670 178.985 ;
        RECT 109.710 178.430 110.015 178.560 ;
        RECT 110.460 178.450 110.990 178.815 ;
        RECT 109.330 177.835 109.595 178.295 ;
        RECT 109.765 178.005 110.015 178.430 ;
        RECT 111.160 178.280 111.330 178.895 ;
        RECT 110.225 178.110 111.330 178.280 ;
        RECT 111.500 177.835 111.670 178.635 ;
        RECT 111.840 178.335 112.010 179.405 ;
        RECT 112.180 178.505 112.370 179.225 ;
        RECT 112.540 178.475 112.860 179.435 ;
        RECT 113.030 179.475 113.200 179.935 ;
        RECT 113.475 179.855 113.685 180.385 ;
        RECT 113.945 179.645 114.275 180.170 ;
        RECT 114.445 179.775 114.615 180.385 ;
        RECT 114.785 179.730 115.115 180.165 ;
        RECT 114.785 179.645 115.165 179.730 ;
        RECT 114.075 179.475 114.275 179.645 ;
        RECT 114.940 179.605 115.165 179.645 ;
        RECT 113.030 179.145 113.905 179.475 ;
        RECT 114.075 179.145 114.825 179.475 ;
        RECT 111.840 178.005 112.090 178.335 ;
        RECT 113.030 178.305 113.200 179.145 ;
        RECT 114.075 178.940 114.265 179.145 ;
        RECT 114.995 179.025 115.165 179.605 ;
        RECT 114.950 178.975 115.165 179.025 ;
        RECT 113.370 178.565 114.265 178.940 ;
        RECT 114.775 178.895 115.165 178.975 ;
        RECT 112.315 178.135 113.200 178.305 ;
        RECT 113.380 177.835 113.695 178.335 ;
        RECT 113.925 178.005 114.265 178.565 ;
        RECT 114.435 177.835 114.605 178.845 ;
        RECT 114.775 178.050 115.105 178.895 ;
        RECT 116.275 178.805 116.505 180.145 ;
        RECT 116.685 179.305 116.915 180.205 ;
        RECT 117.115 179.605 117.360 180.385 ;
        RECT 117.530 179.845 117.960 180.205 ;
        RECT 118.540 180.015 119.270 180.385 ;
        RECT 117.530 179.655 119.270 179.845 ;
        RECT 117.530 179.425 117.750 179.655 ;
        RECT 116.685 178.625 117.025 179.305 ;
        RECT 116.275 178.425 117.025 178.625 ;
        RECT 117.205 179.125 117.750 179.425 ;
        RECT 116.275 178.035 116.515 178.425 ;
        RECT 116.685 177.835 117.035 178.245 ;
        RECT 117.205 178.015 117.535 179.125 ;
        RECT 117.920 178.855 118.345 179.475 ;
        RECT 118.540 178.855 118.800 179.475 ;
        RECT 119.010 179.145 119.270 179.655 ;
        RECT 117.705 178.485 118.730 178.685 ;
        RECT 117.705 178.015 117.885 178.485 ;
        RECT 118.055 177.835 118.385 178.315 ;
        RECT 118.560 178.015 118.730 178.485 ;
        RECT 118.995 177.835 119.280 178.975 ;
        RECT 119.470 178.015 119.750 180.205 ;
        RECT 120.395 179.660 120.685 180.385 ;
        RECT 120.855 179.840 126.200 180.385 ;
        RECT 126.400 179.995 126.730 180.385 ;
        RECT 122.440 179.010 122.780 179.840 ;
        RECT 126.900 179.825 127.125 180.205 ;
        RECT 120.395 177.835 120.685 179.000 ;
        RECT 124.260 178.270 124.610 179.520 ;
        RECT 126.385 179.145 126.625 179.795 ;
        RECT 126.795 179.645 127.125 179.825 ;
        RECT 126.795 178.975 126.970 179.645 ;
        RECT 127.325 179.475 127.555 180.095 ;
        RECT 127.735 179.655 128.035 180.385 ;
        RECT 128.235 179.575 128.475 180.385 ;
        RECT 128.645 179.575 128.975 180.215 ;
        RECT 129.145 179.575 129.415 180.385 ;
        RECT 129.595 179.615 132.185 180.385 ;
        RECT 132.355 179.645 132.940 180.215 ;
        RECT 133.190 179.815 133.520 180.160 ;
        RECT 133.735 179.985 134.110 180.385 ;
        RECT 134.290 179.815 134.585 180.160 ;
        RECT 133.190 179.645 134.585 179.815 ;
        RECT 134.755 179.645 135.425 180.385 ;
        RECT 127.140 179.145 127.555 179.475 ;
        RECT 127.735 179.145 128.030 179.475 ;
        RECT 128.215 179.145 128.565 179.395 ;
        RECT 128.735 178.975 128.905 179.575 ;
        RECT 129.075 179.145 129.425 179.395 ;
        RECT 129.595 179.095 130.805 179.615 ;
        RECT 126.385 178.785 126.970 178.975 ;
        RECT 120.855 177.835 126.200 178.270 ;
        RECT 126.385 178.015 126.660 178.785 ;
        RECT 127.140 178.615 128.035 178.945 ;
        RECT 126.830 178.445 128.035 178.615 ;
        RECT 126.830 178.015 127.160 178.445 ;
        RECT 127.330 177.835 127.525 178.275 ;
        RECT 127.705 178.015 128.035 178.445 ;
        RECT 128.225 178.805 128.905 178.975 ;
        RECT 128.225 178.020 128.555 178.805 ;
        RECT 129.085 177.835 129.415 178.975 ;
        RECT 130.975 178.925 132.185 179.445 ;
        RECT 132.355 179.145 132.600 179.475 ;
        RECT 132.770 178.975 132.940 179.645 ;
        RECT 133.110 179.145 133.510 179.475 ;
        RECT 133.680 179.145 133.970 179.475 ;
        RECT 129.595 177.835 132.185 178.925 ;
        RECT 132.355 178.805 133.565 178.975 ;
        RECT 132.355 178.005 132.645 178.805 ;
        RECT 132.815 177.835 133.050 178.635 ;
        RECT 133.235 178.175 133.565 178.805 ;
        RECT 133.735 178.400 133.970 179.145 ;
        RECT 134.160 179.145 134.500 179.475 ;
        RECT 134.670 179.145 135.005 179.475 ;
        RECT 134.160 178.400 134.430 179.145 ;
        RECT 135.175 178.975 135.345 179.475 ;
        RECT 135.595 179.400 135.865 180.215 ;
        RECT 134.600 178.805 135.345 178.975 ;
        RECT 134.600 178.175 134.770 178.805 ;
        RECT 133.235 178.005 134.770 178.175 ;
        RECT 134.940 177.835 135.345 178.635 ;
        RECT 135.515 178.005 135.865 179.400 ;
        RECT 136.035 179.925 136.595 180.215 ;
        RECT 136.765 179.925 137.015 180.385 ;
        RECT 136.035 178.555 136.285 179.925 ;
        RECT 137.635 179.755 137.965 180.115 ;
        RECT 136.575 179.565 137.965 179.755 ;
        RECT 138.355 179.575 138.595 180.385 ;
        RECT 138.765 179.575 139.095 180.215 ;
        RECT 139.265 179.575 139.535 180.385 ;
        RECT 139.715 179.840 145.060 180.385 ;
        RECT 136.575 179.475 136.745 179.565 ;
        RECT 136.455 179.145 136.745 179.475 ;
        RECT 136.915 179.145 137.255 179.395 ;
        RECT 137.475 179.145 138.150 179.395 ;
        RECT 138.335 179.145 138.685 179.395 ;
        RECT 136.575 178.895 136.745 179.145 ;
        RECT 136.575 178.725 137.515 178.895 ;
        RECT 137.885 178.785 138.150 179.145 ;
        RECT 138.855 178.975 139.025 179.575 ;
        RECT 139.195 179.145 139.545 179.395 ;
        RECT 141.300 179.010 141.640 179.840 ;
        RECT 145.695 179.635 146.905 180.385 ;
        RECT 138.345 178.805 139.025 178.975 ;
        RECT 136.035 178.005 136.495 178.555 ;
        RECT 136.685 177.835 137.015 178.555 ;
        RECT 137.215 178.175 137.515 178.725 ;
        RECT 137.685 177.835 137.965 178.505 ;
        RECT 138.345 178.020 138.675 178.805 ;
        RECT 139.205 177.835 139.535 178.975 ;
        RECT 143.120 178.270 143.470 179.520 ;
        RECT 145.695 178.925 146.215 179.465 ;
        RECT 146.385 179.095 146.905 179.635 ;
        RECT 139.715 177.835 145.060 178.270 ;
        RECT 145.695 177.835 146.905 178.925 ;
        RECT 17.270 177.665 146.990 177.835 ;
        RECT 17.355 176.575 18.565 177.665 ;
        RECT 18.735 176.575 22.245 177.665 ;
        RECT 22.415 176.575 23.625 177.665 ;
        RECT 17.355 175.865 17.875 176.405 ;
        RECT 18.045 176.035 18.565 176.575 ;
        RECT 18.735 175.885 20.385 176.405 ;
        RECT 20.555 176.055 22.245 176.575 ;
        RECT 17.355 175.115 18.565 175.865 ;
        RECT 18.735 175.115 22.245 175.885 ;
        RECT 22.415 175.865 22.935 176.405 ;
        RECT 23.105 176.035 23.625 176.575 ;
        RECT 23.855 176.525 24.065 177.665 ;
        RECT 24.235 176.515 24.565 177.495 ;
        RECT 24.735 176.525 24.965 177.665 ;
        RECT 25.635 176.945 26.095 177.495 ;
        RECT 26.285 176.945 26.615 177.665 ;
        RECT 22.415 175.115 23.625 175.865 ;
        RECT 23.855 175.115 24.065 175.935 ;
        RECT 24.235 175.915 24.485 176.515 ;
        RECT 24.655 176.105 24.985 176.355 ;
        RECT 24.235 175.285 24.565 175.915 ;
        RECT 24.735 175.115 24.965 175.935 ;
        RECT 25.635 175.575 25.885 176.945 ;
        RECT 26.815 176.775 27.115 177.325 ;
        RECT 27.285 176.995 27.565 177.665 ;
        RECT 26.175 176.605 27.115 176.775 ;
        RECT 26.175 176.355 26.345 176.605 ;
        RECT 27.485 176.355 27.750 176.715 ;
        RECT 27.935 176.575 29.605 177.665 ;
        RECT 26.055 176.025 26.345 176.355 ;
        RECT 26.515 176.105 26.855 176.355 ;
        RECT 27.075 176.105 27.750 176.355 ;
        RECT 26.175 175.935 26.345 176.025 ;
        RECT 26.175 175.745 27.565 175.935 ;
        RECT 25.635 175.285 26.195 175.575 ;
        RECT 26.365 175.115 26.615 175.575 ;
        RECT 27.235 175.385 27.565 175.745 ;
        RECT 27.935 175.885 28.685 176.405 ;
        RECT 28.855 176.055 29.605 176.575 ;
        RECT 30.235 176.500 30.525 177.665 ;
        RECT 30.700 177.275 31.035 177.495 ;
        RECT 32.040 177.285 32.395 177.665 ;
        RECT 30.700 176.655 30.955 177.275 ;
        RECT 31.205 177.115 31.435 177.155 ;
        RECT 32.565 177.115 32.815 177.495 ;
        RECT 31.205 176.915 32.815 177.115 ;
        RECT 31.205 176.825 31.390 176.915 ;
        RECT 31.980 176.905 32.815 176.915 ;
        RECT 33.065 176.885 33.315 177.665 ;
        RECT 33.485 176.815 33.745 177.495 ;
        RECT 31.545 176.715 31.875 176.745 ;
        RECT 31.545 176.655 33.345 176.715 ;
        RECT 30.700 176.545 33.405 176.655 ;
        RECT 30.700 176.485 31.875 176.545 ;
        RECT 33.205 176.510 33.405 176.545 ;
        RECT 30.695 176.105 31.185 176.305 ;
        RECT 31.375 176.105 31.850 176.315 ;
        RECT 27.935 175.115 29.605 175.885 ;
        RECT 30.235 175.115 30.525 175.840 ;
        RECT 30.700 175.115 31.155 175.880 ;
        RECT 31.630 175.705 31.850 176.105 ;
        RECT 32.095 176.105 32.425 176.315 ;
        RECT 32.095 175.705 32.305 176.105 ;
        RECT 32.595 176.070 33.005 176.375 ;
        RECT 33.235 175.935 33.405 176.510 ;
        RECT 33.135 175.815 33.405 175.935 ;
        RECT 32.560 175.770 33.405 175.815 ;
        RECT 32.560 175.645 33.315 175.770 ;
        RECT 32.560 175.495 32.730 175.645 ;
        RECT 33.575 175.615 33.745 176.815 ;
        RECT 33.915 176.485 34.235 177.665 ;
        RECT 34.405 176.645 34.605 177.435 ;
        RECT 34.795 177.075 35.295 177.495 ;
        RECT 35.785 177.205 35.995 177.665 ;
        RECT 34.795 176.865 35.635 177.075 ;
        RECT 34.405 176.475 34.725 176.645 ;
        RECT 33.915 176.105 34.375 176.305 ;
        RECT 34.545 176.275 34.725 176.475 ;
        RECT 34.895 176.445 35.295 176.695 ;
        RECT 34.545 176.105 34.910 176.275 ;
        RECT 35.125 176.025 35.295 176.445 ;
        RECT 31.430 175.285 32.730 175.495 ;
        RECT 32.985 175.115 33.315 175.475 ;
        RECT 33.485 175.285 33.745 175.615 ;
        RECT 33.915 175.855 34.945 175.895 ;
        RECT 35.465 175.855 35.635 176.865 ;
        RECT 33.915 175.725 35.115 175.855 ;
        RECT 33.915 175.310 34.255 175.725 ;
        RECT 34.425 175.115 34.595 175.555 ;
        RECT 34.785 175.505 35.115 175.725 ;
        RECT 35.285 175.675 35.635 175.855 ;
        RECT 35.805 175.695 36.045 177.020 ;
        RECT 36.215 176.525 36.475 177.665 ;
        RECT 36.645 176.515 36.975 177.495 ;
        RECT 37.145 176.525 37.425 177.665 ;
        RECT 37.595 177.230 42.940 177.665 ;
        RECT 36.235 176.105 36.570 176.355 ;
        RECT 36.740 175.915 36.910 176.515 ;
        RECT 37.080 176.085 37.415 176.355 ;
        RECT 34.785 175.325 36.045 175.505 ;
        RECT 36.215 175.285 36.910 175.915 ;
        RECT 37.115 175.115 37.425 175.915 ;
        RECT 39.180 175.660 39.520 176.490 ;
        RECT 41.000 175.980 41.350 177.230 ;
        RECT 43.580 177.155 45.235 177.445 ;
        RECT 43.580 176.815 45.170 176.985 ;
        RECT 45.405 176.865 45.685 177.665 ;
        RECT 43.580 176.525 43.900 176.815 ;
        RECT 45.000 176.695 45.170 176.815 ;
        RECT 43.580 175.785 43.930 176.355 ;
        RECT 44.100 176.025 44.810 176.645 ;
        RECT 45.000 176.525 45.725 176.695 ;
        RECT 45.895 176.525 46.165 177.495 ;
        RECT 46.335 177.110 46.940 177.665 ;
        RECT 47.115 177.155 47.595 177.495 ;
        RECT 47.765 177.120 48.020 177.665 ;
        RECT 46.335 177.010 46.950 177.110 ;
        RECT 46.765 176.985 46.950 177.010 ;
        RECT 45.555 176.355 45.725 176.525 ;
        RECT 44.980 176.025 45.385 176.355 ;
        RECT 45.555 176.025 45.825 176.355 ;
        RECT 45.555 175.855 45.725 176.025 ;
        RECT 44.115 175.685 45.725 175.855 ;
        RECT 45.995 175.790 46.165 176.525 ;
        RECT 46.335 176.390 46.595 176.840 ;
        RECT 46.765 176.740 47.095 176.985 ;
        RECT 47.265 176.665 48.020 176.915 ;
        RECT 48.190 176.795 48.465 177.495 ;
        RECT 47.250 176.630 48.020 176.665 ;
        RECT 47.235 176.620 48.020 176.630 ;
        RECT 47.230 176.605 48.125 176.620 ;
        RECT 47.210 176.590 48.125 176.605 ;
        RECT 47.190 176.580 48.125 176.590 ;
        RECT 47.165 176.570 48.125 176.580 ;
        RECT 47.095 176.540 48.125 176.570 ;
        RECT 47.075 176.510 48.125 176.540 ;
        RECT 47.055 176.480 48.125 176.510 ;
        RECT 47.025 176.455 48.125 176.480 ;
        RECT 46.990 176.420 48.125 176.455 ;
        RECT 46.960 176.415 48.125 176.420 ;
        RECT 46.960 176.410 47.350 176.415 ;
        RECT 46.960 176.400 47.325 176.410 ;
        RECT 46.960 176.395 47.310 176.400 ;
        RECT 46.960 176.390 47.295 176.395 ;
        RECT 46.335 176.385 47.295 176.390 ;
        RECT 46.335 176.375 47.285 176.385 ;
        RECT 46.335 176.370 47.275 176.375 ;
        RECT 46.335 176.360 47.265 176.370 ;
        RECT 46.335 176.350 47.260 176.360 ;
        RECT 46.335 176.345 47.255 176.350 ;
        RECT 46.335 176.330 47.245 176.345 ;
        RECT 46.335 176.315 47.240 176.330 ;
        RECT 46.335 176.290 47.230 176.315 ;
        RECT 46.335 176.220 47.225 176.290 ;
        RECT 37.595 175.115 42.940 175.660 ;
        RECT 43.585 175.115 43.915 175.615 ;
        RECT 44.115 175.335 44.285 175.685 ;
        RECT 44.485 175.115 44.815 175.515 ;
        RECT 44.985 175.335 45.155 175.685 ;
        RECT 45.325 175.115 45.705 175.515 ;
        RECT 45.895 175.445 46.165 175.790 ;
        RECT 46.335 175.665 46.885 176.050 ;
        RECT 47.055 175.495 47.225 176.220 ;
        RECT 46.335 175.325 47.225 175.495 ;
        RECT 47.395 175.820 47.725 176.245 ;
        RECT 47.895 176.020 48.125 176.415 ;
        RECT 47.395 175.335 47.615 175.820 ;
        RECT 48.295 175.765 48.465 176.795 ;
        RECT 48.675 176.525 48.905 177.665 ;
        RECT 49.075 176.515 49.405 177.495 ;
        RECT 49.575 176.525 49.785 177.665 ;
        RECT 50.015 176.575 52.605 177.665 ;
        RECT 48.655 176.105 48.985 176.355 ;
        RECT 47.785 175.115 48.035 175.655 ;
        RECT 48.205 175.285 48.465 175.765 ;
        RECT 48.675 175.115 48.905 175.935 ;
        RECT 49.155 175.915 49.405 176.515 ;
        RECT 49.075 175.285 49.405 175.915 ;
        RECT 49.575 175.115 49.785 175.935 ;
        RECT 50.015 175.885 51.225 176.405 ;
        RECT 51.395 176.055 52.605 176.575 ;
        RECT 53.275 176.525 53.505 177.665 ;
        RECT 53.675 176.515 54.005 177.495 ;
        RECT 54.175 176.525 54.385 177.665 ;
        RECT 54.615 176.575 55.825 177.665 ;
        RECT 53.255 176.105 53.585 176.355 ;
        RECT 50.015 175.115 52.605 175.885 ;
        RECT 53.275 175.115 53.505 175.935 ;
        RECT 53.755 175.915 54.005 176.515 ;
        RECT 53.675 175.285 54.005 175.915 ;
        RECT 54.175 175.115 54.385 175.935 ;
        RECT 54.615 175.865 55.135 176.405 ;
        RECT 55.305 176.035 55.825 176.575 ;
        RECT 55.995 176.500 56.285 177.665 ;
        RECT 56.925 176.525 57.255 177.665 ;
        RECT 57.785 176.695 58.115 177.480 ;
        RECT 58.385 176.995 58.555 177.495 ;
        RECT 58.725 177.165 59.055 177.665 ;
        RECT 58.385 176.825 59.050 176.995 ;
        RECT 57.435 176.525 58.115 176.695 ;
        RECT 56.915 176.105 57.265 176.355 ;
        RECT 57.435 175.925 57.605 176.525 ;
        RECT 57.775 176.105 58.125 176.355 ;
        RECT 58.300 176.005 58.650 176.655 ;
        RECT 54.615 175.115 55.825 175.865 ;
        RECT 55.995 175.115 56.285 175.840 ;
        RECT 56.925 175.115 57.195 175.925 ;
        RECT 57.365 175.285 57.695 175.925 ;
        RECT 57.865 175.115 58.105 175.925 ;
        RECT 58.820 175.835 59.050 176.825 ;
        RECT 58.385 175.665 59.050 175.835 ;
        RECT 58.385 175.375 58.555 175.665 ;
        RECT 58.725 175.115 59.055 175.495 ;
        RECT 59.225 175.375 59.410 177.495 ;
        RECT 59.650 177.205 59.915 177.665 ;
        RECT 60.085 177.070 60.335 177.495 ;
        RECT 60.545 177.220 61.650 177.390 ;
        RECT 60.030 176.940 60.335 177.070 ;
        RECT 59.580 175.745 59.860 176.695 ;
        RECT 60.030 175.835 60.200 176.940 ;
        RECT 60.370 176.155 60.610 176.750 ;
        RECT 60.780 176.685 61.310 177.050 ;
        RECT 60.780 175.985 60.950 176.685 ;
        RECT 61.480 176.605 61.650 177.220 ;
        RECT 61.820 176.865 61.990 177.665 ;
        RECT 62.160 177.165 62.410 177.495 ;
        RECT 62.635 177.195 63.520 177.365 ;
        RECT 61.480 176.515 61.990 176.605 ;
        RECT 60.030 175.705 60.255 175.835 ;
        RECT 60.425 175.765 60.950 175.985 ;
        RECT 61.120 176.345 61.990 176.515 ;
        RECT 59.665 175.115 59.915 175.575 ;
        RECT 60.085 175.565 60.255 175.705 ;
        RECT 61.120 175.565 61.290 176.345 ;
        RECT 61.820 176.275 61.990 176.345 ;
        RECT 61.500 176.095 61.700 176.125 ;
        RECT 62.160 176.095 62.330 177.165 ;
        RECT 62.500 176.275 62.690 176.995 ;
        RECT 61.500 175.795 62.330 176.095 ;
        RECT 62.860 176.065 63.180 177.025 ;
        RECT 60.085 175.395 60.420 175.565 ;
        RECT 60.615 175.395 61.290 175.565 ;
        RECT 61.610 175.115 61.980 175.615 ;
        RECT 62.160 175.565 62.330 175.795 ;
        RECT 62.715 175.735 63.180 176.065 ;
        RECT 63.350 176.355 63.520 177.195 ;
        RECT 63.700 177.165 64.015 177.665 ;
        RECT 64.245 176.935 64.585 177.495 ;
        RECT 63.690 176.560 64.585 176.935 ;
        RECT 64.755 176.655 64.925 177.665 ;
        RECT 64.395 176.355 64.585 176.560 ;
        RECT 65.095 176.605 65.425 177.450 ;
        RECT 65.715 176.605 66.045 177.450 ;
        RECT 66.215 176.655 66.385 177.665 ;
        RECT 66.555 176.935 66.895 177.495 ;
        RECT 67.125 177.165 67.440 177.665 ;
        RECT 67.620 177.195 68.505 177.365 ;
        RECT 65.095 176.525 65.485 176.605 ;
        RECT 65.270 176.475 65.485 176.525 ;
        RECT 63.350 176.025 64.225 176.355 ;
        RECT 64.395 176.025 65.145 176.355 ;
        RECT 63.350 175.565 63.520 176.025 ;
        RECT 64.395 175.855 64.595 176.025 ;
        RECT 65.315 175.895 65.485 176.475 ;
        RECT 65.260 175.855 65.485 175.895 ;
        RECT 62.160 175.395 62.565 175.565 ;
        RECT 62.735 175.395 63.520 175.565 ;
        RECT 63.795 175.115 64.005 175.645 ;
        RECT 64.265 175.330 64.595 175.855 ;
        RECT 65.105 175.770 65.485 175.855 ;
        RECT 65.655 176.525 66.045 176.605 ;
        RECT 66.555 176.560 67.450 176.935 ;
        RECT 65.655 176.475 65.870 176.525 ;
        RECT 65.655 175.895 65.825 176.475 ;
        RECT 66.555 176.355 66.745 176.560 ;
        RECT 67.620 176.355 67.790 177.195 ;
        RECT 68.730 177.165 68.980 177.495 ;
        RECT 65.995 176.025 66.745 176.355 ;
        RECT 66.915 176.025 67.790 176.355 ;
        RECT 65.655 175.855 65.880 175.895 ;
        RECT 66.545 175.855 66.745 176.025 ;
        RECT 65.655 175.770 66.035 175.855 ;
        RECT 64.765 175.115 64.935 175.725 ;
        RECT 65.105 175.335 65.435 175.770 ;
        RECT 65.705 175.335 66.035 175.770 ;
        RECT 66.205 175.115 66.375 175.725 ;
        RECT 66.545 175.330 66.875 175.855 ;
        RECT 67.135 175.115 67.345 175.645 ;
        RECT 67.620 175.565 67.790 176.025 ;
        RECT 67.960 176.065 68.280 177.025 ;
        RECT 68.450 176.275 68.640 176.995 ;
        RECT 68.810 176.095 68.980 177.165 ;
        RECT 69.150 176.865 69.320 177.665 ;
        RECT 69.490 177.220 70.595 177.390 ;
        RECT 69.490 176.605 69.660 177.220 ;
        RECT 70.805 177.070 71.055 177.495 ;
        RECT 71.225 177.205 71.490 177.665 ;
        RECT 69.830 176.685 70.360 177.050 ;
        RECT 70.805 176.940 71.110 177.070 ;
        RECT 69.150 176.515 69.660 176.605 ;
        RECT 69.150 176.345 70.020 176.515 ;
        RECT 69.150 176.275 69.320 176.345 ;
        RECT 69.440 176.095 69.640 176.125 ;
        RECT 67.960 175.735 68.425 176.065 ;
        RECT 68.810 175.795 69.640 176.095 ;
        RECT 68.810 175.565 68.980 175.795 ;
        RECT 67.620 175.395 68.405 175.565 ;
        RECT 68.575 175.395 68.980 175.565 ;
        RECT 69.160 175.115 69.530 175.615 ;
        RECT 69.850 175.565 70.020 176.345 ;
        RECT 70.190 175.985 70.360 176.685 ;
        RECT 70.530 176.155 70.770 176.750 ;
        RECT 70.190 175.765 70.715 175.985 ;
        RECT 70.940 175.835 71.110 176.940 ;
        RECT 70.885 175.705 71.110 175.835 ;
        RECT 71.280 175.745 71.560 176.695 ;
        RECT 70.885 175.565 71.055 175.705 ;
        RECT 69.850 175.395 70.525 175.565 ;
        RECT 70.720 175.395 71.055 175.565 ;
        RECT 71.225 175.115 71.475 175.575 ;
        RECT 71.730 175.375 71.915 177.495 ;
        RECT 72.085 177.165 72.415 177.665 ;
        RECT 72.585 176.995 72.755 177.495 ;
        RECT 73.015 177.230 78.360 177.665 ;
        RECT 72.090 176.825 72.755 176.995 ;
        RECT 72.090 175.835 72.320 176.825 ;
        RECT 72.490 176.005 72.840 176.655 ;
        RECT 72.090 175.665 72.755 175.835 ;
        RECT 72.085 175.115 72.415 175.495 ;
        RECT 72.585 175.375 72.755 175.665 ;
        RECT 74.600 175.660 74.940 176.490 ;
        RECT 76.420 175.980 76.770 177.230 ;
        RECT 78.535 176.575 81.125 177.665 ;
        RECT 78.535 175.885 79.745 176.405 ;
        RECT 79.915 176.055 81.125 176.575 ;
        RECT 81.755 176.500 82.045 177.665 ;
        RECT 82.215 176.575 83.885 177.665 ;
        RECT 84.630 177.035 84.915 177.495 ;
        RECT 85.085 177.205 85.355 177.665 ;
        RECT 84.630 176.815 85.585 177.035 ;
        RECT 82.215 175.885 82.965 176.405 ;
        RECT 83.135 176.055 83.885 176.575 ;
        RECT 84.515 176.085 85.205 176.645 ;
        RECT 85.375 175.915 85.585 176.815 ;
        RECT 73.015 175.115 78.360 175.660 ;
        RECT 78.535 175.115 81.125 175.885 ;
        RECT 81.755 175.115 82.045 175.840 ;
        RECT 82.215 175.115 83.885 175.885 ;
        RECT 84.630 175.745 85.585 175.915 ;
        RECT 85.755 176.645 86.155 177.495 ;
        RECT 86.345 177.035 86.625 177.495 ;
        RECT 87.145 177.205 87.470 177.665 ;
        RECT 86.345 176.815 87.470 177.035 ;
        RECT 85.755 176.085 86.850 176.645 ;
        RECT 87.020 176.355 87.470 176.815 ;
        RECT 87.640 176.525 88.025 177.495 ;
        RECT 88.195 176.575 91.705 177.665 ;
        RECT 91.875 176.575 93.085 177.665 ;
        RECT 93.345 176.995 93.515 177.495 ;
        RECT 93.685 177.165 94.015 177.665 ;
        RECT 93.345 176.825 94.010 176.995 ;
        RECT 84.630 175.285 84.915 175.745 ;
        RECT 85.085 175.115 85.355 175.575 ;
        RECT 85.755 175.285 86.155 176.085 ;
        RECT 87.020 176.025 87.575 176.355 ;
        RECT 87.020 175.915 87.470 176.025 ;
        RECT 86.345 175.745 87.470 175.915 ;
        RECT 87.745 175.855 88.025 176.525 ;
        RECT 86.345 175.285 86.625 175.745 ;
        RECT 87.145 175.115 87.470 175.575 ;
        RECT 87.640 175.285 88.025 175.855 ;
        RECT 88.195 175.885 89.845 176.405 ;
        RECT 90.015 176.055 91.705 176.575 ;
        RECT 88.195 175.115 91.705 175.885 ;
        RECT 91.875 175.865 92.395 176.405 ;
        RECT 92.565 176.035 93.085 176.575 ;
        RECT 93.260 176.005 93.610 176.655 ;
        RECT 91.875 175.115 93.085 175.865 ;
        RECT 93.780 175.835 94.010 176.825 ;
        RECT 93.345 175.665 94.010 175.835 ;
        RECT 93.345 175.375 93.515 175.665 ;
        RECT 93.685 175.115 94.015 175.495 ;
        RECT 94.185 175.375 94.370 177.495 ;
        RECT 94.610 177.205 94.875 177.665 ;
        RECT 95.045 177.070 95.295 177.495 ;
        RECT 95.505 177.220 96.610 177.390 ;
        RECT 94.990 176.940 95.295 177.070 ;
        RECT 94.540 175.745 94.820 176.695 ;
        RECT 94.990 175.835 95.160 176.940 ;
        RECT 95.330 176.155 95.570 176.750 ;
        RECT 95.740 176.685 96.270 177.050 ;
        RECT 95.740 175.985 95.910 176.685 ;
        RECT 96.440 176.605 96.610 177.220 ;
        RECT 96.780 176.865 96.950 177.665 ;
        RECT 97.120 177.165 97.370 177.495 ;
        RECT 97.595 177.195 98.480 177.365 ;
        RECT 96.440 176.515 96.950 176.605 ;
        RECT 94.990 175.705 95.215 175.835 ;
        RECT 95.385 175.765 95.910 175.985 ;
        RECT 96.080 176.345 96.950 176.515 ;
        RECT 94.625 175.115 94.875 175.575 ;
        RECT 95.045 175.565 95.215 175.705 ;
        RECT 96.080 175.565 96.250 176.345 ;
        RECT 96.780 176.275 96.950 176.345 ;
        RECT 96.460 176.095 96.660 176.125 ;
        RECT 97.120 176.095 97.290 177.165 ;
        RECT 97.460 176.275 97.650 176.995 ;
        RECT 96.460 175.795 97.290 176.095 ;
        RECT 97.820 176.065 98.140 177.025 ;
        RECT 95.045 175.395 95.380 175.565 ;
        RECT 95.575 175.395 96.250 175.565 ;
        RECT 96.570 175.115 96.940 175.615 ;
        RECT 97.120 175.565 97.290 175.795 ;
        RECT 97.675 175.735 98.140 176.065 ;
        RECT 98.310 176.355 98.480 177.195 ;
        RECT 98.660 177.165 98.975 177.665 ;
        RECT 99.205 176.935 99.545 177.495 ;
        RECT 98.650 176.560 99.545 176.935 ;
        RECT 99.715 176.655 99.885 177.665 ;
        RECT 99.355 176.355 99.545 176.560 ;
        RECT 100.055 176.605 100.385 177.450 ;
        RECT 100.055 176.525 100.445 176.605 ;
        RECT 100.230 176.475 100.445 176.525 ;
        RECT 98.310 176.025 99.185 176.355 ;
        RECT 99.355 176.025 100.105 176.355 ;
        RECT 98.310 175.565 98.480 176.025 ;
        RECT 99.355 175.855 99.555 176.025 ;
        RECT 100.275 175.895 100.445 176.475 ;
        RECT 100.220 175.855 100.445 175.895 ;
        RECT 97.120 175.395 97.525 175.565 ;
        RECT 97.695 175.395 98.480 175.565 ;
        RECT 98.755 175.115 98.965 175.645 ;
        RECT 99.225 175.330 99.555 175.855 ;
        RECT 100.065 175.770 100.445 175.855 ;
        RECT 100.620 176.525 100.955 177.495 ;
        RECT 101.125 176.525 101.295 177.665 ;
        RECT 101.465 177.325 103.495 177.495 ;
        RECT 100.620 175.855 100.790 176.525 ;
        RECT 101.465 176.355 101.635 177.325 ;
        RECT 100.960 176.025 101.215 176.355 ;
        RECT 101.440 176.025 101.635 176.355 ;
        RECT 101.805 176.985 102.930 177.155 ;
        RECT 101.045 175.855 101.215 176.025 ;
        RECT 101.805 175.855 101.975 176.985 ;
        RECT 99.725 175.115 99.895 175.725 ;
        RECT 100.065 175.335 100.395 175.770 ;
        RECT 100.620 175.285 100.875 175.855 ;
        RECT 101.045 175.685 101.975 175.855 ;
        RECT 102.145 176.645 103.155 176.815 ;
        RECT 102.145 175.845 102.315 176.645 ;
        RECT 102.520 175.965 102.795 176.445 ;
        RECT 102.515 175.795 102.795 175.965 ;
        RECT 101.800 175.650 101.975 175.685 ;
        RECT 101.045 175.115 101.375 175.515 ;
        RECT 101.800 175.285 102.330 175.650 ;
        RECT 102.520 175.285 102.795 175.795 ;
        RECT 102.965 175.285 103.155 176.645 ;
        RECT 103.325 176.660 103.495 177.325 ;
        RECT 103.665 176.905 103.835 177.665 ;
        RECT 104.070 176.905 104.585 177.315 ;
        RECT 103.325 176.470 104.075 176.660 ;
        RECT 104.245 176.095 104.585 176.905 ;
        RECT 105.685 177.055 106.015 177.485 ;
        RECT 106.195 177.225 106.390 177.665 ;
        RECT 106.560 177.055 106.890 177.485 ;
        RECT 105.685 176.885 106.890 177.055 ;
        RECT 105.685 176.555 106.580 176.885 ;
        RECT 107.060 176.715 107.335 177.485 ;
        RECT 106.750 176.525 107.335 176.715 ;
        RECT 103.355 175.925 104.585 176.095 ;
        RECT 105.690 176.025 105.985 176.355 ;
        RECT 106.165 176.025 106.580 176.355 ;
        RECT 103.335 175.115 103.845 175.650 ;
        RECT 104.065 175.320 104.310 175.925 ;
        RECT 105.685 175.115 105.985 175.845 ;
        RECT 106.165 175.405 106.395 176.025 ;
        RECT 106.750 175.855 106.925 176.525 ;
        RECT 107.515 176.500 107.805 177.665 ;
        RECT 108.015 176.525 108.245 177.665 ;
        RECT 108.415 176.515 108.745 177.495 ;
        RECT 108.915 176.525 109.125 177.665 ;
        RECT 109.355 176.525 109.615 177.495 ;
        RECT 109.785 177.240 110.170 177.665 ;
        RECT 110.340 177.070 110.595 177.495 ;
        RECT 109.785 176.875 110.595 177.070 ;
        RECT 106.595 175.675 106.925 175.855 ;
        RECT 107.095 175.705 107.335 176.355 ;
        RECT 107.995 176.105 108.325 176.355 ;
        RECT 106.595 175.295 106.820 175.675 ;
        RECT 106.990 175.115 107.320 175.505 ;
        RECT 107.515 175.115 107.805 175.840 ;
        RECT 108.015 175.115 108.245 175.935 ;
        RECT 108.495 175.915 108.745 176.515 ;
        RECT 108.415 175.285 108.745 175.915 ;
        RECT 108.915 175.115 109.125 175.935 ;
        RECT 109.355 175.855 109.540 176.525 ;
        RECT 109.785 176.355 110.135 176.875 ;
        RECT 110.785 176.705 111.030 177.495 ;
        RECT 111.200 177.240 111.585 177.665 ;
        RECT 111.755 177.070 112.030 177.495 ;
        RECT 109.710 176.025 110.135 176.355 ;
        RECT 110.305 176.525 111.030 176.705 ;
        RECT 111.200 176.875 112.030 177.070 ;
        RECT 110.305 176.025 110.955 176.525 ;
        RECT 111.200 176.355 111.550 176.875 ;
        RECT 112.200 176.705 112.625 177.495 ;
        RECT 112.795 177.240 113.180 177.665 ;
        RECT 113.350 177.070 113.785 177.495 ;
        RECT 111.125 176.025 111.550 176.355 ;
        RECT 111.720 176.525 112.625 176.705 ;
        RECT 112.795 176.900 113.785 177.070 ;
        RECT 111.720 176.025 112.550 176.525 ;
        RECT 112.795 176.355 113.130 176.900 ;
        RECT 112.720 176.025 113.130 176.355 ;
        RECT 113.300 176.025 113.785 176.730 ;
        RECT 113.955 176.525 114.230 177.495 ;
        RECT 114.440 176.865 114.720 177.665 ;
        RECT 114.890 177.155 116.940 177.445 ;
        RECT 114.890 176.815 116.520 176.985 ;
        RECT 114.890 176.695 115.060 176.815 ;
        RECT 114.400 176.525 115.060 176.695 ;
        RECT 109.785 175.855 110.135 176.025 ;
        RECT 110.785 175.855 110.955 176.025 ;
        RECT 111.200 175.855 111.550 176.025 ;
        RECT 112.200 175.855 112.550 176.025 ;
        RECT 112.795 175.855 113.130 176.025 ;
        RECT 109.355 175.285 109.615 175.855 ;
        RECT 109.785 175.685 110.595 175.855 ;
        RECT 109.785 175.115 110.170 175.515 ;
        RECT 110.340 175.285 110.595 175.685 ;
        RECT 110.785 175.285 111.030 175.855 ;
        RECT 111.200 175.685 112.010 175.855 ;
        RECT 111.200 175.115 111.585 175.515 ;
        RECT 111.755 175.285 112.010 175.685 ;
        RECT 112.200 175.285 112.625 175.855 ;
        RECT 112.795 175.685 113.785 175.855 ;
        RECT 112.795 175.115 113.180 175.515 ;
        RECT 113.350 175.285 113.785 175.685 ;
        RECT 113.955 175.790 114.125 176.525 ;
        RECT 114.400 176.355 114.570 176.525 ;
        RECT 114.295 176.025 114.570 176.355 ;
        RECT 114.740 176.025 115.120 176.355 ;
        RECT 115.290 176.025 116.030 176.645 ;
        RECT 116.200 176.525 116.520 176.815 ;
        RECT 116.715 176.355 116.955 176.950 ;
        RECT 117.125 176.590 117.465 177.665 ;
        RECT 117.835 176.995 118.115 177.665 ;
        RECT 118.285 176.775 118.585 177.325 ;
        RECT 118.785 176.945 119.115 177.665 ;
        RECT 119.305 176.945 119.765 177.495 ;
        RECT 117.650 176.355 117.915 176.715 ;
        RECT 118.285 176.605 119.225 176.775 ;
        RECT 119.055 176.355 119.225 176.605 ;
        RECT 116.300 176.025 116.955 176.355 ;
        RECT 114.400 175.855 114.570 176.025 ;
        RECT 113.955 175.445 114.230 175.790 ;
        RECT 114.400 175.685 115.985 175.855 ;
        RECT 114.420 175.115 114.800 175.515 ;
        RECT 114.970 175.335 115.140 175.685 ;
        RECT 115.310 175.115 115.640 175.515 ;
        RECT 115.815 175.335 115.985 175.685 ;
        RECT 116.185 175.115 116.515 175.615 ;
        RECT 116.710 175.335 116.955 176.025 ;
        RECT 117.125 175.785 117.465 176.355 ;
        RECT 117.650 176.105 118.325 176.355 ;
        RECT 118.545 176.105 118.885 176.355 ;
        RECT 119.055 176.025 119.345 176.355 ;
        RECT 119.055 175.935 119.225 176.025 ;
        RECT 117.835 175.745 119.225 175.935 ;
        RECT 117.125 175.115 117.465 175.615 ;
        RECT 117.835 175.385 118.165 175.745 ;
        RECT 119.515 175.575 119.765 176.945 ;
        RECT 119.935 176.525 120.215 177.665 ;
        RECT 120.385 176.515 120.715 177.495 ;
        RECT 120.885 176.525 121.145 177.665 ;
        RECT 121.315 176.575 122.525 177.665 ;
        RECT 119.945 176.085 120.280 176.355 ;
        RECT 120.450 175.915 120.620 176.515 ;
        RECT 120.790 176.105 121.125 176.355 ;
        RECT 118.785 175.115 119.035 175.575 ;
        RECT 119.205 175.285 119.765 175.575 ;
        RECT 119.935 175.115 120.245 175.915 ;
        RECT 120.450 175.285 121.145 175.915 ;
        RECT 121.315 175.865 121.835 176.405 ;
        RECT 122.005 176.035 122.525 176.575 ;
        RECT 122.695 176.525 122.970 177.495 ;
        RECT 123.180 176.865 123.460 177.665 ;
        RECT 123.630 177.155 125.245 177.485 ;
        RECT 123.630 176.815 124.805 176.985 ;
        RECT 123.630 176.695 123.800 176.815 ;
        RECT 123.140 176.525 123.800 176.695 ;
        RECT 121.315 175.115 122.525 175.865 ;
        RECT 122.695 175.790 122.865 176.525 ;
        RECT 123.140 176.355 123.310 176.525 ;
        RECT 124.060 176.355 124.305 176.645 ;
        RECT 124.475 176.525 124.805 176.815 ;
        RECT 125.065 176.355 125.235 176.915 ;
        RECT 125.485 176.525 125.745 177.665 ;
        RECT 126.005 177.045 126.175 177.475 ;
        RECT 126.345 177.215 126.675 177.665 ;
        RECT 126.005 176.815 126.680 177.045 ;
        RECT 123.035 176.025 123.310 176.355 ;
        RECT 123.480 176.025 124.305 176.355 ;
        RECT 124.520 176.025 125.235 176.355 ;
        RECT 125.405 176.105 125.740 176.355 ;
        RECT 123.140 175.855 123.310 176.025 ;
        RECT 124.985 175.935 125.235 176.025 ;
        RECT 122.695 175.445 122.970 175.790 ;
        RECT 123.140 175.685 124.805 175.855 ;
        RECT 123.160 175.115 123.535 175.515 ;
        RECT 123.705 175.335 123.875 175.685 ;
        RECT 124.045 175.115 124.375 175.515 ;
        RECT 124.545 175.285 124.805 175.685 ;
        RECT 124.985 175.515 125.315 175.935 ;
        RECT 125.485 175.115 125.745 175.935 ;
        RECT 125.975 175.795 126.275 176.645 ;
        RECT 126.445 176.165 126.680 176.815 ;
        RECT 126.850 176.505 127.135 177.450 ;
        RECT 127.315 177.195 128.000 177.665 ;
        RECT 127.310 176.675 128.005 176.985 ;
        RECT 128.180 176.610 128.485 177.395 ;
        RECT 126.850 176.355 127.710 176.505 ;
        RECT 126.850 176.335 128.135 176.355 ;
        RECT 126.445 175.835 126.980 176.165 ;
        RECT 127.150 175.975 128.135 176.335 ;
        RECT 126.445 175.685 126.665 175.835 ;
        RECT 125.920 175.115 126.255 175.620 ;
        RECT 126.425 175.310 126.665 175.685 ;
        RECT 127.150 175.640 127.320 175.975 ;
        RECT 128.310 175.805 128.485 176.610 ;
        RECT 128.685 177.055 129.015 177.485 ;
        RECT 129.195 177.225 129.390 177.665 ;
        RECT 129.560 177.055 129.890 177.485 ;
        RECT 128.685 176.885 129.890 177.055 ;
        RECT 128.685 176.555 129.580 176.885 ;
        RECT 130.060 176.715 130.335 177.485 ;
        RECT 129.750 176.525 130.335 176.715 ;
        RECT 130.525 176.525 130.855 177.665 ;
        RECT 131.385 176.695 131.715 177.480 ;
        RECT 131.035 176.525 131.715 176.695 ;
        RECT 131.895 176.575 133.105 177.665 ;
        RECT 128.690 176.025 128.985 176.355 ;
        RECT 129.165 176.025 129.580 176.355 ;
        RECT 126.945 175.445 127.320 175.640 ;
        RECT 126.945 175.300 127.115 175.445 ;
        RECT 127.680 175.115 128.075 175.610 ;
        RECT 128.245 175.285 128.485 175.805 ;
        RECT 128.685 175.115 128.985 175.845 ;
        RECT 129.165 175.405 129.395 176.025 ;
        RECT 129.750 175.855 129.925 176.525 ;
        RECT 129.595 175.675 129.925 175.855 ;
        RECT 130.095 175.705 130.335 176.355 ;
        RECT 130.515 176.105 130.865 176.355 ;
        RECT 131.035 175.925 131.205 176.525 ;
        RECT 131.375 176.105 131.725 176.355 ;
        RECT 129.595 175.295 129.820 175.675 ;
        RECT 129.990 175.115 130.320 175.505 ;
        RECT 130.525 175.115 130.795 175.925 ;
        RECT 130.965 175.285 131.295 175.925 ;
        RECT 131.465 175.115 131.705 175.925 ;
        RECT 131.895 175.865 132.415 176.405 ;
        RECT 132.585 176.035 133.105 176.575 ;
        RECT 133.275 176.500 133.565 177.665 ;
        RECT 133.735 177.155 134.925 177.445 ;
        RECT 133.755 176.815 134.925 176.985 ;
        RECT 135.095 176.865 135.375 177.665 ;
        RECT 133.755 176.525 134.080 176.815 ;
        RECT 134.755 176.695 134.925 176.815 ;
        RECT 134.250 176.355 134.445 176.645 ;
        RECT 134.755 176.525 135.415 176.695 ;
        RECT 135.585 176.525 135.860 177.495 ;
        RECT 136.035 176.525 136.295 177.665 ;
        RECT 135.245 176.355 135.415 176.525 ;
        RECT 133.735 176.025 134.080 176.355 ;
        RECT 134.250 176.025 135.075 176.355 ;
        RECT 135.245 176.025 135.520 176.355 ;
        RECT 131.895 175.115 133.105 175.865 ;
        RECT 135.245 175.855 135.415 176.025 ;
        RECT 133.275 175.115 133.565 175.840 ;
        RECT 133.750 175.685 135.415 175.855 ;
        RECT 135.690 175.790 135.860 176.525 ;
        RECT 136.465 176.515 136.795 177.495 ;
        RECT 136.965 176.525 137.245 177.665 ;
        RECT 137.415 177.230 142.760 177.665 ;
        RECT 136.055 176.105 136.390 176.355 ;
        RECT 136.560 175.915 136.730 176.515 ;
        RECT 136.900 176.085 137.235 176.355 ;
        RECT 133.750 175.335 134.005 175.685 ;
        RECT 134.175 175.115 134.505 175.515 ;
        RECT 134.675 175.335 134.845 175.685 ;
        RECT 135.015 175.115 135.395 175.515 ;
        RECT 135.585 175.445 135.860 175.790 ;
        RECT 136.035 175.285 136.730 175.915 ;
        RECT 136.935 175.115 137.245 175.915 ;
        RECT 139.000 175.660 139.340 176.490 ;
        RECT 140.820 175.980 141.170 177.230 ;
        RECT 143.860 176.515 144.120 177.665 ;
        RECT 144.295 176.590 144.550 177.495 ;
        RECT 144.720 176.905 145.050 177.665 ;
        RECT 145.265 176.735 145.435 177.495 ;
        RECT 137.415 175.115 142.760 175.660 ;
        RECT 143.860 175.115 144.120 175.955 ;
        RECT 144.295 175.860 144.465 176.590 ;
        RECT 144.720 176.565 145.435 176.735 ;
        RECT 145.695 176.575 146.905 177.665 ;
        RECT 144.720 176.355 144.890 176.565 ;
        RECT 144.635 176.025 144.890 176.355 ;
        RECT 144.295 175.285 144.550 175.860 ;
        RECT 144.720 175.835 144.890 176.025 ;
        RECT 145.170 176.015 145.525 176.385 ;
        RECT 145.695 176.035 146.215 176.575 ;
        RECT 146.385 175.865 146.905 176.405 ;
        RECT 144.720 175.665 145.435 175.835 ;
        RECT 144.720 175.115 145.050 175.495 ;
        RECT 145.265 175.285 145.435 175.665 ;
        RECT 145.695 175.115 146.905 175.865 ;
        RECT 17.270 174.945 146.990 175.115 ;
        RECT 17.355 174.195 18.565 174.945 ;
        RECT 17.355 173.655 17.875 174.195 ;
        RECT 18.735 174.175 20.405 174.945 ;
        RECT 20.610 174.205 21.225 174.775 ;
        RECT 21.395 174.435 21.610 174.945 ;
        RECT 21.840 174.435 22.120 174.765 ;
        RECT 22.300 174.435 22.540 174.945 ;
        RECT 18.045 173.485 18.565 174.025 ;
        RECT 18.735 173.655 19.485 174.175 ;
        RECT 19.655 173.485 20.405 174.005 ;
        RECT 17.355 172.395 18.565 173.485 ;
        RECT 18.735 172.395 20.405 173.485 ;
        RECT 20.610 173.185 20.925 174.205 ;
        RECT 21.095 173.535 21.265 174.035 ;
        RECT 21.515 173.705 21.780 174.265 ;
        RECT 21.950 173.535 22.120 174.435 ;
        RECT 22.875 174.295 23.135 174.775 ;
        RECT 23.305 174.405 23.555 174.945 ;
        RECT 22.290 173.705 22.645 174.265 ;
        RECT 21.095 173.365 22.520 173.535 ;
        RECT 20.610 172.565 21.145 173.185 ;
        RECT 21.315 172.395 21.645 173.195 ;
        RECT 22.130 173.190 22.520 173.365 ;
        RECT 22.875 173.265 23.045 174.295 ;
        RECT 23.725 174.240 23.945 174.725 ;
        RECT 23.215 173.645 23.445 174.040 ;
        RECT 23.615 173.815 23.945 174.240 ;
        RECT 24.115 174.565 25.005 174.735 ;
        RECT 24.115 173.840 24.285 174.565 ;
        RECT 24.455 174.010 25.005 174.395 ;
        RECT 25.210 174.205 25.825 174.775 ;
        RECT 25.995 174.435 26.210 174.945 ;
        RECT 26.440 174.435 26.720 174.765 ;
        RECT 26.900 174.435 27.140 174.945 ;
        RECT 28.265 174.545 28.595 174.945 ;
        RECT 24.115 173.770 25.005 173.840 ;
        RECT 24.110 173.745 25.005 173.770 ;
        RECT 24.100 173.730 25.005 173.745 ;
        RECT 24.095 173.715 25.005 173.730 ;
        RECT 24.085 173.710 25.005 173.715 ;
        RECT 24.080 173.700 25.005 173.710 ;
        RECT 24.075 173.690 25.005 173.700 ;
        RECT 24.065 173.685 25.005 173.690 ;
        RECT 24.055 173.675 25.005 173.685 ;
        RECT 24.045 173.670 25.005 173.675 ;
        RECT 24.045 173.665 24.380 173.670 ;
        RECT 24.030 173.660 24.380 173.665 ;
        RECT 24.015 173.650 24.380 173.660 ;
        RECT 23.990 173.645 24.380 173.650 ;
        RECT 23.215 173.640 24.380 173.645 ;
        RECT 23.215 173.605 24.350 173.640 ;
        RECT 23.215 173.580 24.315 173.605 ;
        RECT 23.215 173.550 24.285 173.580 ;
        RECT 23.215 173.520 24.265 173.550 ;
        RECT 23.215 173.490 24.245 173.520 ;
        RECT 23.215 173.480 24.175 173.490 ;
        RECT 23.215 173.470 24.150 173.480 ;
        RECT 23.215 173.455 24.130 173.470 ;
        RECT 23.215 173.440 24.110 173.455 ;
        RECT 23.320 173.430 24.105 173.440 ;
        RECT 23.320 173.395 24.090 173.430 ;
        RECT 22.875 172.565 23.150 173.265 ;
        RECT 23.320 173.145 24.075 173.395 ;
        RECT 24.245 173.075 24.575 173.320 ;
        RECT 24.745 173.220 25.005 173.670 ;
        RECT 24.390 173.050 24.575 173.075 ;
        RECT 25.210 173.185 25.525 174.205 ;
        RECT 25.695 173.535 25.865 174.035 ;
        RECT 26.115 173.705 26.380 174.265 ;
        RECT 26.550 173.535 26.720 174.435 ;
        RECT 28.765 174.375 29.095 174.715 ;
        RECT 30.145 174.545 30.475 174.945 ;
        RECT 26.890 173.705 27.245 174.265 ;
        RECT 28.110 174.205 30.475 174.375 ;
        RECT 30.645 174.220 30.975 174.730 ;
        RECT 25.695 173.365 27.120 173.535 ;
        RECT 24.390 172.950 25.005 173.050 ;
        RECT 23.320 172.395 23.575 172.940 ;
        RECT 23.745 172.565 24.225 172.905 ;
        RECT 24.400 172.395 25.005 172.950 ;
        RECT 25.210 172.565 25.745 173.185 ;
        RECT 25.915 172.395 26.245 173.195 ;
        RECT 26.730 173.190 27.120 173.365 ;
        RECT 28.110 173.205 28.280 174.205 ;
        RECT 30.305 174.035 30.475 174.205 ;
        RECT 28.450 173.375 28.695 174.035 ;
        RECT 28.910 173.375 29.175 174.035 ;
        RECT 29.370 173.375 29.655 174.035 ;
        RECT 29.830 173.705 30.135 174.035 ;
        RECT 30.305 173.705 30.615 174.035 ;
        RECT 29.830 173.375 30.045 173.705 ;
        RECT 28.110 173.035 28.565 173.205 ;
        RECT 28.235 172.605 28.565 173.035 ;
        RECT 28.745 173.035 30.035 173.205 ;
        RECT 28.745 172.615 28.995 173.035 ;
        RECT 29.225 172.395 29.555 172.865 ;
        RECT 29.785 172.615 30.035 173.035 ;
        RECT 30.225 172.395 30.475 173.535 ;
        RECT 30.785 173.455 30.975 174.220 ;
        RECT 31.215 174.125 31.425 174.945 ;
        RECT 31.595 174.145 31.925 174.775 ;
        RECT 31.595 173.545 31.845 174.145 ;
        RECT 32.095 174.125 32.325 174.945 ;
        RECT 32.535 174.175 36.045 174.945 ;
        RECT 36.710 174.205 37.325 174.775 ;
        RECT 37.495 174.435 37.710 174.945 ;
        RECT 37.940 174.435 38.220 174.765 ;
        RECT 38.400 174.435 38.640 174.945 ;
        RECT 32.015 173.705 32.345 173.955 ;
        RECT 32.535 173.655 34.185 174.175 ;
        RECT 30.645 172.605 30.975 173.455 ;
        RECT 31.215 172.395 31.425 173.535 ;
        RECT 31.595 172.565 31.925 173.545 ;
        RECT 32.095 172.395 32.325 173.535 ;
        RECT 34.355 173.485 36.045 174.005 ;
        RECT 32.535 172.395 36.045 173.485 ;
        RECT 36.710 173.185 37.025 174.205 ;
        RECT 37.195 173.535 37.365 174.035 ;
        RECT 37.615 173.705 37.880 174.265 ;
        RECT 38.050 173.535 38.220 174.435 ;
        RECT 38.390 173.705 38.745 174.265 ;
        RECT 39.035 174.125 39.245 174.945 ;
        RECT 39.415 174.145 39.745 174.775 ;
        RECT 39.415 173.545 39.665 174.145 ;
        RECT 39.915 174.125 40.145 174.945 ;
        RECT 40.355 174.195 41.565 174.945 ;
        RECT 39.835 173.705 40.165 173.955 ;
        RECT 40.355 173.655 40.875 174.195 ;
        RECT 41.745 174.135 42.015 174.945 ;
        RECT 42.185 174.135 42.515 174.775 ;
        RECT 42.685 174.135 42.925 174.945 ;
        RECT 43.115 174.220 43.405 174.945 ;
        RECT 43.575 174.445 43.835 174.775 ;
        RECT 44.005 174.585 44.335 174.945 ;
        RECT 44.590 174.565 45.890 174.775 ;
        RECT 43.575 174.435 43.805 174.445 ;
        RECT 37.195 173.365 38.620 173.535 ;
        RECT 36.710 172.565 37.245 173.185 ;
        RECT 37.415 172.395 37.745 173.195 ;
        RECT 38.230 173.190 38.620 173.365 ;
        RECT 39.035 172.395 39.245 173.535 ;
        RECT 39.415 172.565 39.745 173.545 ;
        RECT 39.915 172.395 40.145 173.535 ;
        RECT 41.045 173.485 41.565 174.025 ;
        RECT 41.735 173.705 42.085 173.955 ;
        RECT 42.255 173.535 42.425 174.135 ;
        RECT 42.595 173.705 42.945 173.955 ;
        RECT 40.355 172.395 41.565 173.485 ;
        RECT 41.745 172.395 42.075 173.535 ;
        RECT 42.255 173.365 42.935 173.535 ;
        RECT 42.605 172.580 42.935 173.365 ;
        RECT 43.115 172.395 43.405 173.560 ;
        RECT 43.575 173.245 43.745 174.435 ;
        RECT 44.590 174.415 44.760 174.565 ;
        RECT 44.005 174.290 44.760 174.415 ;
        RECT 43.915 174.245 44.760 174.290 ;
        RECT 43.915 174.125 44.185 174.245 ;
        RECT 43.915 173.550 44.085 174.125 ;
        RECT 44.315 173.685 44.725 173.990 ;
        RECT 45.015 173.955 45.225 174.355 ;
        RECT 44.895 173.745 45.225 173.955 ;
        RECT 45.470 173.955 45.690 174.355 ;
        RECT 46.165 174.180 46.620 174.945 ;
        RECT 46.795 174.145 47.490 174.775 ;
        RECT 47.695 174.145 48.005 174.945 ;
        RECT 48.685 174.290 49.015 174.725 ;
        RECT 49.185 174.335 49.355 174.945 ;
        RECT 48.635 174.205 49.015 174.290 ;
        RECT 49.525 174.205 49.855 174.730 ;
        RECT 50.115 174.415 50.325 174.945 ;
        RECT 50.600 174.495 51.385 174.665 ;
        RECT 51.555 174.495 51.960 174.665 ;
        RECT 48.635 174.165 48.860 174.205 ;
        RECT 45.470 173.745 45.945 173.955 ;
        RECT 46.135 173.755 46.625 173.955 ;
        RECT 46.815 173.705 47.150 173.955 ;
        RECT 43.915 173.515 44.115 173.550 ;
        RECT 45.445 173.515 46.620 173.575 ;
        RECT 47.320 173.545 47.490 174.145 ;
        RECT 47.660 173.705 47.995 173.975 ;
        RECT 48.635 173.585 48.805 174.165 ;
        RECT 49.525 174.035 49.725 174.205 ;
        RECT 50.600 174.035 50.770 174.495 ;
        RECT 48.975 173.705 49.725 174.035 ;
        RECT 49.895 173.705 50.770 174.035 ;
        RECT 43.915 173.405 46.620 173.515 ;
        RECT 43.975 173.345 45.775 173.405 ;
        RECT 45.445 173.315 45.775 173.345 ;
        RECT 43.575 172.565 43.835 173.245 ;
        RECT 44.005 172.395 44.255 173.175 ;
        RECT 44.505 173.145 45.340 173.155 ;
        RECT 45.930 173.145 46.115 173.235 ;
        RECT 44.505 172.945 46.115 173.145 ;
        RECT 44.505 172.565 44.755 172.945 ;
        RECT 45.885 172.905 46.115 172.945 ;
        RECT 46.365 172.785 46.620 173.405 ;
        RECT 44.925 172.395 45.280 172.775 ;
        RECT 46.285 172.565 46.620 172.785 ;
        RECT 46.795 172.395 47.055 173.535 ;
        RECT 47.225 172.565 47.555 173.545 ;
        RECT 48.635 173.535 48.850 173.585 ;
        RECT 47.725 172.395 48.005 173.535 ;
        RECT 48.635 173.455 49.025 173.535 ;
        RECT 48.695 172.610 49.025 173.455 ;
        RECT 49.535 173.500 49.725 173.705 ;
        RECT 49.195 172.395 49.365 173.405 ;
        RECT 49.535 173.125 50.430 173.500 ;
        RECT 49.535 172.565 49.875 173.125 ;
        RECT 50.105 172.395 50.420 172.895 ;
        RECT 50.600 172.865 50.770 173.705 ;
        RECT 50.940 173.995 51.405 174.325 ;
        RECT 51.790 174.265 51.960 174.495 ;
        RECT 52.140 174.445 52.510 174.945 ;
        RECT 52.830 174.495 53.505 174.665 ;
        RECT 53.700 174.495 54.035 174.665 ;
        RECT 50.940 173.035 51.260 173.995 ;
        RECT 51.790 173.965 52.620 174.265 ;
        RECT 51.430 173.065 51.620 173.785 ;
        RECT 51.790 172.895 51.960 173.965 ;
        RECT 52.420 173.935 52.620 173.965 ;
        RECT 52.130 173.715 52.300 173.785 ;
        RECT 52.830 173.715 53.000 174.495 ;
        RECT 53.865 174.355 54.035 174.495 ;
        RECT 54.205 174.485 54.455 174.945 ;
        RECT 52.130 173.545 53.000 173.715 ;
        RECT 53.170 174.075 53.695 174.295 ;
        RECT 53.865 174.225 54.090 174.355 ;
        RECT 52.130 173.455 52.640 173.545 ;
        RECT 50.600 172.695 51.485 172.865 ;
        RECT 51.710 172.565 51.960 172.895 ;
        RECT 52.130 172.395 52.300 173.195 ;
        RECT 52.470 172.840 52.640 173.455 ;
        RECT 53.170 173.375 53.340 174.075 ;
        RECT 52.810 173.010 53.340 173.375 ;
        RECT 53.510 173.310 53.750 173.905 ;
        RECT 53.920 173.120 54.090 174.225 ;
        RECT 54.260 173.365 54.540 174.315 ;
        RECT 53.785 172.990 54.090 173.120 ;
        RECT 52.470 172.670 53.575 172.840 ;
        RECT 53.785 172.565 54.035 172.990 ;
        RECT 54.205 172.395 54.470 172.855 ;
        RECT 54.710 172.565 54.895 174.685 ;
        RECT 55.065 174.565 55.395 174.945 ;
        RECT 55.565 174.395 55.735 174.685 ;
        RECT 55.995 174.400 61.340 174.945 ;
        RECT 55.070 174.225 55.735 174.395 ;
        RECT 55.070 173.235 55.300 174.225 ;
        RECT 55.470 173.405 55.820 174.055 ;
        RECT 57.580 173.570 57.920 174.400 ;
        RECT 61.605 174.395 61.775 174.685 ;
        RECT 61.945 174.565 62.275 174.945 ;
        RECT 61.605 174.225 62.270 174.395 ;
        RECT 55.070 173.065 55.735 173.235 ;
        RECT 55.065 172.395 55.395 172.895 ;
        RECT 55.565 172.565 55.735 173.065 ;
        RECT 59.400 172.830 59.750 174.080 ;
        RECT 61.520 173.405 61.870 174.055 ;
        RECT 62.040 173.235 62.270 174.225 ;
        RECT 61.605 173.065 62.270 173.235 ;
        RECT 55.995 172.395 61.340 172.830 ;
        RECT 61.605 172.565 61.775 173.065 ;
        RECT 61.945 172.395 62.275 172.895 ;
        RECT 62.445 172.565 62.630 174.685 ;
        RECT 62.885 174.485 63.135 174.945 ;
        RECT 63.305 174.495 63.640 174.665 ;
        RECT 63.835 174.495 64.510 174.665 ;
        RECT 63.305 174.355 63.475 174.495 ;
        RECT 62.800 173.365 63.080 174.315 ;
        RECT 63.250 174.225 63.475 174.355 ;
        RECT 63.250 173.120 63.420 174.225 ;
        RECT 63.645 174.075 64.170 174.295 ;
        RECT 63.590 173.310 63.830 173.905 ;
        RECT 64.000 173.375 64.170 174.075 ;
        RECT 64.340 173.715 64.510 174.495 ;
        RECT 64.830 174.445 65.200 174.945 ;
        RECT 65.380 174.495 65.785 174.665 ;
        RECT 65.955 174.495 66.740 174.665 ;
        RECT 65.380 174.265 65.550 174.495 ;
        RECT 64.720 173.965 65.550 174.265 ;
        RECT 65.935 173.995 66.400 174.325 ;
        RECT 64.720 173.935 64.920 173.965 ;
        RECT 65.040 173.715 65.210 173.785 ;
        RECT 64.340 173.545 65.210 173.715 ;
        RECT 64.700 173.455 65.210 173.545 ;
        RECT 63.250 172.990 63.555 173.120 ;
        RECT 64.000 173.010 64.530 173.375 ;
        RECT 62.870 172.395 63.135 172.855 ;
        RECT 63.305 172.565 63.555 172.990 ;
        RECT 64.700 172.840 64.870 173.455 ;
        RECT 63.765 172.670 64.870 172.840 ;
        RECT 65.040 172.395 65.210 173.195 ;
        RECT 65.380 172.895 65.550 173.965 ;
        RECT 65.720 173.065 65.910 173.785 ;
        RECT 66.080 173.035 66.400 173.995 ;
        RECT 66.570 174.035 66.740 174.495 ;
        RECT 67.015 174.415 67.225 174.945 ;
        RECT 67.485 174.205 67.815 174.730 ;
        RECT 67.985 174.335 68.155 174.945 ;
        RECT 68.325 174.290 68.655 174.725 ;
        RECT 68.325 174.205 68.705 174.290 ;
        RECT 68.875 174.220 69.165 174.945 ;
        RECT 69.335 174.400 74.680 174.945 ;
        RECT 67.615 174.035 67.815 174.205 ;
        RECT 68.480 174.165 68.705 174.205 ;
        RECT 66.570 173.705 67.445 174.035 ;
        RECT 67.615 173.705 68.365 174.035 ;
        RECT 65.380 172.565 65.630 172.895 ;
        RECT 66.570 172.865 66.740 173.705 ;
        RECT 67.615 173.500 67.805 173.705 ;
        RECT 68.535 173.585 68.705 174.165 ;
        RECT 68.490 173.535 68.705 173.585 ;
        RECT 70.920 173.570 71.260 174.400 ;
        RECT 74.855 174.175 76.525 174.945 ;
        RECT 76.745 174.290 77.075 174.725 ;
        RECT 77.245 174.335 77.415 174.945 ;
        RECT 76.695 174.205 77.075 174.290 ;
        RECT 77.585 174.205 77.915 174.730 ;
        RECT 78.175 174.415 78.385 174.945 ;
        RECT 78.660 174.495 79.445 174.665 ;
        RECT 79.615 174.495 80.020 174.665 ;
        RECT 66.910 173.125 67.805 173.500 ;
        RECT 68.315 173.455 68.705 173.535 ;
        RECT 65.855 172.695 66.740 172.865 ;
        RECT 66.920 172.395 67.235 172.895 ;
        RECT 67.465 172.565 67.805 173.125 ;
        RECT 67.975 172.395 68.145 173.405 ;
        RECT 68.315 172.610 68.645 173.455 ;
        RECT 68.875 172.395 69.165 173.560 ;
        RECT 72.740 172.830 73.090 174.080 ;
        RECT 74.855 173.655 75.605 174.175 ;
        RECT 76.695 174.165 76.920 174.205 ;
        RECT 75.775 173.485 76.525 174.005 ;
        RECT 69.335 172.395 74.680 172.830 ;
        RECT 74.855 172.395 76.525 173.485 ;
        RECT 76.695 173.585 76.865 174.165 ;
        RECT 77.585 174.035 77.785 174.205 ;
        RECT 78.660 174.035 78.830 174.495 ;
        RECT 77.035 173.705 77.785 174.035 ;
        RECT 77.955 173.705 78.830 174.035 ;
        RECT 76.695 173.535 76.910 173.585 ;
        RECT 76.695 173.455 77.085 173.535 ;
        RECT 76.755 172.610 77.085 173.455 ;
        RECT 77.595 173.500 77.785 173.705 ;
        RECT 77.255 172.395 77.425 173.405 ;
        RECT 77.595 173.125 78.490 173.500 ;
        RECT 77.595 172.565 77.935 173.125 ;
        RECT 78.165 172.395 78.480 172.895 ;
        RECT 78.660 172.865 78.830 173.705 ;
        RECT 79.000 173.995 79.465 174.325 ;
        RECT 79.850 174.265 80.020 174.495 ;
        RECT 80.200 174.445 80.570 174.945 ;
        RECT 80.890 174.495 81.565 174.665 ;
        RECT 81.760 174.495 82.095 174.665 ;
        RECT 79.000 173.035 79.320 173.995 ;
        RECT 79.850 173.965 80.680 174.265 ;
        RECT 79.490 173.065 79.680 173.785 ;
        RECT 79.850 172.895 80.020 173.965 ;
        RECT 80.480 173.935 80.680 173.965 ;
        RECT 80.190 173.715 80.360 173.785 ;
        RECT 80.890 173.715 81.060 174.495 ;
        RECT 81.925 174.355 82.095 174.495 ;
        RECT 82.265 174.485 82.515 174.945 ;
        RECT 80.190 173.545 81.060 173.715 ;
        RECT 81.230 174.075 81.755 174.295 ;
        RECT 81.925 174.225 82.150 174.355 ;
        RECT 80.190 173.455 80.700 173.545 ;
        RECT 78.660 172.695 79.545 172.865 ;
        RECT 79.770 172.565 80.020 172.895 ;
        RECT 80.190 172.395 80.360 173.195 ;
        RECT 80.530 172.840 80.700 173.455 ;
        RECT 81.230 173.375 81.400 174.075 ;
        RECT 80.870 173.010 81.400 173.375 ;
        RECT 81.570 173.310 81.810 173.905 ;
        RECT 81.980 173.120 82.150 174.225 ;
        RECT 82.320 173.365 82.600 174.315 ;
        RECT 81.845 172.990 82.150 173.120 ;
        RECT 80.530 172.670 81.635 172.840 ;
        RECT 81.845 172.565 82.095 172.990 ;
        RECT 82.265 172.395 82.530 172.855 ;
        RECT 82.770 172.565 82.955 174.685 ;
        RECT 83.125 174.565 83.455 174.945 ;
        RECT 83.625 174.395 83.795 174.685 ;
        RECT 83.130 174.225 83.795 174.395 ;
        RECT 83.130 173.235 83.360 174.225 ;
        RECT 84.055 174.220 84.315 174.775 ;
        RECT 84.485 174.500 84.915 174.945 ;
        RECT 85.150 174.375 85.320 174.775 ;
        RECT 85.490 174.545 86.210 174.945 ;
        RECT 83.530 173.405 83.880 174.055 ;
        RECT 84.055 173.505 84.230 174.220 ;
        RECT 85.150 174.205 86.030 174.375 ;
        RECT 86.380 174.330 86.550 174.775 ;
        RECT 87.125 174.435 87.525 174.945 ;
        RECT 87.755 174.435 87.995 174.945 ;
        RECT 84.400 173.705 84.655 174.035 ;
        RECT 83.130 173.065 83.795 173.235 ;
        RECT 83.125 172.395 83.455 172.895 ;
        RECT 83.625 172.565 83.795 173.065 ;
        RECT 84.055 172.565 84.315 173.505 ;
        RECT 84.485 173.225 84.655 173.705 ;
        RECT 84.880 173.415 85.210 174.035 ;
        RECT 85.380 173.655 85.670 174.035 ;
        RECT 85.860 173.485 86.030 174.205 ;
        RECT 85.510 173.315 86.030 173.485 ;
        RECT 86.200 174.160 86.550 174.330 ;
        RECT 84.485 173.055 85.245 173.225 ;
        RECT 85.510 173.125 85.680 173.315 ;
        RECT 86.200 173.135 86.370 174.160 ;
        RECT 86.790 173.675 87.050 174.265 ;
        RECT 86.570 173.375 87.050 173.675 ;
        RECT 87.250 173.375 87.510 174.265 ;
        RECT 87.740 173.705 87.995 174.265 ;
        RECT 88.165 174.205 88.495 174.740 ;
        RECT 88.710 174.205 88.880 174.945 ;
        RECT 89.090 174.295 89.420 174.765 ;
        RECT 89.590 174.465 89.760 174.945 ;
        RECT 89.930 174.295 90.260 174.765 ;
        RECT 90.430 174.465 90.600 174.945 ;
        RECT 88.165 173.535 88.345 174.205 ;
        RECT 89.090 174.125 90.785 174.295 ;
        RECT 88.515 173.705 88.890 174.035 ;
        RECT 89.060 173.785 90.270 173.955 ;
        RECT 89.060 173.535 89.265 173.785 ;
        RECT 90.440 173.535 90.785 174.125 ;
        RECT 90.955 174.175 94.465 174.945 ;
        RECT 94.635 174.220 94.925 174.945 ;
        RECT 95.095 174.175 98.605 174.945 ;
        RECT 90.955 173.655 92.605 174.175 ;
        RECT 87.805 173.365 89.265 173.535 ;
        RECT 89.930 173.365 90.785 173.535 ;
        RECT 92.775 173.485 94.465 174.005 ;
        RECT 95.095 173.655 96.745 174.175 ;
        RECT 98.775 174.145 99.085 174.945 ;
        RECT 99.290 174.145 99.985 174.775 ;
        RECT 100.205 174.290 100.535 174.725 ;
        RECT 100.705 174.335 100.875 174.945 ;
        RECT 100.155 174.205 100.535 174.290 ;
        RECT 101.045 174.205 101.375 174.730 ;
        RECT 101.635 174.415 101.845 174.945 ;
        RECT 102.120 174.495 102.905 174.665 ;
        RECT 103.075 174.495 103.480 174.665 ;
        RECT 100.155 174.165 100.380 174.205 ;
        RECT 85.075 172.830 85.245 173.055 ;
        RECT 85.960 172.965 86.370 173.135 ;
        RECT 86.545 173.025 87.485 173.195 ;
        RECT 85.960 172.830 86.215 172.965 ;
        RECT 84.485 172.395 84.815 172.795 ;
        RECT 85.075 172.660 86.215 172.830 ;
        RECT 86.545 172.775 86.715 173.025 ;
        RECT 85.960 172.565 86.215 172.660 ;
        RECT 86.385 172.605 86.715 172.775 ;
        RECT 86.885 172.395 87.135 172.855 ;
        RECT 87.305 172.565 87.485 173.025 ;
        RECT 87.805 172.565 88.165 173.365 ;
        RECT 89.930 173.195 90.260 173.365 ;
        RECT 88.710 172.395 88.880 173.195 ;
        RECT 89.090 173.025 90.260 173.195 ;
        RECT 89.090 172.565 89.420 173.025 ;
        RECT 89.590 172.395 89.760 172.855 ;
        RECT 89.930 172.565 90.260 173.025 ;
        RECT 90.430 172.395 90.600 173.195 ;
        RECT 90.955 172.395 94.465 173.485 ;
        RECT 94.635 172.395 94.925 173.560 ;
        RECT 96.915 173.485 98.605 174.005 ;
        RECT 98.785 173.705 99.120 173.975 ;
        RECT 99.290 173.545 99.460 174.145 ;
        RECT 99.630 173.705 99.965 173.955 ;
        RECT 100.155 173.585 100.325 174.165 ;
        RECT 101.045 174.035 101.245 174.205 ;
        RECT 102.120 174.035 102.290 174.495 ;
        RECT 100.495 173.705 101.245 174.035 ;
        RECT 101.415 173.705 102.290 174.035 ;
        RECT 95.095 172.395 98.605 173.485 ;
        RECT 98.775 172.395 99.055 173.535 ;
        RECT 99.225 172.565 99.555 173.545 ;
        RECT 100.155 173.535 100.370 173.585 ;
        RECT 99.725 172.395 99.985 173.535 ;
        RECT 100.155 173.455 100.545 173.535 ;
        RECT 100.215 172.610 100.545 173.455 ;
        RECT 101.055 173.500 101.245 173.705 ;
        RECT 100.715 172.395 100.885 173.405 ;
        RECT 101.055 173.125 101.950 173.500 ;
        RECT 101.055 172.565 101.395 173.125 ;
        RECT 101.625 172.395 101.940 172.895 ;
        RECT 102.120 172.865 102.290 173.705 ;
        RECT 102.460 173.995 102.925 174.325 ;
        RECT 103.310 174.265 103.480 174.495 ;
        RECT 103.660 174.445 104.030 174.945 ;
        RECT 104.350 174.495 105.025 174.665 ;
        RECT 105.220 174.495 105.555 174.665 ;
        RECT 102.460 173.035 102.780 173.995 ;
        RECT 103.310 173.965 104.140 174.265 ;
        RECT 102.950 173.065 103.140 173.785 ;
        RECT 103.310 172.895 103.480 173.965 ;
        RECT 103.940 173.935 104.140 173.965 ;
        RECT 103.650 173.715 103.820 173.785 ;
        RECT 104.350 173.715 104.520 174.495 ;
        RECT 105.385 174.355 105.555 174.495 ;
        RECT 105.725 174.485 105.975 174.945 ;
        RECT 103.650 173.545 104.520 173.715 ;
        RECT 104.690 174.075 105.215 174.295 ;
        RECT 105.385 174.225 105.610 174.355 ;
        RECT 103.650 173.455 104.160 173.545 ;
        RECT 102.120 172.695 103.005 172.865 ;
        RECT 103.230 172.565 103.480 172.895 ;
        RECT 103.650 172.395 103.820 173.195 ;
        RECT 103.990 172.840 104.160 173.455 ;
        RECT 104.690 173.375 104.860 174.075 ;
        RECT 104.330 173.010 104.860 173.375 ;
        RECT 105.030 173.310 105.270 173.905 ;
        RECT 105.440 173.120 105.610 174.225 ;
        RECT 105.780 173.365 106.060 174.315 ;
        RECT 105.305 172.990 105.610 173.120 ;
        RECT 103.990 172.670 105.095 172.840 ;
        RECT 105.305 172.565 105.555 172.990 ;
        RECT 105.725 172.395 105.990 172.855 ;
        RECT 106.230 172.565 106.415 174.685 ;
        RECT 106.585 174.565 106.915 174.945 ;
        RECT 107.085 174.395 107.255 174.685 ;
        RECT 106.590 174.225 107.255 174.395 ;
        RECT 106.590 173.235 106.820 174.225 ;
        RECT 107.515 174.205 107.900 174.775 ;
        RECT 108.070 174.485 108.395 174.945 ;
        RECT 108.915 174.315 109.195 174.775 ;
        RECT 106.990 173.405 107.340 174.055 ;
        RECT 107.515 173.535 107.795 174.205 ;
        RECT 108.070 174.145 109.195 174.315 ;
        RECT 108.070 174.035 108.520 174.145 ;
        RECT 107.965 173.705 108.520 174.035 ;
        RECT 109.385 173.975 109.785 174.775 ;
        RECT 110.185 174.485 110.455 174.945 ;
        RECT 110.625 174.315 110.910 174.775 ;
        RECT 106.590 173.065 107.255 173.235 ;
        RECT 106.585 172.395 106.915 172.895 ;
        RECT 107.085 172.565 107.255 173.065 ;
        RECT 107.515 172.565 107.900 173.535 ;
        RECT 108.070 173.245 108.520 173.705 ;
        RECT 108.690 173.415 109.785 173.975 ;
        RECT 108.070 173.025 109.195 173.245 ;
        RECT 108.070 172.395 108.395 172.855 ;
        RECT 108.915 172.565 109.195 173.025 ;
        RECT 109.385 172.565 109.785 173.415 ;
        RECT 109.955 174.145 110.910 174.315 ;
        RECT 109.955 173.245 110.165 174.145 ;
        RECT 110.335 173.415 111.025 173.975 ;
        RECT 111.215 173.365 111.445 174.705 ;
        RECT 111.625 173.865 111.855 174.765 ;
        RECT 112.055 174.165 112.300 174.945 ;
        RECT 112.470 174.405 112.900 174.765 ;
        RECT 113.480 174.575 114.210 174.945 ;
        RECT 112.470 174.215 114.210 174.405 ;
        RECT 112.470 173.985 112.690 174.215 ;
        RECT 109.955 173.025 110.910 173.245 ;
        RECT 111.625 173.185 111.965 173.865 ;
        RECT 110.185 172.395 110.455 172.855 ;
        RECT 110.625 172.565 110.910 173.025 ;
        RECT 111.215 172.985 111.965 173.185 ;
        RECT 112.145 173.685 112.690 173.985 ;
        RECT 111.215 172.595 111.455 172.985 ;
        RECT 111.625 172.395 111.975 172.805 ;
        RECT 112.145 172.575 112.475 173.685 ;
        RECT 112.860 173.415 113.285 174.035 ;
        RECT 113.480 173.415 113.740 174.035 ;
        RECT 113.950 173.705 114.210 174.215 ;
        RECT 112.645 173.045 113.670 173.245 ;
        RECT 112.645 172.575 112.825 173.045 ;
        RECT 112.995 172.395 113.325 172.875 ;
        RECT 113.500 172.575 113.670 173.045 ;
        RECT 113.935 172.395 114.220 173.535 ;
        RECT 114.410 172.575 114.690 174.765 ;
        RECT 114.875 174.445 115.215 174.945 ;
        RECT 114.875 173.705 115.215 174.275 ;
        RECT 115.385 174.035 115.630 174.725 ;
        RECT 115.825 174.445 116.155 174.945 ;
        RECT 116.355 174.375 116.525 174.725 ;
        RECT 116.700 174.545 117.030 174.945 ;
        RECT 117.200 174.375 117.370 174.725 ;
        RECT 117.540 174.545 117.920 174.945 ;
        RECT 116.355 174.205 117.940 174.375 ;
        RECT 118.110 174.270 118.385 174.615 ;
        RECT 117.770 174.035 117.940 174.205 ;
        RECT 115.385 173.705 116.040 174.035 ;
        RECT 114.875 172.395 115.215 173.470 ;
        RECT 115.385 173.110 115.625 173.705 ;
        RECT 115.820 173.245 116.140 173.535 ;
        RECT 116.310 173.415 117.050 174.035 ;
        RECT 117.220 173.705 117.600 174.035 ;
        RECT 117.770 173.705 118.045 174.035 ;
        RECT 117.770 173.535 117.940 173.705 ;
        RECT 118.215 173.535 118.385 174.270 ;
        RECT 118.555 174.175 120.225 174.945 ;
        RECT 120.395 174.220 120.685 174.945 ;
        RECT 120.855 174.295 121.115 174.775 ;
        RECT 121.285 174.405 121.535 174.945 ;
        RECT 118.555 173.655 119.305 174.175 ;
        RECT 117.280 173.365 117.940 173.535 ;
        RECT 117.280 173.245 117.450 173.365 ;
        RECT 115.820 173.075 117.450 173.245 ;
        RECT 115.395 172.735 117.450 172.905 ;
        RECT 115.400 172.615 117.450 172.735 ;
        RECT 117.620 172.395 117.900 173.195 ;
        RECT 118.110 172.565 118.385 173.535 ;
        RECT 119.475 173.485 120.225 174.005 ;
        RECT 118.555 172.395 120.225 173.485 ;
        RECT 120.395 172.395 120.685 173.560 ;
        RECT 120.855 173.265 121.025 174.295 ;
        RECT 121.705 174.240 121.925 174.725 ;
        RECT 121.195 173.645 121.425 174.040 ;
        RECT 121.595 173.815 121.925 174.240 ;
        RECT 122.095 174.565 122.985 174.735 ;
        RECT 122.095 173.840 122.265 174.565 ;
        RECT 123.215 174.485 123.460 174.945 ;
        RECT 122.435 174.010 122.985 174.395 ;
        RECT 122.095 173.770 122.985 173.840 ;
        RECT 122.090 173.745 122.985 173.770 ;
        RECT 122.080 173.730 122.985 173.745 ;
        RECT 122.075 173.715 122.985 173.730 ;
        RECT 122.065 173.710 122.985 173.715 ;
        RECT 122.060 173.700 122.985 173.710 ;
        RECT 123.155 173.705 123.470 174.315 ;
        RECT 123.640 173.955 123.890 174.765 ;
        RECT 124.060 174.420 124.320 174.945 ;
        RECT 124.490 174.295 124.750 174.750 ;
        RECT 124.920 174.465 125.180 174.945 ;
        RECT 125.350 174.295 125.610 174.750 ;
        RECT 125.780 174.465 126.040 174.945 ;
        RECT 126.210 174.295 126.470 174.750 ;
        RECT 126.640 174.465 126.900 174.945 ;
        RECT 127.070 174.295 127.330 174.750 ;
        RECT 127.500 174.465 127.800 174.945 ;
        RECT 129.295 174.385 129.625 174.775 ;
        RECT 129.795 174.555 130.980 174.725 ;
        RECT 131.240 174.475 131.410 174.945 ;
        RECT 124.490 174.125 127.800 174.295 ;
        RECT 129.295 174.205 129.805 174.385 ;
        RECT 123.640 173.705 126.660 173.955 ;
        RECT 122.055 173.690 122.985 173.700 ;
        RECT 122.045 173.685 122.985 173.690 ;
        RECT 122.035 173.675 122.985 173.685 ;
        RECT 122.025 173.670 122.985 173.675 ;
        RECT 122.025 173.665 122.360 173.670 ;
        RECT 122.010 173.660 122.360 173.665 ;
        RECT 121.995 173.650 122.360 173.660 ;
        RECT 121.970 173.645 122.360 173.650 ;
        RECT 121.195 173.640 122.360 173.645 ;
        RECT 121.195 173.605 122.330 173.640 ;
        RECT 121.195 173.580 122.295 173.605 ;
        RECT 121.195 173.550 122.265 173.580 ;
        RECT 121.195 173.520 122.245 173.550 ;
        RECT 121.195 173.490 122.225 173.520 ;
        RECT 121.195 173.480 122.155 173.490 ;
        RECT 121.195 173.470 122.130 173.480 ;
        RECT 121.195 173.455 122.110 173.470 ;
        RECT 121.195 173.440 122.090 173.455 ;
        RECT 121.300 173.430 122.085 173.440 ;
        RECT 121.300 173.395 122.070 173.430 ;
        RECT 120.855 172.565 121.130 173.265 ;
        RECT 121.300 173.145 122.055 173.395 ;
        RECT 122.225 173.075 122.555 173.320 ;
        RECT 122.725 173.220 122.985 173.670 ;
        RECT 122.370 173.050 122.555 173.075 ;
        RECT 122.370 172.950 122.985 173.050 ;
        RECT 121.300 172.395 121.555 172.940 ;
        RECT 121.725 172.565 122.205 172.905 ;
        RECT 122.380 172.395 122.985 172.950 ;
        RECT 123.165 172.395 123.460 173.505 ;
        RECT 123.640 172.570 123.890 173.705 ;
        RECT 126.830 173.535 127.800 174.125 ;
        RECT 129.135 173.745 129.465 174.035 ;
        RECT 129.635 173.575 129.805 174.205 ;
        RECT 130.210 174.295 130.595 174.385 ;
        RECT 131.580 174.295 131.910 174.760 ;
        RECT 130.210 174.125 131.910 174.295 ;
        RECT 132.080 174.125 132.250 174.945 ;
        RECT 132.420 174.125 133.105 174.765 ;
        RECT 129.975 173.745 130.305 173.955 ;
        RECT 130.485 173.705 130.865 173.955 ;
        RECT 131.055 173.925 131.540 173.955 ;
        RECT 131.035 173.755 131.540 173.925 ;
        RECT 124.060 172.395 124.320 173.505 ;
        RECT 124.490 173.295 127.800 173.535 ;
        RECT 129.290 173.405 130.375 173.575 ;
        RECT 124.490 172.570 124.750 173.295 ;
        RECT 124.920 172.395 125.180 173.125 ;
        RECT 125.350 172.570 125.610 173.295 ;
        RECT 125.780 172.395 126.040 173.125 ;
        RECT 126.210 172.570 126.470 173.295 ;
        RECT 126.640 172.395 126.900 173.125 ;
        RECT 127.070 172.570 127.330 173.295 ;
        RECT 127.500 172.395 127.795 173.125 ;
        RECT 129.290 172.565 129.590 173.405 ;
        RECT 129.785 172.395 130.035 173.235 ;
        RECT 130.205 173.155 130.375 173.405 ;
        RECT 130.545 173.325 130.865 173.705 ;
        RECT 131.055 173.745 131.540 173.755 ;
        RECT 131.730 173.745 132.180 173.955 ;
        RECT 132.350 173.745 132.685 173.955 ;
        RECT 131.055 173.325 131.430 173.745 ;
        RECT 132.350 173.575 132.520 173.745 ;
        RECT 131.600 173.405 132.520 173.575 ;
        RECT 131.600 173.155 131.770 173.405 ;
        RECT 130.205 172.985 131.770 173.155 ;
        RECT 130.625 172.565 131.430 172.985 ;
        RECT 131.940 172.395 132.270 173.235 ;
        RECT 132.855 173.155 133.105 174.125 ;
        RECT 132.440 172.565 133.105 173.155 ;
        RECT 133.770 174.205 134.385 174.775 ;
        RECT 134.555 174.435 134.770 174.945 ;
        RECT 135.000 174.435 135.280 174.765 ;
        RECT 135.460 174.435 135.700 174.945 ;
        RECT 133.770 173.185 134.085 174.205 ;
        RECT 134.255 173.535 134.425 174.035 ;
        RECT 134.675 173.705 134.940 174.265 ;
        RECT 135.110 173.535 135.280 174.435 ;
        RECT 136.585 174.395 136.755 174.685 ;
        RECT 136.925 174.565 137.255 174.945 ;
        RECT 135.450 173.705 135.805 174.265 ;
        RECT 136.585 174.225 137.250 174.395 ;
        RECT 134.255 173.365 135.680 173.535 ;
        RECT 136.500 173.405 136.850 174.055 ;
        RECT 133.770 172.565 134.305 173.185 ;
        RECT 134.475 172.395 134.805 173.195 ;
        RECT 135.290 173.190 135.680 173.365 ;
        RECT 137.020 173.235 137.250 174.225 ;
        RECT 136.585 173.065 137.250 173.235 ;
        RECT 136.585 172.565 136.755 173.065 ;
        RECT 136.925 172.395 137.255 172.895 ;
        RECT 137.425 172.565 137.610 174.685 ;
        RECT 137.865 174.485 138.115 174.945 ;
        RECT 138.285 174.495 138.620 174.665 ;
        RECT 138.815 174.495 139.490 174.665 ;
        RECT 138.285 174.355 138.455 174.495 ;
        RECT 137.780 173.365 138.060 174.315 ;
        RECT 138.230 174.225 138.455 174.355 ;
        RECT 138.230 173.120 138.400 174.225 ;
        RECT 138.625 174.075 139.150 174.295 ;
        RECT 138.570 173.310 138.810 173.905 ;
        RECT 138.980 173.375 139.150 174.075 ;
        RECT 139.320 173.715 139.490 174.495 ;
        RECT 139.810 174.445 140.180 174.945 ;
        RECT 140.360 174.495 140.765 174.665 ;
        RECT 140.935 174.495 141.720 174.665 ;
        RECT 140.360 174.265 140.530 174.495 ;
        RECT 139.700 173.965 140.530 174.265 ;
        RECT 140.915 173.995 141.380 174.325 ;
        RECT 139.700 173.935 139.900 173.965 ;
        RECT 140.020 173.715 140.190 173.785 ;
        RECT 139.320 173.545 140.190 173.715 ;
        RECT 139.680 173.455 140.190 173.545 ;
        RECT 138.230 172.990 138.535 173.120 ;
        RECT 138.980 173.010 139.510 173.375 ;
        RECT 137.850 172.395 138.115 172.855 ;
        RECT 138.285 172.565 138.535 172.990 ;
        RECT 139.680 172.840 139.850 173.455 ;
        RECT 138.745 172.670 139.850 172.840 ;
        RECT 140.020 172.395 140.190 173.195 ;
        RECT 140.360 172.895 140.530 173.965 ;
        RECT 140.700 173.065 140.890 173.785 ;
        RECT 141.060 173.035 141.380 173.995 ;
        RECT 141.550 174.035 141.720 174.495 ;
        RECT 141.995 174.415 142.205 174.945 ;
        RECT 142.465 174.205 142.795 174.730 ;
        RECT 142.965 174.335 143.135 174.945 ;
        RECT 143.305 174.290 143.635 174.725 ;
        RECT 143.945 174.395 144.115 174.775 ;
        RECT 144.330 174.565 144.660 174.945 ;
        RECT 143.305 174.205 143.685 174.290 ;
        RECT 143.945 174.225 144.660 174.395 ;
        RECT 142.595 174.035 142.795 174.205 ;
        RECT 143.460 174.165 143.685 174.205 ;
        RECT 141.550 173.705 142.425 174.035 ;
        RECT 142.595 173.705 143.345 174.035 ;
        RECT 140.360 172.565 140.610 172.895 ;
        RECT 141.550 172.865 141.720 173.705 ;
        RECT 142.595 173.500 142.785 173.705 ;
        RECT 143.515 173.585 143.685 174.165 ;
        RECT 143.855 173.675 144.210 174.045 ;
        RECT 144.490 174.035 144.660 174.225 ;
        RECT 144.830 174.200 145.085 174.775 ;
        RECT 144.490 173.705 144.745 174.035 ;
        RECT 143.470 173.535 143.685 173.585 ;
        RECT 141.890 173.125 142.785 173.500 ;
        RECT 143.295 173.455 143.685 173.535 ;
        RECT 144.490 173.495 144.660 173.705 ;
        RECT 140.835 172.695 141.720 172.865 ;
        RECT 141.900 172.395 142.215 172.895 ;
        RECT 142.445 172.565 142.785 173.125 ;
        RECT 142.955 172.395 143.125 173.405 ;
        RECT 143.295 172.610 143.625 173.455 ;
        RECT 143.945 173.325 144.660 173.495 ;
        RECT 144.915 173.470 145.085 174.200 ;
        RECT 145.260 174.105 145.520 174.945 ;
        RECT 145.695 174.195 146.905 174.945 ;
        RECT 143.945 172.565 144.115 173.325 ;
        RECT 144.330 172.395 144.660 173.155 ;
        RECT 144.830 172.565 145.085 173.470 ;
        RECT 145.260 172.395 145.520 173.545 ;
        RECT 145.695 173.485 146.215 174.025 ;
        RECT 146.385 173.655 146.905 174.195 ;
        RECT 145.695 172.395 146.905 173.485 ;
        RECT 17.270 172.225 146.990 172.395 ;
        RECT 17.355 171.135 18.565 172.225 ;
        RECT 19.285 171.555 19.455 172.055 ;
        RECT 19.625 171.725 19.955 172.225 ;
        RECT 19.285 171.385 19.950 171.555 ;
        RECT 17.355 170.425 17.875 170.965 ;
        RECT 18.045 170.595 18.565 171.135 ;
        RECT 19.200 170.565 19.550 171.215 ;
        RECT 17.355 169.675 18.565 170.425 ;
        RECT 19.720 170.395 19.950 171.385 ;
        RECT 19.285 170.225 19.950 170.395 ;
        RECT 19.285 169.935 19.455 170.225 ;
        RECT 19.625 169.675 19.955 170.055 ;
        RECT 20.125 169.935 20.310 172.055 ;
        RECT 20.550 171.765 20.815 172.225 ;
        RECT 20.985 171.630 21.235 172.055 ;
        RECT 21.445 171.780 22.550 171.950 ;
        RECT 20.930 171.500 21.235 171.630 ;
        RECT 20.480 170.305 20.760 171.255 ;
        RECT 20.930 170.395 21.100 171.500 ;
        RECT 21.270 170.715 21.510 171.310 ;
        RECT 21.680 171.245 22.210 171.610 ;
        RECT 21.680 170.545 21.850 171.245 ;
        RECT 22.380 171.165 22.550 171.780 ;
        RECT 22.720 171.425 22.890 172.225 ;
        RECT 23.060 171.725 23.310 172.055 ;
        RECT 23.535 171.755 24.420 171.925 ;
        RECT 22.380 171.075 22.890 171.165 ;
        RECT 20.930 170.265 21.155 170.395 ;
        RECT 21.325 170.325 21.850 170.545 ;
        RECT 22.020 170.905 22.890 171.075 ;
        RECT 20.565 169.675 20.815 170.135 ;
        RECT 20.985 170.125 21.155 170.265 ;
        RECT 22.020 170.125 22.190 170.905 ;
        RECT 22.720 170.835 22.890 170.905 ;
        RECT 22.400 170.655 22.600 170.685 ;
        RECT 23.060 170.655 23.230 171.725 ;
        RECT 23.400 170.835 23.590 171.555 ;
        RECT 22.400 170.355 23.230 170.655 ;
        RECT 23.760 170.625 24.080 171.585 ;
        RECT 20.985 169.955 21.320 170.125 ;
        RECT 21.515 169.955 22.190 170.125 ;
        RECT 22.510 169.675 22.880 170.175 ;
        RECT 23.060 170.125 23.230 170.355 ;
        RECT 23.615 170.295 24.080 170.625 ;
        RECT 24.250 170.915 24.420 171.755 ;
        RECT 24.600 171.725 24.915 172.225 ;
        RECT 25.145 171.495 25.485 172.055 ;
        RECT 24.590 171.120 25.485 171.495 ;
        RECT 25.655 171.215 25.825 172.225 ;
        RECT 25.295 170.915 25.485 171.120 ;
        RECT 25.995 171.165 26.325 172.010 ;
        RECT 25.995 171.085 26.385 171.165 ;
        RECT 26.555 171.085 26.815 172.225 ;
        RECT 26.170 171.035 26.385 171.085 ;
        RECT 26.985 171.075 27.315 172.055 ;
        RECT 27.485 171.085 27.765 172.225 ;
        RECT 27.935 171.670 28.540 172.225 ;
        RECT 28.715 171.715 29.195 172.055 ;
        RECT 29.365 171.680 29.620 172.225 ;
        RECT 27.935 171.570 28.550 171.670 ;
        RECT 28.365 171.545 28.550 171.570 ;
        RECT 24.250 170.585 25.125 170.915 ;
        RECT 25.295 170.585 26.045 170.915 ;
        RECT 24.250 170.125 24.420 170.585 ;
        RECT 25.295 170.415 25.495 170.585 ;
        RECT 26.215 170.455 26.385 171.035 ;
        RECT 26.575 170.665 26.910 170.915 ;
        RECT 27.080 170.475 27.250 171.075 ;
        RECT 27.935 170.950 28.195 171.400 ;
        RECT 28.365 171.300 28.695 171.545 ;
        RECT 28.865 171.225 29.620 171.475 ;
        RECT 29.790 171.355 30.065 172.055 ;
        RECT 28.850 171.190 29.620 171.225 ;
        RECT 28.835 171.180 29.620 171.190 ;
        RECT 28.830 171.165 29.725 171.180 ;
        RECT 28.810 171.150 29.725 171.165 ;
        RECT 28.790 171.140 29.725 171.150 ;
        RECT 28.765 171.130 29.725 171.140 ;
        RECT 28.695 171.100 29.725 171.130 ;
        RECT 28.675 171.070 29.725 171.100 ;
        RECT 28.655 171.040 29.725 171.070 ;
        RECT 28.625 171.015 29.725 171.040 ;
        RECT 28.590 170.980 29.725 171.015 ;
        RECT 28.560 170.975 29.725 170.980 ;
        RECT 28.560 170.970 28.950 170.975 ;
        RECT 28.560 170.960 28.925 170.970 ;
        RECT 28.560 170.955 28.910 170.960 ;
        RECT 28.560 170.950 28.895 170.955 ;
        RECT 27.935 170.945 28.895 170.950 ;
        RECT 27.935 170.935 28.885 170.945 ;
        RECT 27.935 170.930 28.875 170.935 ;
        RECT 27.935 170.920 28.865 170.930 ;
        RECT 27.420 170.645 27.755 170.915 ;
        RECT 27.935 170.910 28.860 170.920 ;
        RECT 27.935 170.905 28.855 170.910 ;
        RECT 27.935 170.890 28.845 170.905 ;
        RECT 27.935 170.875 28.840 170.890 ;
        RECT 27.935 170.850 28.830 170.875 ;
        RECT 27.935 170.780 28.825 170.850 ;
        RECT 26.160 170.415 26.385 170.455 ;
        RECT 23.060 169.955 23.465 170.125 ;
        RECT 23.635 169.955 24.420 170.125 ;
        RECT 24.695 169.675 24.905 170.205 ;
        RECT 25.165 169.890 25.495 170.415 ;
        RECT 26.005 170.330 26.385 170.415 ;
        RECT 25.665 169.675 25.835 170.285 ;
        RECT 26.005 169.895 26.335 170.330 ;
        RECT 26.555 169.845 27.250 170.475 ;
        RECT 27.455 169.675 27.765 170.475 ;
        RECT 27.935 170.225 28.485 170.610 ;
        RECT 28.655 170.055 28.825 170.780 ;
        RECT 27.935 169.885 28.825 170.055 ;
        RECT 28.995 170.380 29.325 170.805 ;
        RECT 29.495 170.580 29.725 170.975 ;
        RECT 28.995 169.895 29.215 170.380 ;
        RECT 29.895 170.325 30.065 171.355 ;
        RECT 30.235 171.060 30.525 172.225 ;
        RECT 30.785 171.555 30.955 172.055 ;
        RECT 31.125 171.725 31.455 172.225 ;
        RECT 30.785 171.385 31.450 171.555 ;
        RECT 30.700 170.565 31.050 171.215 ;
        RECT 29.385 169.675 29.635 170.215 ;
        RECT 29.805 169.845 30.065 170.325 ;
        RECT 30.235 169.675 30.525 170.400 ;
        RECT 31.220 170.395 31.450 171.385 ;
        RECT 30.785 170.225 31.450 170.395 ;
        RECT 30.785 169.935 30.955 170.225 ;
        RECT 31.125 169.675 31.455 170.055 ;
        RECT 31.625 169.935 31.810 172.055 ;
        RECT 32.050 171.765 32.315 172.225 ;
        RECT 32.485 171.630 32.735 172.055 ;
        RECT 32.945 171.780 34.050 171.950 ;
        RECT 32.430 171.500 32.735 171.630 ;
        RECT 31.980 170.305 32.260 171.255 ;
        RECT 32.430 170.395 32.600 171.500 ;
        RECT 32.770 170.715 33.010 171.310 ;
        RECT 33.180 171.245 33.710 171.610 ;
        RECT 33.180 170.545 33.350 171.245 ;
        RECT 33.880 171.165 34.050 171.780 ;
        RECT 34.220 171.425 34.390 172.225 ;
        RECT 34.560 171.725 34.810 172.055 ;
        RECT 35.035 171.755 35.920 171.925 ;
        RECT 33.880 171.075 34.390 171.165 ;
        RECT 32.430 170.265 32.655 170.395 ;
        RECT 32.825 170.325 33.350 170.545 ;
        RECT 33.520 170.905 34.390 171.075 ;
        RECT 32.065 169.675 32.315 170.135 ;
        RECT 32.485 170.125 32.655 170.265 ;
        RECT 33.520 170.125 33.690 170.905 ;
        RECT 34.220 170.835 34.390 170.905 ;
        RECT 33.900 170.655 34.100 170.685 ;
        RECT 34.560 170.655 34.730 171.725 ;
        RECT 34.900 170.835 35.090 171.555 ;
        RECT 33.900 170.355 34.730 170.655 ;
        RECT 35.260 170.625 35.580 171.585 ;
        RECT 32.485 169.955 32.820 170.125 ;
        RECT 33.015 169.955 33.690 170.125 ;
        RECT 34.010 169.675 34.380 170.175 ;
        RECT 34.560 170.125 34.730 170.355 ;
        RECT 35.115 170.295 35.580 170.625 ;
        RECT 35.750 170.915 35.920 171.755 ;
        RECT 36.100 171.725 36.415 172.225 ;
        RECT 36.645 171.495 36.985 172.055 ;
        RECT 36.090 171.120 36.985 171.495 ;
        RECT 37.155 171.215 37.325 172.225 ;
        RECT 36.795 170.915 36.985 171.120 ;
        RECT 37.495 171.165 37.825 172.010 ;
        RECT 38.255 171.555 38.535 172.225 ;
        RECT 38.705 171.335 39.005 171.885 ;
        RECT 39.205 171.505 39.535 172.225 ;
        RECT 39.725 171.505 40.185 172.055 ;
        RECT 40.360 171.800 40.695 172.225 ;
        RECT 40.865 171.620 41.050 172.025 ;
        RECT 37.495 171.085 37.885 171.165 ;
        RECT 37.670 171.035 37.885 171.085 ;
        RECT 35.750 170.585 36.625 170.915 ;
        RECT 36.795 170.585 37.545 170.915 ;
        RECT 35.750 170.125 35.920 170.585 ;
        RECT 36.795 170.415 36.995 170.585 ;
        RECT 37.715 170.455 37.885 171.035 ;
        RECT 38.070 170.915 38.335 171.275 ;
        RECT 38.705 171.165 39.645 171.335 ;
        RECT 39.475 170.915 39.645 171.165 ;
        RECT 38.070 170.665 38.745 170.915 ;
        RECT 38.965 170.665 39.305 170.915 ;
        RECT 39.475 170.585 39.765 170.915 ;
        RECT 39.475 170.495 39.645 170.585 ;
        RECT 37.660 170.415 37.885 170.455 ;
        RECT 34.560 169.955 34.965 170.125 ;
        RECT 35.135 169.955 35.920 170.125 ;
        RECT 36.195 169.675 36.405 170.205 ;
        RECT 36.665 169.890 36.995 170.415 ;
        RECT 37.505 170.330 37.885 170.415 ;
        RECT 37.165 169.675 37.335 170.285 ;
        RECT 37.505 169.895 37.835 170.330 ;
        RECT 38.255 170.305 39.645 170.495 ;
        RECT 38.255 169.945 38.585 170.305 ;
        RECT 39.935 170.135 40.185 171.505 ;
        RECT 40.385 171.445 41.050 171.620 ;
        RECT 41.255 171.445 41.585 172.225 ;
        RECT 40.385 170.415 40.725 171.445 ;
        RECT 41.755 171.255 42.025 172.025 ;
        RECT 40.895 171.085 42.025 171.255 ;
        RECT 42.380 171.255 42.770 171.430 ;
        RECT 43.255 171.425 43.585 172.225 ;
        RECT 43.755 171.435 44.290 172.055 ;
        RECT 44.495 171.670 45.100 172.225 ;
        RECT 45.275 171.715 45.755 172.055 ;
        RECT 45.925 171.680 46.180 172.225 ;
        RECT 44.495 171.570 45.110 171.670 ;
        RECT 42.380 171.085 43.805 171.255 ;
        RECT 40.895 170.585 41.145 171.085 ;
        RECT 40.385 170.245 41.070 170.415 ;
        RECT 41.325 170.335 41.685 170.915 ;
        RECT 39.205 169.675 39.455 170.135 ;
        RECT 39.625 169.845 40.185 170.135 ;
        RECT 40.360 169.675 40.695 170.075 ;
        RECT 40.865 169.845 41.070 170.245 ;
        RECT 41.855 170.175 42.025 171.085 ;
        RECT 42.255 170.355 42.610 170.915 ;
        RECT 42.780 170.185 42.950 171.085 ;
        RECT 43.120 170.355 43.385 170.915 ;
        RECT 43.635 170.585 43.805 171.085 ;
        RECT 43.975 170.415 44.290 171.435 ;
        RECT 44.925 171.545 45.110 171.570 ;
        RECT 44.495 170.950 44.755 171.400 ;
        RECT 44.925 171.300 45.255 171.545 ;
        RECT 45.425 171.225 46.180 171.475 ;
        RECT 46.350 171.355 46.625 172.055 ;
        RECT 46.795 171.715 47.095 172.225 ;
        RECT 47.265 171.545 47.595 172.055 ;
        RECT 47.765 171.715 48.395 172.225 ;
        RECT 48.975 171.715 49.355 171.885 ;
        RECT 49.525 171.715 49.825 172.225 ;
        RECT 49.185 171.545 49.355 171.715 ;
        RECT 50.215 171.555 50.495 172.225 ;
        RECT 45.410 171.190 46.180 171.225 ;
        RECT 45.395 171.180 46.180 171.190 ;
        RECT 45.390 171.165 46.285 171.180 ;
        RECT 45.370 171.150 46.285 171.165 ;
        RECT 45.350 171.140 46.285 171.150 ;
        RECT 45.325 171.130 46.285 171.140 ;
        RECT 45.255 171.100 46.285 171.130 ;
        RECT 45.235 171.070 46.285 171.100 ;
        RECT 45.215 171.040 46.285 171.070 ;
        RECT 45.185 171.015 46.285 171.040 ;
        RECT 45.150 170.980 46.285 171.015 ;
        RECT 45.120 170.975 46.285 170.980 ;
        RECT 45.120 170.970 45.510 170.975 ;
        RECT 45.120 170.960 45.485 170.970 ;
        RECT 45.120 170.955 45.470 170.960 ;
        RECT 45.120 170.950 45.455 170.955 ;
        RECT 44.495 170.945 45.455 170.950 ;
        RECT 44.495 170.935 45.445 170.945 ;
        RECT 44.495 170.930 45.435 170.935 ;
        RECT 44.495 170.920 45.425 170.930 ;
        RECT 44.495 170.910 45.420 170.920 ;
        RECT 44.495 170.905 45.415 170.910 ;
        RECT 44.495 170.890 45.405 170.905 ;
        RECT 44.495 170.875 45.400 170.890 ;
        RECT 44.495 170.850 45.390 170.875 ;
        RECT 44.495 170.780 45.385 170.850 ;
        RECT 41.280 169.675 41.555 170.155 ;
        RECT 41.765 169.845 42.025 170.175 ;
        RECT 42.360 169.675 42.600 170.185 ;
        RECT 42.780 169.855 43.060 170.185 ;
        RECT 43.290 169.675 43.505 170.185 ;
        RECT 43.675 169.845 44.290 170.415 ;
        RECT 44.495 170.225 45.045 170.610 ;
        RECT 45.215 170.055 45.385 170.780 ;
        RECT 44.495 169.885 45.385 170.055 ;
        RECT 45.555 170.380 45.885 170.805 ;
        RECT 46.055 170.580 46.285 170.975 ;
        RECT 45.555 169.895 45.775 170.380 ;
        RECT 46.455 170.325 46.625 171.355 ;
        RECT 45.945 169.675 46.195 170.215 ;
        RECT 46.365 169.845 46.625 170.325 ;
        RECT 46.795 171.375 49.015 171.545 ;
        RECT 46.795 170.415 46.965 171.375 ;
        RECT 47.135 171.035 48.675 171.205 ;
        RECT 47.135 170.585 47.380 171.035 ;
        RECT 47.640 170.665 48.335 170.865 ;
        RECT 48.505 170.835 48.675 171.035 ;
        RECT 48.845 171.175 49.015 171.375 ;
        RECT 49.185 171.345 49.845 171.545 ;
        RECT 48.845 171.005 49.505 171.175 ;
        RECT 48.505 170.665 49.105 170.835 ;
        RECT 49.335 170.585 49.505 171.005 ;
        RECT 46.795 169.870 47.260 170.415 ;
        RECT 47.765 169.675 47.935 170.495 ;
        RECT 48.105 170.415 49.015 170.495 ;
        RECT 49.675 170.415 49.845 171.345 ;
        RECT 50.665 171.335 50.965 171.885 ;
        RECT 51.165 171.505 51.495 172.225 ;
        RECT 51.685 171.505 52.145 172.055 ;
        RECT 50.030 170.915 50.295 171.275 ;
        RECT 50.665 171.165 51.605 171.335 ;
        RECT 51.435 170.915 51.605 171.165 ;
        RECT 50.030 170.665 50.705 170.915 ;
        RECT 50.925 170.665 51.265 170.915 ;
        RECT 51.435 170.585 51.725 170.915 ;
        RECT 51.435 170.495 51.605 170.585 ;
        RECT 48.105 170.325 49.355 170.415 ;
        RECT 48.105 169.845 48.435 170.325 ;
        RECT 48.845 170.245 49.355 170.325 ;
        RECT 48.605 169.675 48.955 170.065 ;
        RECT 49.125 169.845 49.355 170.245 ;
        RECT 49.525 169.935 49.845 170.415 ;
        RECT 50.215 170.305 51.605 170.495 ;
        RECT 50.215 169.945 50.545 170.305 ;
        RECT 51.895 170.135 52.145 171.505 ;
        RECT 52.315 171.135 55.825 172.225 ;
        RECT 51.165 169.675 51.415 170.135 ;
        RECT 51.585 169.845 52.145 170.135 ;
        RECT 52.315 170.445 53.965 170.965 ;
        RECT 54.135 170.615 55.825 171.135 ;
        RECT 55.995 171.060 56.285 172.225 ;
        RECT 56.455 171.790 61.800 172.225 ;
        RECT 61.975 171.790 67.320 172.225 ;
        RECT 67.495 171.790 72.840 172.225 ;
        RECT 73.015 171.790 78.360 172.225 ;
        RECT 52.315 169.675 55.825 170.445 ;
        RECT 55.995 169.675 56.285 170.400 ;
        RECT 58.040 170.220 58.380 171.050 ;
        RECT 59.860 170.540 60.210 171.790 ;
        RECT 63.560 170.220 63.900 171.050 ;
        RECT 65.380 170.540 65.730 171.790 ;
        RECT 69.080 170.220 69.420 171.050 ;
        RECT 70.900 170.540 71.250 171.790 ;
        RECT 74.600 170.220 74.940 171.050 ;
        RECT 76.420 170.540 76.770 171.790 ;
        RECT 78.535 171.135 81.125 172.225 ;
        RECT 78.535 170.445 79.745 170.965 ;
        RECT 79.915 170.615 81.125 171.135 ;
        RECT 81.755 171.060 82.045 172.225 ;
        RECT 82.675 170.935 82.945 172.035 ;
        RECT 83.115 171.295 83.390 171.800 ;
        RECT 83.560 171.465 83.890 172.225 ;
        RECT 83.115 171.125 83.605 171.295 ;
        RECT 84.060 171.215 84.385 172.055 ;
        RECT 82.675 170.585 83.125 170.935 ;
        RECT 83.310 170.585 83.605 171.125 ;
        RECT 83.775 171.045 84.385 171.215 ;
        RECT 84.860 171.125 85.235 172.225 ;
        RECT 85.435 171.715 85.695 172.225 ;
        RECT 56.455 169.675 61.800 170.220 ;
        RECT 61.975 169.675 67.320 170.220 ;
        RECT 67.495 169.675 72.840 170.220 ;
        RECT 73.015 169.675 78.360 170.220 ;
        RECT 78.535 169.675 81.125 170.445 ;
        RECT 83.310 170.415 83.480 170.585 ;
        RECT 83.775 170.415 83.945 171.045 ;
        RECT 84.115 170.665 84.615 170.875 ;
        RECT 84.785 170.665 85.265 170.875 ;
        RECT 85.435 170.665 85.775 171.545 ;
        RECT 85.945 170.835 86.115 172.055 ;
        RECT 86.355 171.720 86.970 172.225 ;
        RECT 86.355 171.185 86.605 171.550 ;
        RECT 86.775 171.545 86.970 171.720 ;
        RECT 87.140 171.715 87.615 172.055 ;
        RECT 87.785 171.680 88.000 172.225 ;
        RECT 86.775 171.355 87.105 171.545 ;
        RECT 87.325 171.185 88.040 171.480 ;
        RECT 88.210 171.355 88.485 172.055 ;
        RECT 86.355 171.015 88.145 171.185 ;
        RECT 85.945 170.585 86.740 170.835 ;
        RECT 85.945 170.495 86.195 170.585 ;
        RECT 81.755 169.675 82.045 170.400 ;
        RECT 82.675 169.675 82.950 170.415 ;
        RECT 83.170 170.245 83.480 170.415 ;
        RECT 83.170 170.085 83.360 170.245 ;
        RECT 83.705 170.235 83.945 170.415 ;
        RECT 84.160 170.325 85.255 170.495 ;
        RECT 83.705 169.845 83.875 170.235 ;
        RECT 84.160 170.075 84.330 170.325 ;
        RECT 84.080 169.845 84.410 170.075 ;
        RECT 84.585 169.675 84.755 170.145 ;
        RECT 84.925 169.860 85.255 170.325 ;
        RECT 85.435 169.675 85.695 170.495 ;
        RECT 85.865 170.075 86.195 170.495 ;
        RECT 86.910 170.160 87.165 171.015 ;
        RECT 86.375 169.895 87.165 170.160 ;
        RECT 87.335 170.315 87.745 170.835 ;
        RECT 87.915 170.585 88.145 171.015 ;
        RECT 88.315 170.325 88.485 171.355 ;
        RECT 88.655 171.085 88.915 172.225 ;
        RECT 89.085 171.075 89.415 172.055 ;
        RECT 89.585 171.085 89.865 172.225 ;
        RECT 90.585 171.555 90.755 172.055 ;
        RECT 90.925 171.725 91.255 172.225 ;
        RECT 90.585 171.385 91.250 171.555 ;
        RECT 88.675 170.665 89.010 170.915 ;
        RECT 89.180 170.475 89.350 171.075 ;
        RECT 89.520 170.645 89.855 170.915 ;
        RECT 90.500 170.565 90.850 171.215 ;
        RECT 87.335 169.895 87.535 170.315 ;
        RECT 87.725 169.675 88.055 170.135 ;
        RECT 88.225 169.845 88.485 170.325 ;
        RECT 88.655 169.845 89.350 170.475 ;
        RECT 89.555 169.675 89.865 170.475 ;
        RECT 91.020 170.395 91.250 171.385 ;
        RECT 90.585 170.225 91.250 170.395 ;
        RECT 90.585 169.935 90.755 170.225 ;
        RECT 90.925 169.675 91.255 170.055 ;
        RECT 91.425 169.935 91.610 172.055 ;
        RECT 91.850 171.765 92.115 172.225 ;
        RECT 92.285 171.630 92.535 172.055 ;
        RECT 92.745 171.780 93.850 171.950 ;
        RECT 92.230 171.500 92.535 171.630 ;
        RECT 91.780 170.305 92.060 171.255 ;
        RECT 92.230 170.395 92.400 171.500 ;
        RECT 92.570 170.715 92.810 171.310 ;
        RECT 92.980 171.245 93.510 171.610 ;
        RECT 92.980 170.545 93.150 171.245 ;
        RECT 93.680 171.165 93.850 171.780 ;
        RECT 94.020 171.425 94.190 172.225 ;
        RECT 94.360 171.725 94.610 172.055 ;
        RECT 94.835 171.755 95.720 171.925 ;
        RECT 93.680 171.075 94.190 171.165 ;
        RECT 92.230 170.265 92.455 170.395 ;
        RECT 92.625 170.325 93.150 170.545 ;
        RECT 93.320 170.905 94.190 171.075 ;
        RECT 91.865 169.675 92.115 170.135 ;
        RECT 92.285 170.125 92.455 170.265 ;
        RECT 93.320 170.125 93.490 170.905 ;
        RECT 94.020 170.835 94.190 170.905 ;
        RECT 93.700 170.655 93.900 170.685 ;
        RECT 94.360 170.655 94.530 171.725 ;
        RECT 94.700 170.835 94.890 171.555 ;
        RECT 93.700 170.355 94.530 170.655 ;
        RECT 95.060 170.625 95.380 171.585 ;
        RECT 92.285 169.955 92.620 170.125 ;
        RECT 92.815 169.955 93.490 170.125 ;
        RECT 93.810 169.675 94.180 170.175 ;
        RECT 94.360 170.125 94.530 170.355 ;
        RECT 94.915 170.295 95.380 170.625 ;
        RECT 95.550 170.915 95.720 171.755 ;
        RECT 95.900 171.725 96.215 172.225 ;
        RECT 96.445 171.495 96.785 172.055 ;
        RECT 95.890 171.120 96.785 171.495 ;
        RECT 96.955 171.215 97.125 172.225 ;
        RECT 96.595 170.915 96.785 171.120 ;
        RECT 97.295 171.165 97.625 172.010 ;
        RECT 98.105 171.495 98.400 172.225 ;
        RECT 98.570 171.325 98.830 172.050 ;
        RECT 99.000 171.495 99.260 172.225 ;
        RECT 99.430 171.325 99.690 172.050 ;
        RECT 99.860 171.495 100.120 172.225 ;
        RECT 100.290 171.325 100.550 172.050 ;
        RECT 100.720 171.495 100.980 172.225 ;
        RECT 101.150 171.325 101.410 172.050 ;
        RECT 97.295 171.085 97.685 171.165 ;
        RECT 97.470 171.035 97.685 171.085 ;
        RECT 95.550 170.585 96.425 170.915 ;
        RECT 96.595 170.585 97.345 170.915 ;
        RECT 95.550 170.125 95.720 170.585 ;
        RECT 96.595 170.415 96.795 170.585 ;
        RECT 97.515 170.455 97.685 171.035 ;
        RECT 97.460 170.415 97.685 170.455 ;
        RECT 94.360 169.955 94.765 170.125 ;
        RECT 94.935 169.955 95.720 170.125 ;
        RECT 95.995 169.675 96.205 170.205 ;
        RECT 96.465 169.890 96.795 170.415 ;
        RECT 97.305 170.330 97.685 170.415 ;
        RECT 98.100 171.085 101.410 171.325 ;
        RECT 101.580 171.115 101.840 172.225 ;
        RECT 98.100 170.495 99.070 171.085 ;
        RECT 102.010 170.915 102.260 172.050 ;
        RECT 102.440 171.115 102.735 172.225 ;
        RECT 102.915 171.085 103.300 172.055 ;
        RECT 103.470 171.765 103.795 172.225 ;
        RECT 104.315 171.595 104.595 172.055 ;
        RECT 103.470 171.375 104.595 171.595 ;
        RECT 99.240 170.665 102.260 170.915 ;
        RECT 96.965 169.675 97.135 170.285 ;
        RECT 97.305 169.895 97.635 170.330 ;
        RECT 98.100 170.325 101.410 170.495 ;
        RECT 98.100 169.675 98.400 170.155 ;
        RECT 98.570 169.870 98.830 170.325 ;
        RECT 99.000 169.675 99.260 170.155 ;
        RECT 99.430 169.870 99.690 170.325 ;
        RECT 99.860 169.675 100.120 170.155 ;
        RECT 100.290 169.870 100.550 170.325 ;
        RECT 100.720 169.675 100.980 170.155 ;
        RECT 101.150 169.870 101.410 170.325 ;
        RECT 101.580 169.675 101.840 170.200 ;
        RECT 102.010 169.855 102.260 170.665 ;
        RECT 102.430 170.305 102.745 170.915 ;
        RECT 102.915 170.415 103.195 171.085 ;
        RECT 103.470 170.915 103.920 171.375 ;
        RECT 104.785 171.205 105.185 172.055 ;
        RECT 105.585 171.765 105.855 172.225 ;
        RECT 106.025 171.595 106.310 172.055 ;
        RECT 103.365 170.585 103.920 170.915 ;
        RECT 104.090 170.645 105.185 171.205 ;
        RECT 103.470 170.475 103.920 170.585 ;
        RECT 102.440 169.675 102.685 170.135 ;
        RECT 102.915 169.845 103.300 170.415 ;
        RECT 103.470 170.305 104.595 170.475 ;
        RECT 103.470 169.675 103.795 170.135 ;
        RECT 104.315 169.845 104.595 170.305 ;
        RECT 104.785 169.845 105.185 170.645 ;
        RECT 105.355 171.375 106.310 171.595 ;
        RECT 105.355 170.475 105.565 171.375 ;
        RECT 105.735 170.645 106.425 171.205 ;
        RECT 107.515 171.060 107.805 172.225 ;
        RECT 108.020 171.085 108.315 172.225 ;
        RECT 108.575 171.255 108.905 172.055 ;
        RECT 109.075 171.425 109.245 172.225 ;
        RECT 109.415 171.255 109.745 172.055 ;
        RECT 109.915 171.425 110.085 172.225 ;
        RECT 110.255 171.275 110.585 172.055 ;
        RECT 110.755 171.765 110.925 172.225 ;
        RECT 111.195 171.715 111.455 172.225 ;
        RECT 110.255 171.255 111.025 171.275 ;
        RECT 108.575 171.085 111.025 171.255 ;
        RECT 107.995 170.665 110.505 170.915 ;
        RECT 110.675 170.495 111.025 171.085 ;
        RECT 111.195 170.665 111.535 171.545 ;
        RECT 111.705 170.835 111.875 172.055 ;
        RECT 112.115 171.720 112.730 172.225 ;
        RECT 112.115 171.185 112.365 171.550 ;
        RECT 112.535 171.545 112.730 171.720 ;
        RECT 112.900 171.715 113.375 172.055 ;
        RECT 113.545 171.680 113.760 172.225 ;
        RECT 112.535 171.355 112.865 171.545 ;
        RECT 113.085 171.185 113.800 171.480 ;
        RECT 113.970 171.355 114.245 172.055 ;
        RECT 114.455 171.885 115.595 172.055 ;
        RECT 114.455 171.425 114.755 171.885 ;
        RECT 112.115 171.015 113.905 171.185 ;
        RECT 111.705 170.585 112.500 170.835 ;
        RECT 111.705 170.495 111.955 170.585 ;
        RECT 105.355 170.305 106.310 170.475 ;
        RECT 105.585 169.675 105.855 170.135 ;
        RECT 106.025 169.845 106.310 170.305 ;
        RECT 107.515 169.675 107.805 170.400 ;
        RECT 108.655 170.315 111.025 170.495 ;
        RECT 108.020 169.675 108.285 170.135 ;
        RECT 108.655 169.845 108.825 170.315 ;
        RECT 109.075 169.675 109.245 170.135 ;
        RECT 109.495 169.845 109.665 170.315 ;
        RECT 109.915 169.675 110.085 170.135 ;
        RECT 110.335 169.845 110.505 170.315 ;
        RECT 110.675 169.675 110.925 170.140 ;
        RECT 111.195 169.675 111.455 170.495 ;
        RECT 111.625 170.075 111.955 170.495 ;
        RECT 112.670 170.160 112.925 171.015 ;
        RECT 112.135 169.895 112.925 170.160 ;
        RECT 113.095 170.315 113.505 170.835 ;
        RECT 113.675 170.585 113.905 171.015 ;
        RECT 114.075 170.325 114.245 171.355 ;
        RECT 114.925 171.255 115.255 171.715 ;
        RECT 114.495 171.205 115.255 171.255 ;
        RECT 114.475 171.035 115.255 171.205 ;
        RECT 115.425 171.255 115.595 171.885 ;
        RECT 115.765 171.425 116.095 172.225 ;
        RECT 116.265 171.255 116.540 172.055 ;
        RECT 115.425 171.045 116.540 171.255 ;
        RECT 114.495 170.495 114.710 171.035 ;
        RECT 114.880 170.665 115.650 170.865 ;
        RECT 115.820 170.665 116.540 170.865 ;
        RECT 114.495 170.325 116.095 170.495 ;
        RECT 113.095 169.895 113.295 170.315 ;
        RECT 113.485 169.675 113.815 170.135 ;
        RECT 113.985 169.845 114.245 170.325 ;
        RECT 114.925 170.315 116.095 170.325 ;
        RECT 114.465 169.675 114.755 170.145 ;
        RECT 114.925 169.845 115.255 170.315 ;
        RECT 115.425 169.675 115.595 170.145 ;
        RECT 115.765 169.845 116.095 170.315 ;
        RECT 116.265 169.675 116.540 170.495 ;
        RECT 117.645 169.855 117.905 172.045 ;
        RECT 118.075 171.495 118.415 172.225 ;
        RECT 118.595 171.315 118.865 172.045 ;
        RECT 118.095 171.095 118.865 171.315 ;
        RECT 119.045 171.335 119.275 172.045 ;
        RECT 119.445 171.515 119.775 172.225 ;
        RECT 119.945 171.335 120.205 172.045 ;
        RECT 119.045 171.095 120.205 171.335 ;
        RECT 118.095 170.425 118.385 171.095 ;
        RECT 118.565 170.605 119.030 170.915 ;
        RECT 119.210 170.605 119.735 170.915 ;
        RECT 118.095 170.225 119.325 170.425 ;
        RECT 118.165 169.675 118.835 170.045 ;
        RECT 119.015 169.855 119.325 170.225 ;
        RECT 119.505 169.965 119.735 170.605 ;
        RECT 119.915 170.585 120.215 170.915 ;
        RECT 119.915 169.675 120.205 170.405 ;
        RECT 120.865 169.855 121.125 172.045 ;
        RECT 121.295 171.495 121.635 172.225 ;
        RECT 121.815 171.315 122.085 172.045 ;
        RECT 121.315 171.095 122.085 171.315 ;
        RECT 122.265 171.335 122.495 172.045 ;
        RECT 122.665 171.515 122.995 172.225 ;
        RECT 123.165 171.335 123.425 172.045 ;
        RECT 122.265 171.095 123.425 171.335 ;
        RECT 121.315 170.425 121.605 171.095 ;
        RECT 123.745 171.055 124.075 172.225 ;
        RECT 121.785 170.605 122.250 170.915 ;
        RECT 122.430 170.605 122.955 170.915 ;
        RECT 121.315 170.225 122.545 170.425 ;
        RECT 121.385 169.675 122.055 170.045 ;
        RECT 122.235 169.855 122.545 170.225 ;
        RECT 122.725 169.965 122.955 170.605 ;
        RECT 123.135 170.585 123.435 170.915 ;
        RECT 124.275 170.885 124.605 172.055 ;
        RECT 124.805 171.055 125.135 172.225 ;
        RECT 125.335 170.885 125.695 172.055 ;
        RECT 125.865 171.085 126.195 172.225 ;
        RECT 126.530 171.215 126.830 172.055 ;
        RECT 127.025 171.385 127.275 172.225 ;
        RECT 127.865 171.635 128.670 172.055 ;
        RECT 127.445 171.465 129.010 171.635 ;
        RECT 127.445 171.215 127.615 171.465 ;
        RECT 126.530 171.045 127.615 171.215 ;
        RECT 124.275 170.605 125.695 170.885 ;
        RECT 123.135 169.675 123.425 170.405 ;
        RECT 124.285 169.675 124.615 170.365 ;
        RECT 125.335 170.270 125.695 170.605 ;
        RECT 125.865 170.335 126.205 170.915 ;
        RECT 126.375 170.585 126.705 170.875 ;
        RECT 126.875 170.415 127.045 171.045 ;
        RECT 127.785 170.915 128.105 171.295 ;
        RECT 128.295 171.205 128.670 171.295 ;
        RECT 128.275 171.035 128.670 171.205 ;
        RECT 128.840 171.215 129.010 171.465 ;
        RECT 129.180 171.385 129.510 172.225 ;
        RECT 129.680 171.465 130.345 172.055 ;
        RECT 128.840 171.045 129.760 171.215 ;
        RECT 127.215 170.665 127.545 170.875 ;
        RECT 127.725 170.665 128.105 170.915 ;
        RECT 128.295 170.875 128.670 171.035 ;
        RECT 129.590 170.875 129.760 171.045 ;
        RECT 128.295 170.665 128.780 170.875 ;
        RECT 128.970 170.665 129.420 170.875 ;
        RECT 129.590 170.665 129.925 170.875 ;
        RECT 130.095 170.495 130.345 171.465 ;
        RECT 125.075 169.845 125.695 170.270 ;
        RECT 126.535 170.235 127.045 170.415 ;
        RECT 127.450 170.325 129.150 170.495 ;
        RECT 127.450 170.235 127.835 170.325 ;
        RECT 125.865 169.675 126.195 170.165 ;
        RECT 126.535 169.845 126.865 170.235 ;
        RECT 127.035 169.895 128.220 170.065 ;
        RECT 128.480 169.675 128.650 170.145 ;
        RECT 128.820 169.860 129.150 170.325 ;
        RECT 129.320 169.675 129.490 170.495 ;
        RECT 129.660 169.855 130.345 170.495 ;
        RECT 130.550 171.435 131.085 172.055 ;
        RECT 130.550 170.415 130.865 171.435 ;
        RECT 131.255 171.425 131.585 172.225 ;
        RECT 132.070 171.255 132.460 171.430 ;
        RECT 131.035 171.085 132.460 171.255 ;
        RECT 131.035 170.585 131.205 171.085 ;
        RECT 130.550 169.845 131.165 170.415 ;
        RECT 131.455 170.355 131.720 170.915 ;
        RECT 131.890 170.185 132.060 171.085 ;
        RECT 133.275 171.060 133.565 172.225 ;
        RECT 133.735 171.715 134.925 172.005 ;
        RECT 133.755 171.375 134.925 171.545 ;
        RECT 135.095 171.425 135.375 172.225 ;
        RECT 133.755 171.085 134.080 171.375 ;
        RECT 134.755 171.255 134.925 171.375 ;
        RECT 134.250 170.915 134.445 171.205 ;
        RECT 134.755 171.085 135.415 171.255 ;
        RECT 135.585 171.085 135.860 172.055 ;
        RECT 136.035 171.135 137.245 172.225 ;
        RECT 135.245 170.915 135.415 171.085 ;
        RECT 132.230 170.355 132.585 170.915 ;
        RECT 133.735 170.585 134.080 170.915 ;
        RECT 134.250 170.585 135.075 170.915 ;
        RECT 135.245 170.585 135.520 170.915 ;
        RECT 135.245 170.415 135.415 170.585 ;
        RECT 131.335 169.675 131.550 170.185 ;
        RECT 131.780 169.855 132.060 170.185 ;
        RECT 132.240 169.675 132.480 170.185 ;
        RECT 133.275 169.675 133.565 170.400 ;
        RECT 133.750 170.245 135.415 170.415 ;
        RECT 135.690 170.350 135.860 171.085 ;
        RECT 133.750 169.895 134.005 170.245 ;
        RECT 134.175 169.675 134.505 170.075 ;
        RECT 134.675 169.895 134.845 170.245 ;
        RECT 135.015 169.675 135.395 170.075 ;
        RECT 135.585 170.005 135.860 170.350 ;
        RECT 136.035 170.425 136.555 170.965 ;
        RECT 136.725 170.595 137.245 171.135 ;
        RECT 137.420 171.085 137.755 172.055 ;
        RECT 137.925 171.085 138.095 172.225 ;
        RECT 138.265 171.885 140.295 172.055 ;
        RECT 136.035 169.675 137.245 170.425 ;
        RECT 137.420 170.415 137.590 171.085 ;
        RECT 138.265 170.915 138.435 171.885 ;
        RECT 137.760 170.585 138.015 170.915 ;
        RECT 138.240 170.585 138.435 170.915 ;
        RECT 138.605 171.545 139.730 171.715 ;
        RECT 137.845 170.415 138.015 170.585 ;
        RECT 138.605 170.415 138.775 171.545 ;
        RECT 137.420 169.845 137.675 170.415 ;
        RECT 137.845 170.245 138.775 170.415 ;
        RECT 138.945 171.205 139.955 171.375 ;
        RECT 138.945 170.405 139.115 171.205 ;
        RECT 139.320 170.525 139.595 171.005 ;
        RECT 139.315 170.355 139.595 170.525 ;
        RECT 138.600 170.210 138.775 170.245 ;
        RECT 137.845 169.675 138.175 170.075 ;
        RECT 138.600 169.845 139.130 170.210 ;
        RECT 139.320 169.845 139.595 170.355 ;
        RECT 139.765 169.845 139.955 171.205 ;
        RECT 140.125 171.220 140.295 171.885 ;
        RECT 140.465 171.465 140.635 172.225 ;
        RECT 140.870 171.465 141.385 171.875 ;
        RECT 140.125 171.030 140.875 171.220 ;
        RECT 141.045 170.655 141.385 171.465 ;
        RECT 140.155 170.485 141.385 170.655 ;
        RECT 141.555 171.085 141.940 172.055 ;
        RECT 142.110 171.765 142.435 172.225 ;
        RECT 142.955 171.595 143.235 172.055 ;
        RECT 142.110 171.375 143.235 171.595 ;
        RECT 140.135 169.675 140.645 170.210 ;
        RECT 140.865 169.880 141.110 170.485 ;
        RECT 141.555 170.415 141.835 171.085 ;
        RECT 142.110 170.915 142.560 171.375 ;
        RECT 143.425 171.205 143.825 172.055 ;
        RECT 144.225 171.765 144.495 172.225 ;
        RECT 144.665 171.595 144.950 172.055 ;
        RECT 142.005 170.585 142.560 170.915 ;
        RECT 142.730 170.645 143.825 171.205 ;
        RECT 142.110 170.475 142.560 170.585 ;
        RECT 141.555 169.845 141.940 170.415 ;
        RECT 142.110 170.305 143.235 170.475 ;
        RECT 142.110 169.675 142.435 170.135 ;
        RECT 142.955 169.845 143.235 170.305 ;
        RECT 143.425 169.845 143.825 170.645 ;
        RECT 143.995 171.375 144.950 171.595 ;
        RECT 143.995 170.475 144.205 171.375 ;
        RECT 144.375 170.645 145.065 171.205 ;
        RECT 145.695 171.135 146.905 172.225 ;
        RECT 145.695 170.595 146.215 171.135 ;
        RECT 143.995 170.305 144.950 170.475 ;
        RECT 146.385 170.425 146.905 170.965 ;
        RECT 144.225 169.675 144.495 170.135 ;
        RECT 144.665 169.845 144.950 170.305 ;
        RECT 145.695 169.675 146.905 170.425 ;
        RECT 17.270 169.505 146.990 169.675 ;
        RECT 17.355 168.755 18.565 169.505 ;
        RECT 18.735 168.755 19.945 169.505 ;
        RECT 20.115 168.855 20.375 169.335 ;
        RECT 20.545 168.965 20.795 169.505 ;
        RECT 17.355 168.215 17.875 168.755 ;
        RECT 18.045 168.045 18.565 168.585 ;
        RECT 18.735 168.215 19.255 168.755 ;
        RECT 19.425 168.045 19.945 168.585 ;
        RECT 17.355 166.955 18.565 168.045 ;
        RECT 18.735 166.955 19.945 168.045 ;
        RECT 20.115 167.825 20.285 168.855 ;
        RECT 20.965 168.800 21.185 169.285 ;
        RECT 20.455 168.205 20.685 168.600 ;
        RECT 20.855 168.375 21.185 168.800 ;
        RECT 21.355 169.125 22.245 169.295 ;
        RECT 21.355 168.400 21.525 169.125 ;
        RECT 22.505 168.955 22.675 169.245 ;
        RECT 22.845 169.125 23.175 169.505 ;
        RECT 21.695 168.570 22.245 168.955 ;
        RECT 22.505 168.785 23.170 168.955 ;
        RECT 21.355 168.330 22.245 168.400 ;
        RECT 21.350 168.305 22.245 168.330 ;
        RECT 21.340 168.290 22.245 168.305 ;
        RECT 21.335 168.275 22.245 168.290 ;
        RECT 21.325 168.270 22.245 168.275 ;
        RECT 21.320 168.260 22.245 168.270 ;
        RECT 21.315 168.250 22.245 168.260 ;
        RECT 21.305 168.245 22.245 168.250 ;
        RECT 21.295 168.235 22.245 168.245 ;
        RECT 21.285 168.230 22.245 168.235 ;
        RECT 21.285 168.225 21.620 168.230 ;
        RECT 21.270 168.220 21.620 168.225 ;
        RECT 21.255 168.210 21.620 168.220 ;
        RECT 21.230 168.205 21.620 168.210 ;
        RECT 20.455 168.200 21.620 168.205 ;
        RECT 20.455 168.165 21.590 168.200 ;
        RECT 20.455 168.140 21.555 168.165 ;
        RECT 20.455 168.110 21.525 168.140 ;
        RECT 20.455 168.080 21.505 168.110 ;
        RECT 20.455 168.050 21.485 168.080 ;
        RECT 20.455 168.040 21.415 168.050 ;
        RECT 20.455 168.030 21.390 168.040 ;
        RECT 20.455 168.015 21.370 168.030 ;
        RECT 20.455 168.000 21.350 168.015 ;
        RECT 20.560 167.990 21.345 168.000 ;
        RECT 20.560 167.955 21.330 167.990 ;
        RECT 20.115 167.125 20.390 167.825 ;
        RECT 20.560 167.705 21.315 167.955 ;
        RECT 21.485 167.635 21.815 167.880 ;
        RECT 21.985 167.780 22.245 168.230 ;
        RECT 22.420 167.965 22.770 168.615 ;
        RECT 22.940 167.795 23.170 168.785 ;
        RECT 21.630 167.610 21.815 167.635 ;
        RECT 22.505 167.625 23.170 167.795 ;
        RECT 21.630 167.510 22.245 167.610 ;
        RECT 20.560 166.955 20.815 167.500 ;
        RECT 20.985 167.125 21.465 167.465 ;
        RECT 21.640 166.955 22.245 167.510 ;
        RECT 22.505 167.125 22.675 167.625 ;
        RECT 22.845 166.955 23.175 167.455 ;
        RECT 23.345 167.125 23.530 169.245 ;
        RECT 23.785 169.045 24.035 169.505 ;
        RECT 24.205 169.055 24.540 169.225 ;
        RECT 24.735 169.055 25.410 169.225 ;
        RECT 24.205 168.915 24.375 169.055 ;
        RECT 23.700 167.925 23.980 168.875 ;
        RECT 24.150 168.785 24.375 168.915 ;
        RECT 24.150 167.680 24.320 168.785 ;
        RECT 24.545 168.635 25.070 168.855 ;
        RECT 24.490 167.870 24.730 168.465 ;
        RECT 24.900 167.935 25.070 168.635 ;
        RECT 25.240 168.275 25.410 169.055 ;
        RECT 25.730 169.005 26.100 169.505 ;
        RECT 26.280 169.055 26.685 169.225 ;
        RECT 26.855 169.055 27.640 169.225 ;
        RECT 26.280 168.825 26.450 169.055 ;
        RECT 25.620 168.525 26.450 168.825 ;
        RECT 26.835 168.555 27.300 168.885 ;
        RECT 25.620 168.495 25.820 168.525 ;
        RECT 25.940 168.275 26.110 168.345 ;
        RECT 25.240 168.105 26.110 168.275 ;
        RECT 25.600 168.015 26.110 168.105 ;
        RECT 24.150 167.550 24.455 167.680 ;
        RECT 24.900 167.570 25.430 167.935 ;
        RECT 23.770 166.955 24.035 167.415 ;
        RECT 24.205 167.125 24.455 167.550 ;
        RECT 25.600 167.400 25.770 168.015 ;
        RECT 24.665 167.230 25.770 167.400 ;
        RECT 25.940 166.955 26.110 167.755 ;
        RECT 26.280 167.455 26.450 168.525 ;
        RECT 26.620 167.625 26.810 168.345 ;
        RECT 26.980 167.595 27.300 168.555 ;
        RECT 27.470 168.595 27.640 169.055 ;
        RECT 27.915 168.975 28.125 169.505 ;
        RECT 28.385 168.765 28.715 169.290 ;
        RECT 28.885 168.895 29.055 169.505 ;
        RECT 29.225 168.850 29.555 169.285 ;
        RECT 29.775 169.125 30.665 169.295 ;
        RECT 29.225 168.765 29.605 168.850 ;
        RECT 28.515 168.595 28.715 168.765 ;
        RECT 29.380 168.725 29.605 168.765 ;
        RECT 27.470 168.265 28.345 168.595 ;
        RECT 28.515 168.265 29.265 168.595 ;
        RECT 26.280 167.125 26.530 167.455 ;
        RECT 27.470 167.425 27.640 168.265 ;
        RECT 28.515 168.060 28.705 168.265 ;
        RECT 29.435 168.145 29.605 168.725 ;
        RECT 29.775 168.570 30.325 168.955 ;
        RECT 30.495 168.400 30.665 169.125 ;
        RECT 29.390 168.095 29.605 168.145 ;
        RECT 27.810 167.685 28.705 168.060 ;
        RECT 29.215 168.015 29.605 168.095 ;
        RECT 29.775 168.330 30.665 168.400 ;
        RECT 30.835 168.800 31.055 169.285 ;
        RECT 31.225 168.965 31.475 169.505 ;
        RECT 31.645 168.855 31.905 169.335 ;
        RECT 30.835 168.375 31.165 168.800 ;
        RECT 29.775 168.305 30.670 168.330 ;
        RECT 29.775 168.290 30.680 168.305 ;
        RECT 29.775 168.275 30.685 168.290 ;
        RECT 29.775 168.270 30.695 168.275 ;
        RECT 29.775 168.260 30.700 168.270 ;
        RECT 29.775 168.250 30.705 168.260 ;
        RECT 29.775 168.245 30.715 168.250 ;
        RECT 29.775 168.235 30.725 168.245 ;
        RECT 29.775 168.230 30.735 168.235 ;
        RECT 26.755 167.255 27.640 167.425 ;
        RECT 27.820 166.955 28.135 167.455 ;
        RECT 28.365 167.125 28.705 167.685 ;
        RECT 28.875 166.955 29.045 167.965 ;
        RECT 29.215 167.170 29.545 168.015 ;
        RECT 29.775 167.780 30.035 168.230 ;
        RECT 30.400 168.225 30.735 168.230 ;
        RECT 30.400 168.220 30.750 168.225 ;
        RECT 30.400 168.210 30.765 168.220 ;
        RECT 30.400 168.205 30.790 168.210 ;
        RECT 31.335 168.205 31.565 168.600 ;
        RECT 30.400 168.200 31.565 168.205 ;
        RECT 30.430 168.165 31.565 168.200 ;
        RECT 30.465 168.140 31.565 168.165 ;
        RECT 30.495 168.110 31.565 168.140 ;
        RECT 30.515 168.080 31.565 168.110 ;
        RECT 30.535 168.050 31.565 168.080 ;
        RECT 30.605 168.040 31.565 168.050 ;
        RECT 30.630 168.030 31.565 168.040 ;
        RECT 30.650 168.015 31.565 168.030 ;
        RECT 30.670 168.000 31.565 168.015 ;
        RECT 30.675 167.990 31.460 168.000 ;
        RECT 30.690 167.955 31.460 167.990 ;
        RECT 30.205 167.635 30.535 167.880 ;
        RECT 30.705 167.705 31.460 167.955 ;
        RECT 31.735 167.825 31.905 168.855 ;
        RECT 32.075 168.735 34.665 169.505 ;
        RECT 35.385 168.955 35.555 169.245 ;
        RECT 35.725 169.125 36.055 169.505 ;
        RECT 35.385 168.785 36.050 168.955 ;
        RECT 32.075 168.215 33.285 168.735 ;
        RECT 33.455 168.045 34.665 168.565 ;
        RECT 30.205 167.610 30.390 167.635 ;
        RECT 29.775 167.510 30.390 167.610 ;
        RECT 29.775 166.955 30.380 167.510 ;
        RECT 30.555 167.125 31.035 167.465 ;
        RECT 31.205 166.955 31.460 167.500 ;
        RECT 31.630 167.125 31.905 167.825 ;
        RECT 32.075 166.955 34.665 168.045 ;
        RECT 35.300 167.965 35.650 168.615 ;
        RECT 35.820 167.795 36.050 168.785 ;
        RECT 35.385 167.625 36.050 167.795 ;
        RECT 35.385 167.125 35.555 167.625 ;
        RECT 35.725 166.955 36.055 167.455 ;
        RECT 36.225 167.125 36.410 169.245 ;
        RECT 36.665 169.045 36.915 169.505 ;
        RECT 37.085 169.055 37.420 169.225 ;
        RECT 37.615 169.055 38.290 169.225 ;
        RECT 37.085 168.915 37.255 169.055 ;
        RECT 36.580 167.925 36.860 168.875 ;
        RECT 37.030 168.785 37.255 168.915 ;
        RECT 37.030 167.680 37.200 168.785 ;
        RECT 37.425 168.635 37.950 168.855 ;
        RECT 37.370 167.870 37.610 168.465 ;
        RECT 37.780 167.935 37.950 168.635 ;
        RECT 38.120 168.275 38.290 169.055 ;
        RECT 38.610 169.005 38.980 169.505 ;
        RECT 39.160 169.055 39.565 169.225 ;
        RECT 39.735 169.055 40.520 169.225 ;
        RECT 39.160 168.825 39.330 169.055 ;
        RECT 38.500 168.525 39.330 168.825 ;
        RECT 39.715 168.555 40.180 168.885 ;
        RECT 38.500 168.495 38.700 168.525 ;
        RECT 38.820 168.275 38.990 168.345 ;
        RECT 38.120 168.105 38.990 168.275 ;
        RECT 38.480 168.015 38.990 168.105 ;
        RECT 37.030 167.550 37.335 167.680 ;
        RECT 37.780 167.570 38.310 167.935 ;
        RECT 36.650 166.955 36.915 167.415 ;
        RECT 37.085 167.125 37.335 167.550 ;
        RECT 38.480 167.400 38.650 168.015 ;
        RECT 37.545 167.230 38.650 167.400 ;
        RECT 38.820 166.955 38.990 167.755 ;
        RECT 39.160 167.455 39.330 168.525 ;
        RECT 39.500 167.625 39.690 168.345 ;
        RECT 39.860 167.595 40.180 168.555 ;
        RECT 40.350 168.595 40.520 169.055 ;
        RECT 40.795 168.975 41.005 169.505 ;
        RECT 41.265 168.765 41.595 169.290 ;
        RECT 41.765 168.895 41.935 169.505 ;
        RECT 42.105 168.850 42.435 169.285 ;
        RECT 42.105 168.765 42.485 168.850 ;
        RECT 43.115 168.780 43.405 169.505 ;
        RECT 41.395 168.595 41.595 168.765 ;
        RECT 42.260 168.725 42.485 168.765 ;
        RECT 40.350 168.265 41.225 168.595 ;
        RECT 41.395 168.265 42.145 168.595 ;
        RECT 39.160 167.125 39.410 167.455 ;
        RECT 40.350 167.425 40.520 168.265 ;
        RECT 41.395 168.060 41.585 168.265 ;
        RECT 42.315 168.145 42.485 168.725 ;
        RECT 43.575 168.755 44.785 169.505 ;
        RECT 45.005 168.850 45.335 169.285 ;
        RECT 45.505 168.895 45.675 169.505 ;
        RECT 44.955 168.765 45.335 168.850 ;
        RECT 45.845 168.765 46.175 169.290 ;
        RECT 46.435 168.975 46.645 169.505 ;
        RECT 46.920 169.055 47.705 169.225 ;
        RECT 47.875 169.055 48.280 169.225 ;
        RECT 43.575 168.215 44.095 168.755 ;
        RECT 44.955 168.725 45.180 168.765 ;
        RECT 42.270 168.095 42.485 168.145 ;
        RECT 40.690 167.685 41.585 168.060 ;
        RECT 42.095 168.015 42.485 168.095 ;
        RECT 39.635 167.255 40.520 167.425 ;
        RECT 40.700 166.955 41.015 167.455 ;
        RECT 41.245 167.125 41.585 167.685 ;
        RECT 41.755 166.955 41.925 167.965 ;
        RECT 42.095 167.170 42.425 168.015 ;
        RECT 43.115 166.955 43.405 168.120 ;
        RECT 44.265 168.045 44.785 168.585 ;
        RECT 43.575 166.955 44.785 168.045 ;
        RECT 44.955 168.145 45.125 168.725 ;
        RECT 45.845 168.595 46.045 168.765 ;
        RECT 46.920 168.595 47.090 169.055 ;
        RECT 45.295 168.265 46.045 168.595 ;
        RECT 46.215 168.265 47.090 168.595 ;
        RECT 44.955 168.095 45.170 168.145 ;
        RECT 44.955 168.015 45.345 168.095 ;
        RECT 45.015 167.170 45.345 168.015 ;
        RECT 45.855 168.060 46.045 168.265 ;
        RECT 45.515 166.955 45.685 167.965 ;
        RECT 45.855 167.685 46.750 168.060 ;
        RECT 45.855 167.125 46.195 167.685 ;
        RECT 46.425 166.955 46.740 167.455 ;
        RECT 46.920 167.425 47.090 168.265 ;
        RECT 47.260 168.555 47.725 168.885 ;
        RECT 48.110 168.825 48.280 169.055 ;
        RECT 48.460 169.005 48.830 169.505 ;
        RECT 49.150 169.055 49.825 169.225 ;
        RECT 50.020 169.055 50.355 169.225 ;
        RECT 47.260 167.595 47.580 168.555 ;
        RECT 48.110 168.525 48.940 168.825 ;
        RECT 47.750 167.625 47.940 168.345 ;
        RECT 48.110 167.455 48.280 168.525 ;
        RECT 48.740 168.495 48.940 168.525 ;
        RECT 48.450 168.275 48.620 168.345 ;
        RECT 49.150 168.275 49.320 169.055 ;
        RECT 50.185 168.915 50.355 169.055 ;
        RECT 50.525 169.045 50.775 169.505 ;
        RECT 48.450 168.105 49.320 168.275 ;
        RECT 49.490 168.635 50.015 168.855 ;
        RECT 50.185 168.785 50.410 168.915 ;
        RECT 48.450 168.015 48.960 168.105 ;
        RECT 46.920 167.255 47.805 167.425 ;
        RECT 48.030 167.125 48.280 167.455 ;
        RECT 48.450 166.955 48.620 167.755 ;
        RECT 48.790 167.400 48.960 168.015 ;
        RECT 49.490 167.935 49.660 168.635 ;
        RECT 49.130 167.570 49.660 167.935 ;
        RECT 49.830 167.870 50.070 168.465 ;
        RECT 50.240 167.680 50.410 168.785 ;
        RECT 50.580 167.925 50.860 168.875 ;
        RECT 50.105 167.550 50.410 167.680 ;
        RECT 48.790 167.230 49.895 167.400 ;
        RECT 50.105 167.125 50.355 167.550 ;
        RECT 50.525 166.955 50.790 167.415 ;
        RECT 51.030 167.125 51.215 169.245 ;
        RECT 51.385 169.125 51.715 169.505 ;
        RECT 51.885 168.955 52.055 169.245 ;
        RECT 52.315 168.960 57.660 169.505 ;
        RECT 51.390 168.785 52.055 168.955 ;
        RECT 51.390 167.795 51.620 168.785 ;
        RECT 51.790 167.965 52.140 168.615 ;
        RECT 53.900 168.130 54.240 168.960 ;
        RECT 57.835 168.735 61.345 169.505 ;
        RECT 51.390 167.625 52.055 167.795 ;
        RECT 51.385 166.955 51.715 167.455 ;
        RECT 51.885 167.125 52.055 167.625 ;
        RECT 55.720 167.390 56.070 168.640 ;
        RECT 57.835 168.215 59.485 168.735 ;
        RECT 62.035 168.685 62.245 169.505 ;
        RECT 62.415 168.705 62.745 169.335 ;
        RECT 59.655 168.045 61.345 168.565 ;
        RECT 62.415 168.105 62.665 168.705 ;
        RECT 62.915 168.685 63.145 169.505 ;
        RECT 64.275 168.765 64.660 169.335 ;
        RECT 64.830 169.045 65.155 169.505 ;
        RECT 65.675 168.875 65.955 169.335 ;
        RECT 62.835 168.265 63.165 168.515 ;
        RECT 52.315 166.955 57.660 167.390 ;
        RECT 57.835 166.955 61.345 168.045 ;
        RECT 62.035 166.955 62.245 168.095 ;
        RECT 62.415 167.125 62.745 168.105 ;
        RECT 64.275 168.095 64.555 168.765 ;
        RECT 64.830 168.705 65.955 168.875 ;
        RECT 64.830 168.595 65.280 168.705 ;
        RECT 64.725 168.265 65.280 168.595 ;
        RECT 66.145 168.535 66.545 169.335 ;
        RECT 66.945 169.045 67.215 169.505 ;
        RECT 67.385 168.875 67.670 169.335 ;
        RECT 62.915 166.955 63.145 168.095 ;
        RECT 64.275 167.125 64.660 168.095 ;
        RECT 64.830 167.805 65.280 168.265 ;
        RECT 65.450 167.975 66.545 168.535 ;
        RECT 64.830 167.585 65.955 167.805 ;
        RECT 64.830 166.955 65.155 167.415 ;
        RECT 65.675 167.125 65.955 167.585 ;
        RECT 66.145 167.125 66.545 167.975 ;
        RECT 66.715 168.705 67.670 168.875 ;
        RECT 68.875 168.780 69.165 169.505 ;
        RECT 69.335 168.960 74.680 169.505 ;
        RECT 66.715 167.805 66.925 168.705 ;
        RECT 67.095 167.975 67.785 168.535 ;
        RECT 70.920 168.130 71.260 168.960 ;
        RECT 74.855 168.735 78.365 169.505 ;
        RECT 79.570 168.875 79.855 169.335 ;
        RECT 80.025 169.045 80.295 169.505 ;
        RECT 66.715 167.585 67.670 167.805 ;
        RECT 66.945 166.955 67.215 167.415 ;
        RECT 67.385 167.125 67.670 167.585 ;
        RECT 68.875 166.955 69.165 168.120 ;
        RECT 72.740 167.390 73.090 168.640 ;
        RECT 74.855 168.215 76.505 168.735 ;
        RECT 79.570 168.705 80.525 168.875 ;
        RECT 76.675 168.045 78.365 168.565 ;
        RECT 69.335 166.955 74.680 167.390 ;
        RECT 74.855 166.955 78.365 168.045 ;
        RECT 79.455 167.975 80.145 168.535 ;
        RECT 80.315 167.805 80.525 168.705 ;
        RECT 79.570 167.585 80.525 167.805 ;
        RECT 80.695 168.535 81.095 169.335 ;
        RECT 81.285 168.875 81.565 169.335 ;
        RECT 82.085 169.045 82.410 169.505 ;
        RECT 81.285 168.705 82.410 168.875 ;
        RECT 82.580 168.765 82.965 169.335 ;
        RECT 81.960 168.595 82.410 168.705 ;
        RECT 80.695 167.975 81.790 168.535 ;
        RECT 81.960 168.265 82.515 168.595 ;
        RECT 79.570 167.125 79.855 167.585 ;
        RECT 80.025 166.955 80.295 167.415 ;
        RECT 80.695 167.125 81.095 167.975 ;
        RECT 81.960 167.805 82.410 168.265 ;
        RECT 82.685 168.095 82.965 168.765 ;
        RECT 83.135 168.735 86.645 169.505 ;
        RECT 86.865 168.985 87.120 169.285 ;
        RECT 87.290 169.105 87.620 169.505 ;
        RECT 86.815 168.935 87.120 168.985 ;
        RECT 87.790 168.935 87.960 169.285 ;
        RECT 88.260 169.025 88.430 169.505 ;
        RECT 88.665 168.995 89.015 169.325 ;
        RECT 89.185 169.025 89.355 169.505 ;
        RECT 86.815 168.855 87.960 168.935 ;
        RECT 86.815 168.825 88.525 168.855 ;
        RECT 86.815 168.765 88.675 168.825 ;
        RECT 83.135 168.215 84.785 168.735 ;
        RECT 81.285 167.585 82.410 167.805 ;
        RECT 81.285 167.125 81.565 167.585 ;
        RECT 82.085 166.955 82.410 167.415 ;
        RECT 82.580 167.125 82.965 168.095 ;
        RECT 84.955 168.045 86.645 168.565 ;
        RECT 83.135 166.955 86.645 168.045 ;
        RECT 86.815 168.095 86.985 168.765 ;
        RECT 87.790 168.685 88.675 168.765 ;
        RECT 88.355 168.655 88.675 168.685 ;
        RECT 87.160 168.265 87.460 168.595 ;
        RECT 86.815 167.665 87.120 168.095 ;
        RECT 87.290 167.805 87.460 168.265 ;
        RECT 87.720 167.975 88.255 168.515 ;
        RECT 88.505 168.265 88.675 168.655 ;
        RECT 88.845 168.095 89.015 168.995 ;
        RECT 89.605 168.855 89.865 169.300 ;
        RECT 88.620 167.890 89.015 168.095 ;
        RECT 89.185 168.685 89.865 168.855 ;
        RECT 90.500 168.685 90.775 169.505 ;
        RECT 90.945 168.865 91.275 169.335 ;
        RECT 91.445 169.035 91.615 169.505 ;
        RECT 91.785 168.865 92.115 169.335 ;
        RECT 92.285 169.035 92.455 169.505 ;
        RECT 92.625 168.865 92.955 169.335 ;
        RECT 93.125 169.035 93.295 169.505 ;
        RECT 93.465 168.865 93.795 169.335 ;
        RECT 93.965 169.035 94.250 169.505 ;
        RECT 90.945 168.685 94.465 168.865 ;
        RECT 94.635 168.780 94.925 169.505 ;
        RECT 95.260 168.995 95.500 169.505 ;
        RECT 95.680 168.995 95.960 169.325 ;
        RECT 96.190 168.995 96.405 169.505 ;
        RECT 87.290 167.720 88.400 167.805 ;
        RECT 89.185 167.780 89.355 168.685 ;
        RECT 89.525 167.950 89.865 168.515 ;
        RECT 90.550 168.315 92.210 168.515 ;
        RECT 92.530 168.315 93.895 168.515 ;
        RECT 94.065 168.145 94.465 168.685 ;
        RECT 95.155 168.265 95.510 168.825 ;
        RECT 90.500 167.925 92.535 168.135 ;
        RECT 89.185 167.720 89.865 167.780 ;
        RECT 87.290 167.635 89.865 167.720 ;
        RECT 88.230 167.550 89.865 167.635 ;
        RECT 86.815 167.225 88.015 167.465 ;
        RECT 88.195 166.955 88.525 167.380 ;
        RECT 89.040 166.955 89.400 167.380 ;
        RECT 89.605 167.370 89.865 167.550 ;
        RECT 90.500 167.125 90.775 167.925 ;
        RECT 90.945 166.955 91.275 167.755 ;
        RECT 91.445 167.125 91.615 167.925 ;
        RECT 91.785 166.955 92.035 167.755 ;
        RECT 92.205 167.295 92.535 167.925 ;
        RECT 92.705 167.845 94.465 168.145 ;
        RECT 92.705 167.465 92.875 167.845 ;
        RECT 93.045 167.295 93.375 167.655 ;
        RECT 93.545 167.465 93.715 167.845 ;
        RECT 93.885 167.295 94.300 167.675 ;
        RECT 92.205 167.125 94.300 167.295 ;
        RECT 94.635 166.955 94.925 168.120 ;
        RECT 95.680 168.095 95.850 168.995 ;
        RECT 96.020 168.265 96.285 168.825 ;
        RECT 96.575 168.765 97.190 169.335 ;
        RECT 96.535 168.095 96.705 168.595 ;
        RECT 95.280 167.925 96.705 168.095 ;
        RECT 95.280 167.750 95.670 167.925 ;
        RECT 96.155 166.955 96.485 167.755 ;
        RECT 96.875 167.745 97.190 168.765 ;
        RECT 97.855 168.885 98.120 169.335 ;
        RECT 98.290 169.055 98.580 169.505 ;
        RECT 98.750 168.885 99.040 169.335 ;
        RECT 97.855 168.715 99.040 168.885 ;
        RECT 99.220 168.595 99.465 169.200 ;
        RECT 97.875 167.930 98.205 168.515 ;
        RECT 98.375 168.265 98.860 168.515 ;
        RECT 99.205 168.265 99.465 168.595 ;
        RECT 99.715 168.265 99.985 169.200 ;
        RECT 100.165 168.515 100.375 169.200 ;
        RECT 100.545 168.855 100.885 169.335 ;
        RECT 101.065 169.025 101.375 169.505 ;
        RECT 100.545 168.685 101.215 168.855 ;
        RECT 101.045 168.595 101.215 168.685 ;
        RECT 100.165 168.265 100.645 168.515 ;
        RECT 101.045 168.265 101.385 168.595 ;
        RECT 96.655 167.125 97.190 167.745 ;
        RECT 97.855 166.955 98.180 167.755 ;
        RECT 98.375 167.175 98.560 168.265 ;
        RECT 101.045 168.095 101.215 168.265 ;
        RECT 98.730 167.925 101.215 168.095 ;
        RECT 98.730 167.125 98.980 167.925 ;
        RECT 99.150 166.955 99.890 167.755 ;
        RECT 100.075 167.125 100.405 167.925 ;
        RECT 100.575 166.955 101.385 167.755 ;
        RECT 101.555 167.125 101.815 169.335 ;
        RECT 101.995 168.765 102.380 169.335 ;
        RECT 102.550 169.045 102.875 169.505 ;
        RECT 103.395 168.875 103.675 169.335 ;
        RECT 101.995 168.095 102.275 168.765 ;
        RECT 102.550 168.705 103.675 168.875 ;
        RECT 102.550 168.595 103.000 168.705 ;
        RECT 102.445 168.265 103.000 168.595 ;
        RECT 103.865 168.535 104.265 169.335 ;
        RECT 104.665 169.045 104.935 169.505 ;
        RECT 105.105 168.875 105.390 169.335 ;
        RECT 101.995 167.125 102.380 168.095 ;
        RECT 102.550 167.805 103.000 168.265 ;
        RECT 103.170 167.975 104.265 168.535 ;
        RECT 102.550 167.585 103.675 167.805 ;
        RECT 102.550 166.955 102.875 167.415 ;
        RECT 103.395 167.125 103.675 167.585 ;
        RECT 103.865 167.125 104.265 167.975 ;
        RECT 104.435 168.705 105.390 168.875 ;
        RECT 105.675 169.005 105.935 169.335 ;
        RECT 106.105 169.145 106.435 169.505 ;
        RECT 106.690 169.125 107.990 169.335 ;
        RECT 105.675 168.995 105.905 169.005 ;
        RECT 104.435 167.805 104.645 168.705 ;
        RECT 104.815 167.975 105.505 168.535 ;
        RECT 105.675 167.805 105.845 168.995 ;
        RECT 106.690 168.975 106.860 169.125 ;
        RECT 106.105 168.850 106.860 168.975 ;
        RECT 106.015 168.805 106.860 168.850 ;
        RECT 106.015 168.685 106.285 168.805 ;
        RECT 106.015 168.110 106.185 168.685 ;
        RECT 106.415 168.245 106.825 168.550 ;
        RECT 107.115 168.515 107.325 168.915 ;
        RECT 106.995 168.305 107.325 168.515 ;
        RECT 107.570 168.515 107.790 168.915 ;
        RECT 108.265 168.740 108.720 169.505 ;
        RECT 110.085 168.705 110.345 169.505 ;
        RECT 110.515 168.855 110.845 169.335 ;
        RECT 111.015 169.025 111.205 169.505 ;
        RECT 111.375 169.085 113.425 169.335 ;
        RECT 111.375 168.855 111.635 169.085 ;
        RECT 113.595 169.065 113.875 169.505 ;
        RECT 114.065 168.975 114.255 169.335 ;
        RECT 114.425 169.145 114.755 169.505 ;
        RECT 114.925 168.975 115.115 169.220 ;
        RECT 110.515 168.685 111.635 168.855 ;
        RECT 111.805 168.895 113.435 168.915 ;
        RECT 114.065 168.895 115.115 168.975 ;
        RECT 111.805 168.725 115.115 168.895 ;
        RECT 115.285 168.785 115.620 169.505 ;
        RECT 111.805 168.695 114.110 168.725 ;
        RECT 107.570 168.305 108.045 168.515 ;
        RECT 108.235 168.315 108.725 168.515 ;
        RECT 106.015 168.075 106.215 168.110 ;
        RECT 107.545 168.075 108.720 168.135 ;
        RECT 106.015 167.965 108.720 168.075 ;
        RECT 106.075 167.905 107.875 167.965 ;
        RECT 107.545 167.875 107.875 167.905 ;
        RECT 104.435 167.585 105.390 167.805 ;
        RECT 104.665 166.955 104.935 167.415 ;
        RECT 105.105 167.125 105.390 167.585 ;
        RECT 105.675 167.125 105.935 167.805 ;
        RECT 106.105 166.955 106.355 167.735 ;
        RECT 106.605 167.705 107.440 167.715 ;
        RECT 108.030 167.705 108.215 167.795 ;
        RECT 106.605 167.505 108.215 167.705 ;
        RECT 106.605 167.125 106.855 167.505 ;
        RECT 107.985 167.465 108.215 167.505 ;
        RECT 108.465 167.345 108.720 167.965 ;
        RECT 110.240 168.110 111.485 168.515 ;
        RECT 111.710 168.280 113.145 168.525 ;
        RECT 113.315 168.110 113.660 168.525 ;
        RECT 110.240 167.885 113.660 168.110 ;
        RECT 113.830 168.005 114.110 168.695 ;
        RECT 115.835 168.685 116.065 169.505 ;
        RECT 116.235 168.705 116.565 169.335 ;
        RECT 115.310 168.555 115.620 168.595 ;
        RECT 114.280 168.175 115.620 168.555 ;
        RECT 115.815 168.265 116.145 168.515 ;
        RECT 116.315 168.105 116.565 168.705 ;
        RECT 116.735 168.685 116.945 169.505 ;
        RECT 117.175 168.705 117.870 169.335 ;
        RECT 118.075 168.705 118.385 169.505 ;
        RECT 119.015 168.705 119.325 169.505 ;
        RECT 119.530 168.705 120.225 169.335 ;
        RECT 120.395 168.780 120.685 169.505 ;
        RECT 120.870 168.935 121.125 169.285 ;
        RECT 121.295 169.105 121.625 169.505 ;
        RECT 121.795 168.935 121.965 169.285 ;
        RECT 122.135 169.105 122.515 169.505 ;
        RECT 120.870 168.765 122.535 168.935 ;
        RECT 122.705 168.830 122.980 169.175 ;
        RECT 123.215 169.045 123.460 169.505 ;
        RECT 117.195 168.265 117.530 168.515 ;
        RECT 117.700 168.105 117.870 168.705 ;
        RECT 118.040 168.265 118.375 168.535 ;
        RECT 119.025 168.265 119.360 168.535 ;
        RECT 119.530 168.105 119.700 168.705 ;
        RECT 122.365 168.595 122.535 168.765 ;
        RECT 119.870 168.265 120.205 168.515 ;
        RECT 120.855 168.265 121.200 168.595 ;
        RECT 121.370 168.265 122.195 168.595 ;
        RECT 122.365 168.265 122.640 168.595 ;
        RECT 113.830 167.885 115.130 168.005 ;
        RECT 107.025 166.955 107.380 167.335 ;
        RECT 108.385 167.125 108.720 167.345 ;
        RECT 110.085 167.485 113.795 167.715 ;
        RECT 113.965 167.555 115.130 167.885 ;
        RECT 110.085 167.125 110.345 167.485 ;
        RECT 110.515 166.955 110.845 167.315 ;
        RECT 111.025 167.125 111.205 167.485 ;
        RECT 111.375 166.955 111.705 167.315 ;
        RECT 111.875 167.125 112.065 167.485 ;
        RECT 112.235 166.955 112.565 167.315 ;
        RECT 112.735 167.125 112.925 167.485 ;
        RECT 113.595 167.385 113.795 167.485 ;
        RECT 113.595 167.375 114.755 167.385 ;
        RECT 115.335 167.375 115.530 167.795 ;
        RECT 113.095 166.955 113.425 167.315 ;
        RECT 113.595 167.125 115.530 167.375 ;
        RECT 115.835 166.955 116.065 168.095 ;
        RECT 116.235 167.125 116.565 168.105 ;
        RECT 116.735 166.955 116.945 168.095 ;
        RECT 117.175 166.955 117.435 168.095 ;
        RECT 117.605 167.125 117.935 168.105 ;
        RECT 118.105 166.955 118.385 168.095 ;
        RECT 119.015 166.955 119.295 168.095 ;
        RECT 119.465 167.125 119.795 168.105 ;
        RECT 119.965 166.955 120.225 168.095 ;
        RECT 120.395 166.955 120.685 168.120 ;
        RECT 120.875 167.805 121.200 168.095 ;
        RECT 121.370 167.975 121.565 168.265 ;
        RECT 122.365 168.095 122.535 168.265 ;
        RECT 122.810 168.095 122.980 168.830 ;
        RECT 123.155 168.265 123.470 168.875 ;
        RECT 123.640 168.515 123.890 169.325 ;
        RECT 124.060 168.980 124.320 169.505 ;
        RECT 124.490 168.855 124.750 169.310 ;
        RECT 124.920 169.025 125.180 169.505 ;
        RECT 125.350 168.855 125.610 169.310 ;
        RECT 125.780 169.025 126.040 169.505 ;
        RECT 126.210 168.855 126.470 169.310 ;
        RECT 126.640 169.025 126.900 169.505 ;
        RECT 127.070 168.855 127.330 169.310 ;
        RECT 127.500 169.025 127.800 169.505 ;
        RECT 124.490 168.685 127.800 168.855 ;
        RECT 128.420 168.725 128.920 169.335 ;
        RECT 123.640 168.265 126.660 168.515 ;
        RECT 121.875 167.925 122.535 168.095 ;
        RECT 121.875 167.805 122.045 167.925 ;
        RECT 120.875 167.635 122.045 167.805 ;
        RECT 120.855 167.175 122.045 167.465 ;
        RECT 122.215 166.955 122.495 167.755 ;
        RECT 122.705 167.125 122.980 168.095 ;
        RECT 123.165 166.955 123.460 168.065 ;
        RECT 123.640 167.130 123.890 168.265 ;
        RECT 126.830 168.095 127.800 168.685 ;
        RECT 128.215 168.265 128.565 168.515 ;
        RECT 128.750 168.095 128.920 168.725 ;
        RECT 129.550 168.855 129.880 169.335 ;
        RECT 130.050 169.045 130.275 169.505 ;
        RECT 130.445 168.855 130.775 169.335 ;
        RECT 129.550 168.685 130.775 168.855 ;
        RECT 130.965 168.705 131.215 169.505 ;
        RECT 131.385 168.705 131.725 169.335 ;
        RECT 131.900 168.740 132.355 169.505 ;
        RECT 132.630 169.125 133.930 169.335 ;
        RECT 134.185 169.145 134.515 169.505 ;
        RECT 133.760 168.975 133.930 169.125 ;
        RECT 134.685 169.005 134.945 169.335 ;
        RECT 134.715 168.995 134.945 169.005 ;
        RECT 131.495 168.655 131.725 168.705 ;
        RECT 129.090 168.315 129.420 168.515 ;
        RECT 129.590 168.315 129.920 168.515 ;
        RECT 130.090 168.315 130.510 168.515 ;
        RECT 130.685 168.345 131.380 168.515 ;
        RECT 130.685 168.095 130.855 168.345 ;
        RECT 131.550 168.095 131.725 168.655 ;
        RECT 132.830 168.515 133.050 168.915 ;
        RECT 131.895 168.315 132.385 168.515 ;
        RECT 132.575 168.305 133.050 168.515 ;
        RECT 133.295 168.515 133.505 168.915 ;
        RECT 133.760 168.850 134.515 168.975 ;
        RECT 133.760 168.805 134.605 168.850 ;
        RECT 134.335 168.685 134.605 168.805 ;
        RECT 133.295 168.305 133.625 168.515 ;
        RECT 133.795 168.245 134.205 168.550 ;
        RECT 124.060 166.955 124.320 168.065 ;
        RECT 124.490 167.855 127.800 168.095 ;
        RECT 128.420 167.925 130.855 168.095 ;
        RECT 124.490 167.130 124.750 167.855 ;
        RECT 124.920 166.955 125.180 167.685 ;
        RECT 125.350 167.130 125.610 167.855 ;
        RECT 125.780 166.955 126.040 167.685 ;
        RECT 126.210 167.130 126.470 167.855 ;
        RECT 126.640 166.955 126.900 167.685 ;
        RECT 127.070 167.130 127.330 167.855 ;
        RECT 127.500 166.955 127.795 167.685 ;
        RECT 128.420 167.125 128.750 167.925 ;
        RECT 128.920 166.955 129.250 167.755 ;
        RECT 129.550 167.125 129.880 167.925 ;
        RECT 130.525 166.955 130.775 167.755 ;
        RECT 131.045 166.955 131.215 168.095 ;
        RECT 131.385 167.125 131.725 168.095 ;
        RECT 131.900 168.075 133.075 168.135 ;
        RECT 134.435 168.110 134.605 168.685 ;
        RECT 134.405 168.075 134.605 168.110 ;
        RECT 131.900 167.965 134.605 168.075 ;
        RECT 131.900 167.345 132.155 167.965 ;
        RECT 132.745 167.905 134.545 167.965 ;
        RECT 132.745 167.875 133.075 167.905 ;
        RECT 134.775 167.805 134.945 168.995 ;
        RECT 135.665 168.955 135.835 169.245 ;
        RECT 136.005 169.125 136.335 169.505 ;
        RECT 135.665 168.785 136.330 168.955 ;
        RECT 135.580 167.965 135.930 168.615 ;
        RECT 132.405 167.705 132.590 167.795 ;
        RECT 133.180 167.705 134.015 167.715 ;
        RECT 132.405 167.505 134.015 167.705 ;
        RECT 132.405 167.465 132.635 167.505 ;
        RECT 131.900 167.125 132.235 167.345 ;
        RECT 133.240 166.955 133.595 167.335 ;
        RECT 133.765 167.125 134.015 167.505 ;
        RECT 134.265 166.955 134.515 167.735 ;
        RECT 134.685 167.125 134.945 167.805 ;
        RECT 136.100 167.795 136.330 168.785 ;
        RECT 135.665 167.625 136.330 167.795 ;
        RECT 135.665 167.125 135.835 167.625 ;
        RECT 136.005 166.955 136.335 167.455 ;
        RECT 136.505 167.125 136.690 169.245 ;
        RECT 136.945 169.045 137.195 169.505 ;
        RECT 137.365 169.055 137.700 169.225 ;
        RECT 137.895 169.055 138.570 169.225 ;
        RECT 137.365 168.915 137.535 169.055 ;
        RECT 136.860 167.925 137.140 168.875 ;
        RECT 137.310 168.785 137.535 168.915 ;
        RECT 137.310 167.680 137.480 168.785 ;
        RECT 137.705 168.635 138.230 168.855 ;
        RECT 137.650 167.870 137.890 168.465 ;
        RECT 138.060 167.935 138.230 168.635 ;
        RECT 138.400 168.275 138.570 169.055 ;
        RECT 138.890 169.005 139.260 169.505 ;
        RECT 139.440 169.055 139.845 169.225 ;
        RECT 140.015 169.055 140.800 169.225 ;
        RECT 139.440 168.825 139.610 169.055 ;
        RECT 138.780 168.525 139.610 168.825 ;
        RECT 139.995 168.555 140.460 168.885 ;
        RECT 138.780 168.495 138.980 168.525 ;
        RECT 139.100 168.275 139.270 168.345 ;
        RECT 138.400 168.105 139.270 168.275 ;
        RECT 138.760 168.015 139.270 168.105 ;
        RECT 137.310 167.550 137.615 167.680 ;
        RECT 138.060 167.570 138.590 167.935 ;
        RECT 136.930 166.955 137.195 167.415 ;
        RECT 137.365 167.125 137.615 167.550 ;
        RECT 138.760 167.400 138.930 168.015 ;
        RECT 137.825 167.230 138.930 167.400 ;
        RECT 139.100 166.955 139.270 167.755 ;
        RECT 139.440 167.455 139.610 168.525 ;
        RECT 139.780 167.625 139.970 168.345 ;
        RECT 140.140 167.595 140.460 168.555 ;
        RECT 140.630 168.595 140.800 169.055 ;
        RECT 141.075 168.975 141.285 169.505 ;
        RECT 141.545 168.765 141.875 169.290 ;
        RECT 142.045 168.895 142.215 169.505 ;
        RECT 142.385 168.850 142.715 169.285 ;
        RECT 143.945 168.955 144.115 169.335 ;
        RECT 144.330 169.125 144.660 169.505 ;
        RECT 142.385 168.765 142.765 168.850 ;
        RECT 143.945 168.785 144.660 168.955 ;
        RECT 141.675 168.595 141.875 168.765 ;
        RECT 142.540 168.725 142.765 168.765 ;
        RECT 140.630 168.265 141.505 168.595 ;
        RECT 141.675 168.265 142.425 168.595 ;
        RECT 139.440 167.125 139.690 167.455 ;
        RECT 140.630 167.425 140.800 168.265 ;
        RECT 141.675 168.060 141.865 168.265 ;
        RECT 142.595 168.145 142.765 168.725 ;
        RECT 143.855 168.235 144.210 168.605 ;
        RECT 144.490 168.595 144.660 168.785 ;
        RECT 144.830 168.760 145.085 169.335 ;
        RECT 144.490 168.265 144.745 168.595 ;
        RECT 142.550 168.095 142.765 168.145 ;
        RECT 140.970 167.685 141.865 168.060 ;
        RECT 142.375 168.015 142.765 168.095 ;
        RECT 144.490 168.055 144.660 168.265 ;
        RECT 139.915 167.255 140.800 167.425 ;
        RECT 140.980 166.955 141.295 167.455 ;
        RECT 141.525 167.125 141.865 167.685 ;
        RECT 142.035 166.955 142.205 167.965 ;
        RECT 142.375 167.170 142.705 168.015 ;
        RECT 143.945 167.885 144.660 168.055 ;
        RECT 144.915 168.030 145.085 168.760 ;
        RECT 145.260 168.665 145.520 169.505 ;
        RECT 145.695 168.755 146.905 169.505 ;
        RECT 143.945 167.125 144.115 167.885 ;
        RECT 144.330 166.955 144.660 167.715 ;
        RECT 144.830 167.125 145.085 168.030 ;
        RECT 145.260 166.955 145.520 168.105 ;
        RECT 145.695 168.045 146.215 168.585 ;
        RECT 146.385 168.215 146.905 168.755 ;
        RECT 145.695 166.955 146.905 168.045 ;
        RECT 17.270 166.785 146.990 166.955 ;
        RECT 17.355 165.695 18.565 166.785 ;
        RECT 18.735 166.350 24.080 166.785 ;
        RECT 24.255 166.350 29.600 166.785 ;
        RECT 17.355 164.985 17.875 165.525 ;
        RECT 18.045 165.155 18.565 165.695 ;
        RECT 17.355 164.235 18.565 164.985 ;
        RECT 20.320 164.780 20.660 165.610 ;
        RECT 22.140 165.100 22.490 166.350 ;
        RECT 25.840 164.780 26.180 165.610 ;
        RECT 27.660 165.100 28.010 166.350 ;
        RECT 30.235 165.620 30.525 166.785 ;
        RECT 30.695 166.350 36.040 166.785 ;
        RECT 18.735 164.235 24.080 164.780 ;
        RECT 24.255 164.235 29.600 164.780 ;
        RECT 30.235 164.235 30.525 164.960 ;
        RECT 32.280 164.780 32.620 165.610 ;
        RECT 34.100 165.100 34.450 166.350 ;
        RECT 36.675 165.915 36.950 166.615 ;
        RECT 37.120 166.240 37.375 166.785 ;
        RECT 37.545 166.275 38.025 166.615 ;
        RECT 38.200 166.230 38.805 166.785 ;
        RECT 38.975 166.350 44.320 166.785 ;
        RECT 44.495 166.350 49.840 166.785 ;
        RECT 50.015 166.350 55.360 166.785 ;
        RECT 38.190 166.130 38.805 166.230 ;
        RECT 38.190 166.105 38.375 166.130 ;
        RECT 36.675 164.885 36.845 165.915 ;
        RECT 37.120 165.785 37.875 166.035 ;
        RECT 38.045 165.860 38.375 166.105 ;
        RECT 37.120 165.750 37.890 165.785 ;
        RECT 37.120 165.740 37.905 165.750 ;
        RECT 37.015 165.725 37.910 165.740 ;
        RECT 37.015 165.710 37.930 165.725 ;
        RECT 37.015 165.700 37.950 165.710 ;
        RECT 37.015 165.690 37.975 165.700 ;
        RECT 37.015 165.660 38.045 165.690 ;
        RECT 37.015 165.630 38.065 165.660 ;
        RECT 37.015 165.600 38.085 165.630 ;
        RECT 37.015 165.575 38.115 165.600 ;
        RECT 37.015 165.540 38.150 165.575 ;
        RECT 37.015 165.535 38.180 165.540 ;
        RECT 37.015 165.140 37.245 165.535 ;
        RECT 37.790 165.530 38.180 165.535 ;
        RECT 37.815 165.520 38.180 165.530 ;
        RECT 37.830 165.515 38.180 165.520 ;
        RECT 37.845 165.510 38.180 165.515 ;
        RECT 38.545 165.510 38.805 165.960 ;
        RECT 37.845 165.505 38.805 165.510 ;
        RECT 37.855 165.495 38.805 165.505 ;
        RECT 37.865 165.490 38.805 165.495 ;
        RECT 37.875 165.480 38.805 165.490 ;
        RECT 37.880 165.470 38.805 165.480 ;
        RECT 37.885 165.465 38.805 165.470 ;
        RECT 37.895 165.450 38.805 165.465 ;
        RECT 37.900 165.435 38.805 165.450 ;
        RECT 37.910 165.410 38.805 165.435 ;
        RECT 37.415 164.940 37.745 165.365 ;
        RECT 30.695 164.235 36.040 164.780 ;
        RECT 36.675 164.405 36.935 164.885 ;
        RECT 37.105 164.235 37.355 164.775 ;
        RECT 37.525 164.455 37.745 164.940 ;
        RECT 37.915 165.340 38.805 165.410 ;
        RECT 37.915 164.615 38.085 165.340 ;
        RECT 38.255 164.785 38.805 165.170 ;
        RECT 40.560 164.780 40.900 165.610 ;
        RECT 42.380 165.100 42.730 166.350 ;
        RECT 46.080 164.780 46.420 165.610 ;
        RECT 47.900 165.100 48.250 166.350 ;
        RECT 51.600 164.780 51.940 165.610 ;
        RECT 53.420 165.100 53.770 166.350 ;
        RECT 55.995 165.620 56.285 166.785 ;
        RECT 56.455 165.695 58.125 166.785 ;
        RECT 58.870 166.155 59.155 166.615 ;
        RECT 59.325 166.325 59.595 166.785 ;
        RECT 58.870 165.935 59.825 166.155 ;
        RECT 56.455 165.005 57.205 165.525 ;
        RECT 57.375 165.175 58.125 165.695 ;
        RECT 58.755 165.205 59.445 165.765 ;
        RECT 59.615 165.035 59.825 165.935 ;
        RECT 37.915 164.445 38.805 164.615 ;
        RECT 38.975 164.235 44.320 164.780 ;
        RECT 44.495 164.235 49.840 164.780 ;
        RECT 50.015 164.235 55.360 164.780 ;
        RECT 55.995 164.235 56.285 164.960 ;
        RECT 56.455 164.235 58.125 165.005 ;
        RECT 58.870 164.865 59.825 165.035 ;
        RECT 59.995 165.765 60.395 166.615 ;
        RECT 60.585 166.155 60.865 166.615 ;
        RECT 61.385 166.325 61.710 166.785 ;
        RECT 60.585 165.935 61.710 166.155 ;
        RECT 59.995 165.205 61.090 165.765 ;
        RECT 61.260 165.475 61.710 165.935 ;
        RECT 61.880 165.645 62.265 166.615 ;
        RECT 58.870 164.405 59.155 164.865 ;
        RECT 59.325 164.235 59.595 164.695 ;
        RECT 59.995 164.405 60.395 165.205 ;
        RECT 61.260 165.145 61.815 165.475 ;
        RECT 61.260 165.035 61.710 165.145 ;
        RECT 60.585 164.865 61.710 165.035 ;
        RECT 61.985 164.975 62.265 165.645 ;
        RECT 60.585 164.405 60.865 164.865 ;
        RECT 61.385 164.235 61.710 164.695 ;
        RECT 61.880 164.405 62.265 164.975 ;
        RECT 62.445 164.415 62.705 166.605 ;
        RECT 62.875 166.055 63.215 166.785 ;
        RECT 63.395 165.875 63.665 166.605 ;
        RECT 62.895 165.655 63.665 165.875 ;
        RECT 63.845 165.895 64.075 166.605 ;
        RECT 64.245 166.075 64.575 166.785 ;
        RECT 64.745 165.895 65.005 166.605 ;
        RECT 63.845 165.655 65.005 165.895 ;
        RECT 66.150 165.995 66.685 166.615 ;
        RECT 62.895 164.985 63.185 165.655 ;
        RECT 63.365 165.165 63.830 165.475 ;
        RECT 64.010 165.165 64.535 165.475 ;
        RECT 62.895 164.785 64.125 164.985 ;
        RECT 62.965 164.235 63.635 164.605 ;
        RECT 63.815 164.415 64.125 164.785 ;
        RECT 64.305 164.525 64.535 165.165 ;
        RECT 64.715 165.145 65.015 165.475 ;
        RECT 66.150 164.975 66.465 165.995 ;
        RECT 66.855 165.985 67.185 166.785 ;
        RECT 68.420 166.360 68.755 166.785 ;
        RECT 68.925 166.180 69.110 166.585 ;
        RECT 68.445 166.005 69.110 166.180 ;
        RECT 69.315 166.005 69.645 166.785 ;
        RECT 67.670 165.815 68.060 165.990 ;
        RECT 66.635 165.645 68.060 165.815 ;
        RECT 66.635 165.145 66.805 165.645 ;
        RECT 64.715 164.235 65.005 164.965 ;
        RECT 66.150 164.405 66.765 164.975 ;
        RECT 67.055 164.915 67.320 165.475 ;
        RECT 67.490 164.745 67.660 165.645 ;
        RECT 67.830 164.915 68.185 165.475 ;
        RECT 68.445 164.975 68.785 166.005 ;
        RECT 69.815 165.815 70.085 166.585 ;
        RECT 68.955 165.645 70.085 165.815 ;
        RECT 70.265 165.815 70.595 166.600 ;
        RECT 70.265 165.645 70.945 165.815 ;
        RECT 71.125 165.645 71.455 166.785 ;
        RECT 71.725 166.115 71.895 166.615 ;
        RECT 72.065 166.285 72.395 166.785 ;
        RECT 71.725 165.945 72.390 166.115 ;
        RECT 68.955 165.145 69.205 165.645 ;
        RECT 68.445 164.805 69.130 164.975 ;
        RECT 69.385 164.895 69.745 165.475 ;
        RECT 66.935 164.235 67.150 164.745 ;
        RECT 67.380 164.415 67.660 164.745 ;
        RECT 67.840 164.235 68.080 164.745 ;
        RECT 68.420 164.235 68.755 164.635 ;
        RECT 68.925 164.405 69.130 164.805 ;
        RECT 69.915 164.735 70.085 165.645 ;
        RECT 70.255 165.225 70.605 165.475 ;
        RECT 70.775 165.045 70.945 165.645 ;
        RECT 71.115 165.225 71.465 165.475 ;
        RECT 71.640 165.125 71.990 165.775 ;
        RECT 69.340 164.235 69.615 164.715 ;
        RECT 69.825 164.405 70.085 164.735 ;
        RECT 70.275 164.235 70.515 165.045 ;
        RECT 70.685 164.405 71.015 165.045 ;
        RECT 71.185 164.235 71.455 165.045 ;
        RECT 72.160 164.955 72.390 165.945 ;
        RECT 71.725 164.785 72.390 164.955 ;
        RECT 71.725 164.495 71.895 164.785 ;
        RECT 72.065 164.235 72.395 164.615 ;
        RECT 72.565 164.495 72.750 166.615 ;
        RECT 72.990 166.325 73.255 166.785 ;
        RECT 73.425 166.190 73.675 166.615 ;
        RECT 73.885 166.340 74.990 166.510 ;
        RECT 73.370 166.060 73.675 166.190 ;
        RECT 72.920 164.865 73.200 165.815 ;
        RECT 73.370 164.955 73.540 166.060 ;
        RECT 73.710 165.275 73.950 165.870 ;
        RECT 74.120 165.805 74.650 166.170 ;
        RECT 74.120 165.105 74.290 165.805 ;
        RECT 74.820 165.725 74.990 166.340 ;
        RECT 75.160 165.985 75.330 166.785 ;
        RECT 75.500 166.285 75.750 166.615 ;
        RECT 75.975 166.315 76.860 166.485 ;
        RECT 74.820 165.635 75.330 165.725 ;
        RECT 73.370 164.825 73.595 164.955 ;
        RECT 73.765 164.885 74.290 165.105 ;
        RECT 74.460 165.465 75.330 165.635 ;
        RECT 73.005 164.235 73.255 164.695 ;
        RECT 73.425 164.685 73.595 164.825 ;
        RECT 74.460 164.685 74.630 165.465 ;
        RECT 75.160 165.395 75.330 165.465 ;
        RECT 74.840 165.215 75.040 165.245 ;
        RECT 75.500 165.215 75.670 166.285 ;
        RECT 75.840 165.395 76.030 166.115 ;
        RECT 74.840 164.915 75.670 165.215 ;
        RECT 76.200 165.185 76.520 166.145 ;
        RECT 73.425 164.515 73.760 164.685 ;
        RECT 73.955 164.515 74.630 164.685 ;
        RECT 74.950 164.235 75.320 164.735 ;
        RECT 75.500 164.685 75.670 164.915 ;
        RECT 76.055 164.855 76.520 165.185 ;
        RECT 76.690 165.475 76.860 166.315 ;
        RECT 77.040 166.285 77.355 166.785 ;
        RECT 77.585 166.055 77.925 166.615 ;
        RECT 77.030 165.680 77.925 166.055 ;
        RECT 78.095 165.775 78.265 166.785 ;
        RECT 77.735 165.475 77.925 165.680 ;
        RECT 78.435 165.725 78.765 166.570 ;
        RECT 78.995 165.915 79.270 166.615 ;
        RECT 79.440 166.240 79.695 166.785 ;
        RECT 79.865 166.275 80.345 166.615 ;
        RECT 80.520 166.230 81.125 166.785 ;
        RECT 80.510 166.130 81.125 166.230 ;
        RECT 80.510 166.105 80.695 166.130 ;
        RECT 78.435 165.645 78.825 165.725 ;
        RECT 78.610 165.595 78.825 165.645 ;
        RECT 76.690 165.145 77.565 165.475 ;
        RECT 77.735 165.145 78.485 165.475 ;
        RECT 76.690 164.685 76.860 165.145 ;
        RECT 77.735 164.975 77.935 165.145 ;
        RECT 78.655 165.015 78.825 165.595 ;
        RECT 78.600 164.975 78.825 165.015 ;
        RECT 75.500 164.515 75.905 164.685 ;
        RECT 76.075 164.515 76.860 164.685 ;
        RECT 77.135 164.235 77.345 164.765 ;
        RECT 77.605 164.450 77.935 164.975 ;
        RECT 78.445 164.890 78.825 164.975 ;
        RECT 78.105 164.235 78.275 164.845 ;
        RECT 78.445 164.455 78.775 164.890 ;
        RECT 78.995 164.885 79.165 165.915 ;
        RECT 79.440 165.785 80.195 166.035 ;
        RECT 80.365 165.860 80.695 166.105 ;
        RECT 79.440 165.750 80.210 165.785 ;
        RECT 79.440 165.740 80.225 165.750 ;
        RECT 79.335 165.725 80.230 165.740 ;
        RECT 79.335 165.710 80.250 165.725 ;
        RECT 79.335 165.700 80.270 165.710 ;
        RECT 79.335 165.690 80.295 165.700 ;
        RECT 79.335 165.660 80.365 165.690 ;
        RECT 79.335 165.630 80.385 165.660 ;
        RECT 79.335 165.600 80.405 165.630 ;
        RECT 79.335 165.575 80.435 165.600 ;
        RECT 79.335 165.540 80.470 165.575 ;
        RECT 79.335 165.535 80.500 165.540 ;
        RECT 79.335 165.140 79.565 165.535 ;
        RECT 80.110 165.530 80.500 165.535 ;
        RECT 80.135 165.520 80.500 165.530 ;
        RECT 80.150 165.515 80.500 165.520 ;
        RECT 80.165 165.510 80.500 165.515 ;
        RECT 80.865 165.510 81.125 165.960 ;
        RECT 81.755 165.620 82.045 166.785 ;
        RECT 82.215 166.350 87.560 166.785 ;
        RECT 87.735 166.350 93.080 166.785 ;
        RECT 80.165 165.505 81.125 165.510 ;
        RECT 80.175 165.495 81.125 165.505 ;
        RECT 80.185 165.490 81.125 165.495 ;
        RECT 80.195 165.480 81.125 165.490 ;
        RECT 80.200 165.470 81.125 165.480 ;
        RECT 80.205 165.465 81.125 165.470 ;
        RECT 80.215 165.450 81.125 165.465 ;
        RECT 80.220 165.435 81.125 165.450 ;
        RECT 80.230 165.410 81.125 165.435 ;
        RECT 79.735 164.940 80.065 165.365 ;
        RECT 79.815 164.915 80.065 164.940 ;
        RECT 78.995 164.405 79.255 164.885 ;
        RECT 79.425 164.235 79.675 164.775 ;
        RECT 79.845 164.455 80.065 164.915 ;
        RECT 80.235 165.340 81.125 165.410 ;
        RECT 80.235 164.615 80.405 165.340 ;
        RECT 80.575 164.785 81.125 165.170 ;
        RECT 80.235 164.445 81.125 164.615 ;
        RECT 81.755 164.235 82.045 164.960 ;
        RECT 83.800 164.780 84.140 165.610 ;
        RECT 85.620 165.100 85.970 166.350 ;
        RECT 89.320 164.780 89.660 165.610 ;
        RECT 91.140 165.100 91.490 166.350 ;
        RECT 93.255 165.695 96.765 166.785 ;
        RECT 93.255 165.005 94.905 165.525 ;
        RECT 95.075 165.175 96.765 165.695 ;
        RECT 97.405 165.815 97.735 166.600 ;
        RECT 97.405 165.645 98.085 165.815 ;
        RECT 98.265 165.645 98.595 166.785 ;
        RECT 98.775 166.350 104.120 166.785 ;
        RECT 97.395 165.225 97.745 165.475 ;
        RECT 97.915 165.045 98.085 165.645 ;
        RECT 98.255 165.225 98.605 165.475 ;
        RECT 82.215 164.235 87.560 164.780 ;
        RECT 87.735 164.235 93.080 164.780 ;
        RECT 93.255 164.235 96.765 165.005 ;
        RECT 97.415 164.235 97.655 165.045 ;
        RECT 97.825 164.405 98.155 165.045 ;
        RECT 98.325 164.235 98.595 165.045 ;
        RECT 100.360 164.780 100.700 165.610 ;
        RECT 102.180 165.100 102.530 166.350 ;
        RECT 104.295 165.695 106.885 166.785 ;
        RECT 104.295 165.005 105.505 165.525 ;
        RECT 105.675 165.175 106.885 165.695 ;
        RECT 107.515 165.620 107.805 166.785 ;
        RECT 107.975 165.695 111.485 166.785 ;
        RECT 112.230 166.155 112.515 166.615 ;
        RECT 112.685 166.325 112.955 166.785 ;
        RECT 112.230 165.935 113.185 166.155 ;
        RECT 107.975 165.005 109.625 165.525 ;
        RECT 109.795 165.175 111.485 165.695 ;
        RECT 112.115 165.205 112.805 165.765 ;
        RECT 112.975 165.035 113.185 165.935 ;
        RECT 98.775 164.235 104.120 164.780 ;
        RECT 104.295 164.235 106.885 165.005 ;
        RECT 107.515 164.235 107.805 164.960 ;
        RECT 107.975 164.235 111.485 165.005 ;
        RECT 112.230 164.865 113.185 165.035 ;
        RECT 113.355 165.765 113.755 166.615 ;
        RECT 113.945 166.155 114.225 166.615 ;
        RECT 114.745 166.325 115.070 166.785 ;
        RECT 113.945 165.935 115.070 166.155 ;
        RECT 113.355 165.205 114.450 165.765 ;
        RECT 114.620 165.475 115.070 165.935 ;
        RECT 115.240 165.645 115.625 166.615 ;
        RECT 115.795 165.645 116.085 166.785 ;
        RECT 116.880 166.445 118.245 166.615 ;
        RECT 116.880 166.235 117.210 166.445 ;
        RECT 116.255 165.985 117.210 166.235 ;
        RECT 112.230 164.405 112.515 164.865 ;
        RECT 112.685 164.235 112.955 164.695 ;
        RECT 113.355 164.405 113.755 165.205 ;
        RECT 114.620 165.145 115.175 165.475 ;
        RECT 114.620 165.035 115.070 165.145 ;
        RECT 113.945 164.865 115.070 165.035 ;
        RECT 115.345 164.975 115.625 165.645 ;
        RECT 115.795 165.145 116.070 165.475 ;
        RECT 113.945 164.405 114.225 164.865 ;
        RECT 114.745 164.235 115.070 164.695 ;
        RECT 115.240 164.405 115.625 164.975 ;
        RECT 116.255 164.975 116.425 165.985 ;
        RECT 116.595 165.145 116.950 165.810 ;
        RECT 117.135 165.145 117.410 165.810 ;
        RECT 117.580 165.475 117.905 166.275 ;
        RECT 118.075 165.815 118.245 166.445 ;
        RECT 118.415 165.985 118.705 166.785 ;
        RECT 118.075 165.645 118.750 165.815 ;
        RECT 118.920 165.645 119.305 166.605 ;
        RECT 119.475 165.695 121.145 166.785 ;
        RECT 118.580 165.475 118.750 165.645 ;
        RECT 117.580 165.145 117.925 165.475 ;
        RECT 118.135 165.225 118.385 165.475 ;
        RECT 118.580 165.225 118.945 165.475 ;
        RECT 118.215 165.145 118.385 165.225 ;
        RECT 118.755 165.145 118.945 165.225 ;
        RECT 119.130 164.975 119.305 165.645 ;
        RECT 115.795 164.615 116.085 164.885 ;
        RECT 116.255 164.785 116.680 164.975 ;
        RECT 116.850 164.805 118.250 164.975 ;
        RECT 116.850 164.615 117.180 164.805 ;
        RECT 115.795 164.405 117.180 164.615 ;
        RECT 117.415 164.235 117.745 164.635 ;
        RECT 117.920 164.405 118.250 164.805 ;
        RECT 118.455 164.235 118.625 164.795 ;
        RECT 118.795 164.405 119.305 164.975 ;
        RECT 119.475 165.005 120.225 165.525 ;
        RECT 120.395 165.175 121.145 165.695 ;
        RECT 121.785 165.645 122.115 166.785 ;
        RECT 122.645 165.815 122.975 166.600 ;
        RECT 123.155 165.950 123.500 166.785 ;
        RECT 122.295 165.645 122.975 165.815 ;
        RECT 123.675 165.780 123.930 166.585 ;
        RECT 124.100 165.950 124.360 166.785 ;
        RECT 124.535 165.780 124.790 166.585 ;
        RECT 124.960 165.950 125.220 166.785 ;
        RECT 125.390 165.780 125.650 166.585 ;
        RECT 125.820 165.950 126.205 166.785 ;
        RECT 127.020 165.815 127.410 165.990 ;
        RECT 127.895 165.985 128.225 166.785 ;
        RECT 128.395 165.995 128.930 166.615 ;
        RECT 129.145 166.065 129.475 166.785 ;
        RECT 121.775 165.225 122.125 165.475 ;
        RECT 122.295 165.045 122.465 165.645 ;
        RECT 123.175 165.610 126.205 165.780 ;
        RECT 127.020 165.645 128.445 165.815 ;
        RECT 122.635 165.225 122.985 165.475 ;
        RECT 123.175 165.045 123.345 165.610 ;
        RECT 123.515 165.215 125.730 165.440 ;
        RECT 125.905 165.045 126.205 165.610 ;
        RECT 119.475 164.235 121.145 165.005 ;
        RECT 121.785 164.235 122.055 165.045 ;
        RECT 122.225 164.405 122.555 165.045 ;
        RECT 122.725 164.235 122.965 165.045 ;
        RECT 123.175 164.875 126.205 165.045 ;
        RECT 126.895 164.915 127.250 165.475 ;
        RECT 123.635 164.235 123.930 164.705 ;
        RECT 124.100 164.430 124.360 164.875 ;
        RECT 124.530 164.235 124.790 164.705 ;
        RECT 124.960 164.430 125.215 164.875 ;
        RECT 127.420 164.745 127.590 165.645 ;
        RECT 127.760 164.915 128.025 165.475 ;
        RECT 128.275 165.145 128.445 165.645 ;
        RECT 128.615 164.975 128.930 165.995 ;
        RECT 129.135 165.425 129.365 165.765 ;
        RECT 129.655 165.425 129.870 166.540 ;
        RECT 130.065 165.840 130.395 166.615 ;
        RECT 130.565 166.010 131.275 166.785 ;
        RECT 130.065 165.625 131.215 165.840 ;
        RECT 129.135 165.225 129.465 165.425 ;
        RECT 129.655 165.245 130.105 165.425 ;
        RECT 129.775 165.225 130.105 165.245 ;
        RECT 130.275 165.225 130.745 165.455 ;
        RECT 130.930 165.055 131.215 165.625 ;
        RECT 131.445 165.180 131.725 166.615 ;
        RECT 131.895 165.695 133.105 166.785 ;
        RECT 125.385 164.235 125.685 164.705 ;
        RECT 127.000 164.235 127.240 164.745 ;
        RECT 127.420 164.415 127.700 164.745 ;
        RECT 127.930 164.235 128.145 164.745 ;
        RECT 128.315 164.405 128.930 164.975 ;
        RECT 129.135 164.865 130.315 165.055 ;
        RECT 129.135 164.405 129.475 164.865 ;
        RECT 129.985 164.785 130.315 164.865 ;
        RECT 130.505 164.865 131.215 165.055 ;
        RECT 130.505 164.725 130.805 164.865 ;
        RECT 130.490 164.715 130.805 164.725 ;
        RECT 130.480 164.705 130.805 164.715 ;
        RECT 130.470 164.700 130.805 164.705 ;
        RECT 129.645 164.235 129.815 164.695 ;
        RECT 130.465 164.690 130.805 164.700 ;
        RECT 130.460 164.685 130.805 164.690 ;
        RECT 130.455 164.675 130.805 164.685 ;
        RECT 130.450 164.670 130.805 164.675 ;
        RECT 130.445 164.405 130.805 164.670 ;
        RECT 131.045 164.235 131.215 164.695 ;
        RECT 131.385 164.405 131.725 165.180 ;
        RECT 131.895 164.985 132.415 165.525 ;
        RECT 132.585 165.155 133.105 165.695 ;
        RECT 133.275 165.620 133.565 166.785 ;
        RECT 133.740 165.985 133.995 166.785 ;
        RECT 134.195 165.935 134.525 166.615 ;
        RECT 133.740 165.445 133.985 165.805 ;
        RECT 134.175 165.655 134.525 165.935 ;
        RECT 134.175 165.275 134.345 165.655 ;
        RECT 134.705 165.475 134.900 166.525 ;
        RECT 135.080 165.645 135.400 166.785 ;
        RECT 135.665 165.855 135.835 166.615 ;
        RECT 136.015 166.025 136.345 166.785 ;
        RECT 135.665 165.685 136.330 165.855 ;
        RECT 136.515 165.710 136.785 166.615 ;
        RECT 136.160 165.540 136.330 165.685 ;
        RECT 133.825 165.105 134.345 165.275 ;
        RECT 134.515 165.145 134.900 165.475 ;
        RECT 135.080 165.425 135.340 165.475 ;
        RECT 135.080 165.255 135.345 165.425 ;
        RECT 135.080 165.145 135.340 165.255 ;
        RECT 135.595 165.135 135.925 165.505 ;
        RECT 136.160 165.210 136.445 165.540 ;
        RECT 131.895 164.235 133.105 164.985 ;
        RECT 133.275 164.235 133.565 164.960 ;
        RECT 133.825 164.540 133.995 165.105 ;
        RECT 136.160 164.955 136.330 165.210 ;
        RECT 134.185 164.765 135.400 164.935 ;
        RECT 134.185 164.460 134.415 164.765 ;
        RECT 134.585 164.235 134.915 164.595 ;
        RECT 135.110 164.415 135.400 164.765 ;
        RECT 135.665 164.785 136.330 164.955 ;
        RECT 136.615 164.910 136.785 165.710 ;
        RECT 135.665 164.405 135.835 164.785 ;
        RECT 136.015 164.235 136.345 164.615 ;
        RECT 136.525 164.405 136.785 164.910 ;
        RECT 136.960 165.645 137.295 166.615 ;
        RECT 137.465 165.645 137.635 166.785 ;
        RECT 137.805 166.445 139.835 166.615 ;
        RECT 136.960 164.975 137.130 165.645 ;
        RECT 137.805 165.475 137.975 166.445 ;
        RECT 137.300 165.145 137.555 165.475 ;
        RECT 137.780 165.145 137.975 165.475 ;
        RECT 138.145 166.105 139.270 166.275 ;
        RECT 137.385 164.975 137.555 165.145 ;
        RECT 138.145 164.975 138.315 166.105 ;
        RECT 136.960 164.405 137.215 164.975 ;
        RECT 137.385 164.805 138.315 164.975 ;
        RECT 138.485 165.765 139.495 165.935 ;
        RECT 138.485 164.965 138.655 165.765 ;
        RECT 138.860 165.085 139.135 165.565 ;
        RECT 138.855 164.915 139.135 165.085 ;
        RECT 138.140 164.770 138.315 164.805 ;
        RECT 137.385 164.235 137.715 164.635 ;
        RECT 138.140 164.405 138.670 164.770 ;
        RECT 138.860 164.405 139.135 164.915 ;
        RECT 139.305 164.405 139.495 165.765 ;
        RECT 139.665 165.780 139.835 166.445 ;
        RECT 140.005 166.025 140.175 166.785 ;
        RECT 140.410 166.025 140.925 166.435 ;
        RECT 139.665 165.590 140.415 165.780 ;
        RECT 140.585 165.215 140.925 166.025 ;
        RECT 139.695 165.045 140.925 165.215 ;
        RECT 141.095 165.645 141.480 166.615 ;
        RECT 141.650 166.325 141.975 166.785 ;
        RECT 142.495 166.155 142.775 166.615 ;
        RECT 141.650 165.935 142.775 166.155 ;
        RECT 139.675 164.235 140.185 164.770 ;
        RECT 140.405 164.440 140.650 165.045 ;
        RECT 141.095 164.975 141.375 165.645 ;
        RECT 141.650 165.475 142.100 165.935 ;
        RECT 142.965 165.765 143.365 166.615 ;
        RECT 143.765 166.325 144.035 166.785 ;
        RECT 144.205 166.155 144.490 166.615 ;
        RECT 141.545 165.145 142.100 165.475 ;
        RECT 142.270 165.205 143.365 165.765 ;
        RECT 141.650 165.035 142.100 165.145 ;
        RECT 141.095 164.405 141.480 164.975 ;
        RECT 141.650 164.865 142.775 165.035 ;
        RECT 141.650 164.235 141.975 164.695 ;
        RECT 142.495 164.405 142.775 164.865 ;
        RECT 142.965 164.405 143.365 165.205 ;
        RECT 143.535 165.935 144.490 166.155 ;
        RECT 143.535 165.035 143.745 165.935 ;
        RECT 143.915 165.205 144.605 165.765 ;
        RECT 145.695 165.695 146.905 166.785 ;
        RECT 145.695 165.155 146.215 165.695 ;
        RECT 143.535 164.865 144.490 165.035 ;
        RECT 146.385 164.985 146.905 165.525 ;
        RECT 143.765 164.235 144.035 164.695 ;
        RECT 144.205 164.405 144.490 164.865 ;
        RECT 145.695 164.235 146.905 164.985 ;
        RECT 17.270 164.065 146.990 164.235 ;
        RECT 17.355 163.315 18.565 164.065 ;
        RECT 18.825 163.515 18.995 163.895 ;
        RECT 19.210 163.685 19.540 164.065 ;
        RECT 18.825 163.345 19.540 163.515 ;
        RECT 17.355 162.775 17.875 163.315 ;
        RECT 18.045 162.605 18.565 163.145 ;
        RECT 18.735 162.795 19.090 163.165 ;
        RECT 19.370 163.155 19.540 163.345 ;
        RECT 19.710 163.320 19.965 163.895 ;
        RECT 19.370 162.825 19.625 163.155 ;
        RECT 19.370 162.615 19.540 162.825 ;
        RECT 17.355 161.515 18.565 162.605 ;
        RECT 18.825 162.445 19.540 162.615 ;
        RECT 19.795 162.590 19.965 163.320 ;
        RECT 20.140 163.225 20.400 164.065 ;
        RECT 20.575 163.520 25.920 164.065 ;
        RECT 26.095 163.520 31.440 164.065 ;
        RECT 31.615 163.520 36.960 164.065 ;
        RECT 37.135 163.520 42.480 164.065 ;
        RECT 22.160 162.690 22.500 163.520 ;
        RECT 18.825 161.685 18.995 162.445 ;
        RECT 19.210 161.515 19.540 162.275 ;
        RECT 19.710 161.685 19.965 162.590 ;
        RECT 20.140 161.515 20.400 162.665 ;
        RECT 23.980 161.950 24.330 163.200 ;
        RECT 27.680 162.690 28.020 163.520 ;
        RECT 29.500 161.950 29.850 163.200 ;
        RECT 33.200 162.690 33.540 163.520 ;
        RECT 35.020 161.950 35.370 163.200 ;
        RECT 38.720 162.690 39.060 163.520 ;
        RECT 43.115 163.340 43.405 164.065 ;
        RECT 43.575 163.520 48.920 164.065 ;
        RECT 49.095 163.520 54.440 164.065 ;
        RECT 40.540 161.950 40.890 163.200 ;
        RECT 45.160 162.690 45.500 163.520 ;
        RECT 20.575 161.515 25.920 161.950 ;
        RECT 26.095 161.515 31.440 161.950 ;
        RECT 31.615 161.515 36.960 161.950 ;
        RECT 37.135 161.515 42.480 161.950 ;
        RECT 43.115 161.515 43.405 162.680 ;
        RECT 46.980 161.950 47.330 163.200 ;
        RECT 50.680 162.690 51.020 163.520 ;
        RECT 54.615 163.315 55.825 164.065 ;
        RECT 56.275 163.435 56.655 163.885 ;
        RECT 52.500 161.950 52.850 163.200 ;
        RECT 54.615 162.775 55.135 163.315 ;
        RECT 55.305 162.605 55.825 163.145 ;
        RECT 43.575 161.515 48.920 161.950 ;
        RECT 49.095 161.515 54.440 161.950 ;
        RECT 54.615 161.515 55.825 162.605 ;
        RECT 56.015 162.485 56.245 163.175 ;
        RECT 56.425 162.985 56.655 163.435 ;
        RECT 56.835 163.285 57.065 164.065 ;
        RECT 57.245 163.355 57.675 163.885 ;
        RECT 57.245 163.105 57.490 163.355 ;
        RECT 57.855 163.155 58.065 163.775 ;
        RECT 58.235 163.335 58.565 164.065 ;
        RECT 58.845 163.515 59.015 163.805 ;
        RECT 59.185 163.685 59.515 164.065 ;
        RECT 58.845 163.345 59.510 163.515 ;
        RECT 56.425 162.305 56.765 162.985 ;
        RECT 56.005 162.105 56.765 162.305 ;
        RECT 56.955 162.805 57.490 163.105 ;
        RECT 57.670 162.805 58.065 163.155 ;
        RECT 58.260 162.805 58.550 163.155 ;
        RECT 56.005 161.715 56.265 162.105 ;
        RECT 56.435 161.515 56.765 161.925 ;
        RECT 56.955 161.695 57.285 162.805 ;
        RECT 57.455 162.425 58.495 162.625 ;
        RECT 58.760 162.525 59.110 163.175 ;
        RECT 57.455 161.695 57.645 162.425 ;
        RECT 57.815 161.515 58.145 162.245 ;
        RECT 58.325 161.695 58.495 162.425 ;
        RECT 59.280 162.355 59.510 163.345 ;
        RECT 58.845 162.185 59.510 162.355 ;
        RECT 58.845 161.685 59.015 162.185 ;
        RECT 59.185 161.515 59.515 162.015 ;
        RECT 59.685 161.685 59.870 163.805 ;
        RECT 60.125 163.605 60.375 164.065 ;
        RECT 60.545 163.615 60.880 163.785 ;
        RECT 61.075 163.615 61.750 163.785 ;
        RECT 60.545 163.475 60.715 163.615 ;
        RECT 60.040 162.485 60.320 163.435 ;
        RECT 60.490 163.345 60.715 163.475 ;
        RECT 60.490 162.240 60.660 163.345 ;
        RECT 60.885 163.195 61.410 163.415 ;
        RECT 60.830 162.430 61.070 163.025 ;
        RECT 61.240 162.495 61.410 163.195 ;
        RECT 61.580 162.835 61.750 163.615 ;
        RECT 62.070 163.565 62.440 164.065 ;
        RECT 62.620 163.615 63.025 163.785 ;
        RECT 63.195 163.615 63.980 163.785 ;
        RECT 62.620 163.385 62.790 163.615 ;
        RECT 61.960 163.085 62.790 163.385 ;
        RECT 63.175 163.115 63.640 163.445 ;
        RECT 61.960 163.055 62.160 163.085 ;
        RECT 62.280 162.835 62.450 162.905 ;
        RECT 61.580 162.665 62.450 162.835 ;
        RECT 61.940 162.575 62.450 162.665 ;
        RECT 60.490 162.110 60.795 162.240 ;
        RECT 61.240 162.130 61.770 162.495 ;
        RECT 60.110 161.515 60.375 161.975 ;
        RECT 60.545 161.685 60.795 162.110 ;
        RECT 61.940 161.960 62.110 162.575 ;
        RECT 61.005 161.790 62.110 161.960 ;
        RECT 62.280 161.515 62.450 162.315 ;
        RECT 62.620 162.015 62.790 163.085 ;
        RECT 62.960 162.185 63.150 162.905 ;
        RECT 63.320 162.155 63.640 163.115 ;
        RECT 63.810 163.155 63.980 163.615 ;
        RECT 64.255 163.535 64.465 164.065 ;
        RECT 64.725 163.325 65.055 163.850 ;
        RECT 65.225 163.455 65.395 164.065 ;
        RECT 65.565 163.410 65.895 163.845 ;
        RECT 66.120 163.560 66.455 164.065 ;
        RECT 66.625 163.495 66.865 163.870 ;
        RECT 67.145 163.735 67.315 163.880 ;
        RECT 67.145 163.540 67.520 163.735 ;
        RECT 67.880 163.570 68.275 164.065 ;
        RECT 65.565 163.325 65.945 163.410 ;
        RECT 64.855 163.155 65.055 163.325 ;
        RECT 65.720 163.285 65.945 163.325 ;
        RECT 63.810 162.825 64.685 163.155 ;
        RECT 64.855 162.825 65.605 163.155 ;
        RECT 62.620 161.685 62.870 162.015 ;
        RECT 63.810 161.985 63.980 162.825 ;
        RECT 64.855 162.620 65.045 162.825 ;
        RECT 65.775 162.705 65.945 163.285 ;
        RECT 65.730 162.655 65.945 162.705 ;
        RECT 64.150 162.245 65.045 162.620 ;
        RECT 65.555 162.575 65.945 162.655 ;
        RECT 63.095 161.815 63.980 161.985 ;
        RECT 64.160 161.515 64.475 162.015 ;
        RECT 64.705 161.685 65.045 162.245 ;
        RECT 65.215 161.515 65.385 162.525 ;
        RECT 65.555 161.730 65.885 162.575 ;
        RECT 66.175 162.535 66.475 163.385 ;
        RECT 66.645 163.345 66.865 163.495 ;
        RECT 66.645 163.015 67.180 163.345 ;
        RECT 67.350 163.205 67.520 163.540 ;
        RECT 68.445 163.375 68.685 163.895 ;
        RECT 66.645 162.365 66.880 163.015 ;
        RECT 67.350 162.845 68.335 163.205 ;
        RECT 66.205 162.135 66.880 162.365 ;
        RECT 67.050 162.825 68.335 162.845 ;
        RECT 67.050 162.675 67.910 162.825 ;
        RECT 66.205 161.705 66.375 162.135 ;
        RECT 66.545 161.515 66.875 161.965 ;
        RECT 67.050 161.730 67.335 162.675 ;
        RECT 68.510 162.570 68.685 163.375 ;
        RECT 68.875 163.340 69.165 164.065 ;
        RECT 69.335 163.435 69.675 163.895 ;
        RECT 69.845 163.605 70.015 164.065 ;
        RECT 70.645 163.630 71.005 163.895 ;
        RECT 70.650 163.625 71.005 163.630 ;
        RECT 70.655 163.615 71.005 163.625 ;
        RECT 70.660 163.610 71.005 163.615 ;
        RECT 70.665 163.600 71.005 163.610 ;
        RECT 71.245 163.605 71.415 164.065 ;
        RECT 70.670 163.595 71.005 163.600 ;
        RECT 70.680 163.585 71.005 163.595 ;
        RECT 70.690 163.575 71.005 163.585 ;
        RECT 70.185 163.435 70.515 163.515 ;
        RECT 69.335 163.245 70.515 163.435 ;
        RECT 70.705 163.435 71.005 163.575 ;
        RECT 70.705 163.245 71.415 163.435 ;
        RECT 69.335 162.875 69.665 163.075 ;
        RECT 69.975 163.055 70.305 163.075 ;
        RECT 69.855 162.875 70.305 163.055 ;
        RECT 67.510 162.195 68.205 162.505 ;
        RECT 67.515 161.515 68.200 161.985 ;
        RECT 68.380 161.785 68.685 162.570 ;
        RECT 68.875 161.515 69.165 162.680 ;
        RECT 69.335 162.535 69.565 162.875 ;
        RECT 69.345 161.515 69.675 162.235 ;
        RECT 69.855 161.760 70.070 162.875 ;
        RECT 70.475 162.845 70.945 163.075 ;
        RECT 71.130 162.675 71.415 163.245 ;
        RECT 71.585 163.120 71.925 163.895 ;
        RECT 72.210 163.435 72.495 163.895 ;
        RECT 72.665 163.605 72.935 164.065 ;
        RECT 72.210 163.265 73.165 163.435 ;
        RECT 70.265 162.460 71.415 162.675 ;
        RECT 70.265 161.685 70.595 162.460 ;
        RECT 70.765 161.515 71.475 162.290 ;
        RECT 71.645 161.685 71.925 163.120 ;
        RECT 72.095 162.535 72.785 163.095 ;
        RECT 72.955 162.365 73.165 163.265 ;
        RECT 72.210 162.145 73.165 162.365 ;
        RECT 73.335 163.095 73.735 163.895 ;
        RECT 73.925 163.435 74.205 163.895 ;
        RECT 74.725 163.605 75.050 164.065 ;
        RECT 73.925 163.265 75.050 163.435 ;
        RECT 75.220 163.325 75.605 163.895 ;
        RECT 75.865 163.515 76.035 163.805 ;
        RECT 76.205 163.685 76.535 164.065 ;
        RECT 75.865 163.345 76.530 163.515 ;
        RECT 74.600 163.155 75.050 163.265 ;
        RECT 73.335 162.535 74.430 163.095 ;
        RECT 74.600 162.825 75.155 163.155 ;
        RECT 72.210 161.685 72.495 162.145 ;
        RECT 72.665 161.515 72.935 161.975 ;
        RECT 73.335 161.685 73.735 162.535 ;
        RECT 74.600 162.365 75.050 162.825 ;
        RECT 75.325 162.655 75.605 163.325 ;
        RECT 73.925 162.145 75.050 162.365 ;
        RECT 73.925 161.685 74.205 162.145 ;
        RECT 74.725 161.515 75.050 161.975 ;
        RECT 75.220 161.685 75.605 162.655 ;
        RECT 75.780 162.525 76.130 163.175 ;
        RECT 76.300 162.355 76.530 163.345 ;
        RECT 75.865 162.185 76.530 162.355 ;
        RECT 75.865 161.685 76.035 162.185 ;
        RECT 76.205 161.515 76.535 162.015 ;
        RECT 76.705 161.685 76.890 163.805 ;
        RECT 77.145 163.605 77.395 164.065 ;
        RECT 77.565 163.615 77.900 163.785 ;
        RECT 78.095 163.615 78.770 163.785 ;
        RECT 77.565 163.475 77.735 163.615 ;
        RECT 77.060 162.485 77.340 163.435 ;
        RECT 77.510 163.345 77.735 163.475 ;
        RECT 77.510 162.240 77.680 163.345 ;
        RECT 77.905 163.195 78.430 163.415 ;
        RECT 77.850 162.430 78.090 163.025 ;
        RECT 78.260 162.495 78.430 163.195 ;
        RECT 78.600 162.835 78.770 163.615 ;
        RECT 79.090 163.565 79.460 164.065 ;
        RECT 79.640 163.615 80.045 163.785 ;
        RECT 80.215 163.615 81.000 163.785 ;
        RECT 79.640 163.385 79.810 163.615 ;
        RECT 78.980 163.085 79.810 163.385 ;
        RECT 80.195 163.115 80.660 163.445 ;
        RECT 78.980 163.055 79.180 163.085 ;
        RECT 79.300 162.835 79.470 162.905 ;
        RECT 78.600 162.665 79.470 162.835 ;
        RECT 78.960 162.575 79.470 162.665 ;
        RECT 77.510 162.110 77.815 162.240 ;
        RECT 78.260 162.130 78.790 162.495 ;
        RECT 77.130 161.515 77.395 161.975 ;
        RECT 77.565 161.685 77.815 162.110 ;
        RECT 78.960 161.960 79.130 162.575 ;
        RECT 78.025 161.790 79.130 161.960 ;
        RECT 79.300 161.515 79.470 162.315 ;
        RECT 79.640 162.015 79.810 163.085 ;
        RECT 79.980 162.185 80.170 162.905 ;
        RECT 80.340 162.155 80.660 163.115 ;
        RECT 80.830 163.155 81.000 163.615 ;
        RECT 81.275 163.535 81.485 164.065 ;
        RECT 81.745 163.325 82.075 163.850 ;
        RECT 82.245 163.455 82.415 164.065 ;
        RECT 82.585 163.410 82.915 163.845 ;
        RECT 82.585 163.325 82.965 163.410 ;
        RECT 81.875 163.155 82.075 163.325 ;
        RECT 82.740 163.285 82.965 163.325 ;
        RECT 80.830 162.825 81.705 163.155 ;
        RECT 81.875 162.825 82.625 163.155 ;
        RECT 79.640 161.685 79.890 162.015 ;
        RECT 80.830 161.985 81.000 162.825 ;
        RECT 81.875 162.620 82.065 162.825 ;
        RECT 82.795 162.705 82.965 163.285 ;
        RECT 82.750 162.655 82.965 162.705 ;
        RECT 81.170 162.245 82.065 162.620 ;
        RECT 82.575 162.575 82.965 162.655 ;
        RECT 83.135 163.325 83.520 163.895 ;
        RECT 83.690 163.605 84.015 164.065 ;
        RECT 84.535 163.435 84.815 163.895 ;
        RECT 83.135 162.655 83.415 163.325 ;
        RECT 83.690 163.265 84.815 163.435 ;
        RECT 83.690 163.155 84.140 163.265 ;
        RECT 83.585 162.825 84.140 163.155 ;
        RECT 85.005 163.095 85.405 163.895 ;
        RECT 85.805 163.605 86.075 164.065 ;
        RECT 86.245 163.435 86.530 163.895 ;
        RECT 86.835 163.555 87.075 164.065 ;
        RECT 87.245 163.555 87.535 163.895 ;
        RECT 87.765 163.555 88.080 164.065 ;
        RECT 80.115 161.815 81.000 161.985 ;
        RECT 81.180 161.515 81.495 162.015 ;
        RECT 81.725 161.685 82.065 162.245 ;
        RECT 82.235 161.515 82.405 162.525 ;
        RECT 82.575 161.730 82.905 162.575 ;
        RECT 83.135 161.685 83.520 162.655 ;
        RECT 83.690 162.365 84.140 162.825 ;
        RECT 84.310 162.535 85.405 163.095 ;
        RECT 83.690 162.145 84.815 162.365 ;
        RECT 83.690 161.515 84.015 161.975 ;
        RECT 84.535 161.685 84.815 162.145 ;
        RECT 85.005 161.685 85.405 162.535 ;
        RECT 85.575 163.265 86.530 163.435 ;
        RECT 85.575 162.365 85.785 163.265 ;
        RECT 85.955 162.535 86.645 163.095 ;
        RECT 86.880 163.045 87.075 163.385 ;
        RECT 86.875 162.875 87.075 163.045 ;
        RECT 86.880 162.825 87.075 162.875 ;
        RECT 87.245 162.655 87.425 163.555 ;
        RECT 88.250 163.495 88.420 163.765 ;
        RECT 88.590 163.665 88.920 164.065 ;
        RECT 90.515 163.595 90.810 164.065 ;
        RECT 87.595 162.825 88.005 163.385 ;
        RECT 88.250 163.325 88.945 163.495 ;
        RECT 90.980 163.425 91.240 163.870 ;
        RECT 91.410 163.595 91.670 164.065 ;
        RECT 91.840 163.425 92.095 163.870 ;
        RECT 92.265 163.595 92.565 164.065 ;
        RECT 88.175 162.655 88.345 163.155 ;
        RECT 86.885 162.485 88.345 162.655 ;
        RECT 85.575 162.145 86.530 162.365 ;
        RECT 86.885 162.310 87.245 162.485 ;
        RECT 88.515 162.315 88.945 163.325 ;
        RECT 90.055 163.255 93.085 163.425 ;
        RECT 90.055 162.690 90.225 163.255 ;
        RECT 90.395 162.860 92.610 163.085 ;
        RECT 92.785 162.690 93.085 163.255 ;
        RECT 93.255 163.315 94.465 164.065 ;
        RECT 94.635 163.340 94.925 164.065 ;
        RECT 95.095 163.520 100.440 164.065 ;
        RECT 93.255 162.775 93.775 163.315 ;
        RECT 90.055 162.520 93.085 162.690 ;
        RECT 93.945 162.605 94.465 163.145 ;
        RECT 96.680 162.690 97.020 163.520 ;
        RECT 100.615 163.295 102.285 164.065 ;
        RECT 103.005 163.515 103.175 163.805 ;
        RECT 103.345 163.685 103.675 164.065 ;
        RECT 103.005 163.345 103.670 163.515 ;
        RECT 85.805 161.515 86.075 161.975 ;
        RECT 86.245 161.685 86.530 162.145 ;
        RECT 87.830 161.515 88.000 162.315 ;
        RECT 88.170 162.145 88.945 162.315 ;
        RECT 88.170 161.685 88.500 162.145 ;
        RECT 88.670 161.515 88.840 161.975 ;
        RECT 90.035 161.515 90.380 162.350 ;
        RECT 90.555 161.715 90.810 162.520 ;
        RECT 90.980 161.515 91.240 162.350 ;
        RECT 91.415 161.715 91.670 162.520 ;
        RECT 91.840 161.515 92.100 162.350 ;
        RECT 92.270 161.715 92.530 162.520 ;
        RECT 92.700 161.515 93.085 162.350 ;
        RECT 93.255 161.515 94.465 162.605 ;
        RECT 94.635 161.515 94.925 162.680 ;
        RECT 98.500 161.950 98.850 163.200 ;
        RECT 100.615 162.775 101.365 163.295 ;
        RECT 101.535 162.605 102.285 163.125 ;
        RECT 95.095 161.515 100.440 161.950 ;
        RECT 100.615 161.515 102.285 162.605 ;
        RECT 102.920 162.525 103.270 163.175 ;
        RECT 103.440 162.355 103.670 163.345 ;
        RECT 103.005 162.185 103.670 162.355 ;
        RECT 103.005 161.685 103.175 162.185 ;
        RECT 103.345 161.515 103.675 162.015 ;
        RECT 103.845 161.685 104.030 163.805 ;
        RECT 104.285 163.605 104.535 164.065 ;
        RECT 104.705 163.615 105.040 163.785 ;
        RECT 105.235 163.615 105.910 163.785 ;
        RECT 104.705 163.475 104.875 163.615 ;
        RECT 104.200 162.485 104.480 163.435 ;
        RECT 104.650 163.345 104.875 163.475 ;
        RECT 104.650 162.240 104.820 163.345 ;
        RECT 105.045 163.195 105.570 163.415 ;
        RECT 104.990 162.430 105.230 163.025 ;
        RECT 105.400 162.495 105.570 163.195 ;
        RECT 105.740 162.835 105.910 163.615 ;
        RECT 106.230 163.565 106.600 164.065 ;
        RECT 106.780 163.615 107.185 163.785 ;
        RECT 107.355 163.615 108.140 163.785 ;
        RECT 106.780 163.385 106.950 163.615 ;
        RECT 106.120 163.085 106.950 163.385 ;
        RECT 107.335 163.115 107.800 163.445 ;
        RECT 106.120 163.055 106.320 163.085 ;
        RECT 106.440 162.835 106.610 162.905 ;
        RECT 105.740 162.665 106.610 162.835 ;
        RECT 106.100 162.575 106.610 162.665 ;
        RECT 104.650 162.110 104.955 162.240 ;
        RECT 105.400 162.130 105.930 162.495 ;
        RECT 104.270 161.515 104.535 161.975 ;
        RECT 104.705 161.685 104.955 162.110 ;
        RECT 106.100 161.960 106.270 162.575 ;
        RECT 105.165 161.790 106.270 161.960 ;
        RECT 106.440 161.515 106.610 162.315 ;
        RECT 106.780 162.015 106.950 163.085 ;
        RECT 107.120 162.185 107.310 162.905 ;
        RECT 107.480 162.155 107.800 163.115 ;
        RECT 107.970 163.155 108.140 163.615 ;
        RECT 108.415 163.535 108.625 164.065 ;
        RECT 108.885 163.325 109.215 163.850 ;
        RECT 109.385 163.455 109.555 164.065 ;
        RECT 109.725 163.410 110.055 163.845 ;
        RECT 111.195 163.565 111.455 163.895 ;
        RECT 111.625 163.705 111.955 164.065 ;
        RECT 112.210 163.685 113.510 163.895 ;
        RECT 111.195 163.555 111.425 163.565 ;
        RECT 109.725 163.325 110.105 163.410 ;
        RECT 109.015 163.155 109.215 163.325 ;
        RECT 109.880 163.285 110.105 163.325 ;
        RECT 107.970 162.825 108.845 163.155 ;
        RECT 109.015 162.825 109.765 163.155 ;
        RECT 106.780 161.685 107.030 162.015 ;
        RECT 107.970 161.985 108.140 162.825 ;
        RECT 109.015 162.620 109.205 162.825 ;
        RECT 109.935 162.705 110.105 163.285 ;
        RECT 109.890 162.655 110.105 162.705 ;
        RECT 108.310 162.245 109.205 162.620 ;
        RECT 109.715 162.575 110.105 162.655 ;
        RECT 107.255 161.815 108.140 161.985 ;
        RECT 108.320 161.515 108.635 162.015 ;
        RECT 108.865 161.685 109.205 162.245 ;
        RECT 109.375 161.515 109.545 162.525 ;
        RECT 109.715 161.730 110.045 162.575 ;
        RECT 111.195 162.365 111.365 163.555 ;
        RECT 112.210 163.535 112.380 163.685 ;
        RECT 111.625 163.410 112.380 163.535 ;
        RECT 111.535 163.365 112.380 163.410 ;
        RECT 111.535 163.245 111.805 163.365 ;
        RECT 111.535 162.670 111.705 163.245 ;
        RECT 111.935 162.805 112.345 163.110 ;
        RECT 112.635 163.075 112.845 163.475 ;
        RECT 112.515 162.865 112.845 163.075 ;
        RECT 113.090 163.075 113.310 163.475 ;
        RECT 113.785 163.300 114.240 164.065 ;
        RECT 114.420 163.390 114.695 163.735 ;
        RECT 114.885 163.665 115.265 164.065 ;
        RECT 115.435 163.495 115.605 163.845 ;
        RECT 115.775 163.665 116.105 164.065 ;
        RECT 116.275 163.495 116.530 163.845 ;
        RECT 113.090 162.865 113.565 163.075 ;
        RECT 113.755 162.875 114.245 163.075 ;
        RECT 111.535 162.635 111.735 162.670 ;
        RECT 113.065 162.635 114.240 162.695 ;
        RECT 111.535 162.525 114.240 162.635 ;
        RECT 111.595 162.465 113.395 162.525 ;
        RECT 113.065 162.435 113.395 162.465 ;
        RECT 111.195 161.685 111.455 162.365 ;
        RECT 111.625 161.515 111.875 162.295 ;
        RECT 112.125 162.265 112.960 162.275 ;
        RECT 113.550 162.265 113.735 162.355 ;
        RECT 112.125 162.065 113.735 162.265 ;
        RECT 112.125 161.685 112.375 162.065 ;
        RECT 113.505 162.025 113.735 162.065 ;
        RECT 113.985 161.905 114.240 162.525 ;
        RECT 112.545 161.515 112.900 161.895 ;
        RECT 113.905 161.685 114.240 161.905 ;
        RECT 114.420 162.655 114.590 163.390 ;
        RECT 114.865 163.325 116.530 163.495 ;
        RECT 114.865 163.155 115.035 163.325 ;
        RECT 116.755 163.245 116.985 164.065 ;
        RECT 117.155 163.265 117.485 163.895 ;
        RECT 114.760 162.825 115.035 163.155 ;
        RECT 115.205 162.825 116.030 163.155 ;
        RECT 116.200 162.825 116.545 163.155 ;
        RECT 116.735 162.825 117.065 163.075 ;
        RECT 114.865 162.655 115.035 162.825 ;
        RECT 114.420 161.685 114.695 162.655 ;
        RECT 114.865 162.485 115.525 162.655 ;
        RECT 115.835 162.535 116.030 162.825 ;
        RECT 117.235 162.665 117.485 163.265 ;
        RECT 117.655 163.245 117.865 164.065 ;
        RECT 118.260 163.555 118.500 164.065 ;
        RECT 118.680 163.555 118.960 163.885 ;
        RECT 119.190 163.555 119.405 164.065 ;
        RECT 118.155 162.825 118.510 163.385 ;
        RECT 115.355 162.365 115.525 162.485 ;
        RECT 116.200 162.365 116.525 162.655 ;
        RECT 114.905 161.515 115.185 162.315 ;
        RECT 115.355 162.195 116.525 162.365 ;
        RECT 115.355 161.735 116.545 162.025 ;
        RECT 116.755 161.515 116.985 162.655 ;
        RECT 117.155 161.685 117.485 162.665 ;
        RECT 118.680 162.655 118.850 163.555 ;
        RECT 119.020 162.825 119.285 163.385 ;
        RECT 119.575 163.325 120.190 163.895 ;
        RECT 120.395 163.340 120.685 164.065 ;
        RECT 119.535 162.655 119.705 163.155 ;
        RECT 117.655 161.515 117.865 162.655 ;
        RECT 118.280 162.485 119.705 162.655 ;
        RECT 118.280 162.310 118.670 162.485 ;
        RECT 119.155 161.515 119.485 162.315 ;
        RECT 119.875 162.305 120.190 163.325 ;
        RECT 120.860 163.300 121.315 164.065 ;
        RECT 121.590 163.685 122.890 163.895 ;
        RECT 123.145 163.705 123.475 164.065 ;
        RECT 122.720 163.535 122.890 163.685 ;
        RECT 123.645 163.565 123.905 163.895 ;
        RECT 123.675 163.555 123.905 163.565 ;
        RECT 121.790 163.075 122.010 163.475 ;
        RECT 120.855 162.875 121.345 163.075 ;
        RECT 121.535 162.865 122.010 163.075 ;
        RECT 122.255 163.075 122.465 163.475 ;
        RECT 122.720 163.410 123.475 163.535 ;
        RECT 122.720 163.365 123.565 163.410 ;
        RECT 123.295 163.245 123.565 163.365 ;
        RECT 122.255 162.865 122.585 163.075 ;
        RECT 122.755 162.805 123.165 163.110 ;
        RECT 119.655 161.685 120.190 162.305 ;
        RECT 120.395 161.515 120.685 162.680 ;
        RECT 120.860 162.635 122.035 162.695 ;
        RECT 123.395 162.670 123.565 163.245 ;
        RECT 123.365 162.635 123.565 162.670 ;
        RECT 120.860 162.525 123.565 162.635 ;
        RECT 120.860 161.905 121.115 162.525 ;
        RECT 121.705 162.465 123.505 162.525 ;
        RECT 121.705 162.435 122.035 162.465 ;
        RECT 123.735 162.365 123.905 163.555 ;
        RECT 124.075 163.520 129.420 164.065 ;
        RECT 125.660 162.690 126.000 163.520 ;
        RECT 129.685 163.515 129.855 163.895 ;
        RECT 130.035 163.685 130.365 164.065 ;
        RECT 129.685 163.345 130.350 163.515 ;
        RECT 130.545 163.390 130.805 163.895 ;
        RECT 121.365 162.265 121.550 162.355 ;
        RECT 122.140 162.265 122.975 162.275 ;
        RECT 121.365 162.065 122.975 162.265 ;
        RECT 121.365 162.025 121.595 162.065 ;
        RECT 120.860 161.685 121.195 161.905 ;
        RECT 122.200 161.515 122.555 161.895 ;
        RECT 122.725 161.685 122.975 162.065 ;
        RECT 123.225 161.515 123.475 162.295 ;
        RECT 123.645 161.685 123.905 162.365 ;
        RECT 127.480 161.950 127.830 163.200 ;
        RECT 129.615 162.795 129.945 163.165 ;
        RECT 130.180 163.090 130.350 163.345 ;
        RECT 130.180 162.760 130.465 163.090 ;
        RECT 130.180 162.615 130.350 162.760 ;
        RECT 129.685 162.445 130.350 162.615 ;
        RECT 130.635 162.590 130.805 163.390 ;
        RECT 130.980 163.225 131.240 164.065 ;
        RECT 131.415 163.320 131.670 163.895 ;
        RECT 131.840 163.685 132.170 164.065 ;
        RECT 132.385 163.515 132.555 163.895 ;
        RECT 131.840 163.345 132.555 163.515 ;
        RECT 124.075 161.515 129.420 161.950 ;
        RECT 129.685 161.685 129.855 162.445 ;
        RECT 130.035 161.515 130.365 162.275 ;
        RECT 130.535 161.685 130.805 162.590 ;
        RECT 130.980 161.515 131.240 162.665 ;
        RECT 131.415 162.590 131.585 163.320 ;
        RECT 131.840 163.155 132.010 163.345 ;
        RECT 132.820 163.225 133.080 164.065 ;
        RECT 133.255 163.320 133.510 163.895 ;
        RECT 133.680 163.685 134.010 164.065 ;
        RECT 134.225 163.515 134.395 163.895 ;
        RECT 133.680 163.345 134.395 163.515 ;
        RECT 131.755 162.825 132.010 163.155 ;
        RECT 131.840 162.615 132.010 162.825 ;
        RECT 132.290 162.795 132.645 163.165 ;
        RECT 131.415 161.685 131.670 162.590 ;
        RECT 131.840 162.445 132.555 162.615 ;
        RECT 131.840 161.515 132.170 162.275 ;
        RECT 132.385 161.685 132.555 162.445 ;
        RECT 132.820 161.515 133.080 162.665 ;
        RECT 133.255 162.590 133.425 163.320 ;
        RECT 133.680 163.155 133.850 163.345 ;
        RECT 134.660 163.325 134.915 163.895 ;
        RECT 135.085 163.665 135.415 164.065 ;
        RECT 135.840 163.530 136.370 163.895 ;
        RECT 135.840 163.495 136.015 163.530 ;
        RECT 135.085 163.325 136.015 163.495 ;
        RECT 133.595 162.825 133.850 163.155 ;
        RECT 133.680 162.615 133.850 162.825 ;
        RECT 134.130 162.795 134.485 163.165 ;
        RECT 134.660 162.655 134.830 163.325 ;
        RECT 135.085 163.155 135.255 163.325 ;
        RECT 135.000 162.825 135.255 163.155 ;
        RECT 135.480 162.825 135.675 163.155 ;
        RECT 133.255 161.685 133.510 162.590 ;
        RECT 133.680 162.445 134.395 162.615 ;
        RECT 133.680 161.515 134.010 162.275 ;
        RECT 134.225 161.685 134.395 162.445 ;
        RECT 134.660 161.685 134.995 162.655 ;
        RECT 135.165 161.515 135.335 162.655 ;
        RECT 135.505 161.855 135.675 162.825 ;
        RECT 135.845 162.195 136.015 163.325 ;
        RECT 136.185 162.535 136.355 163.335 ;
        RECT 136.560 163.045 136.835 163.895 ;
        RECT 136.555 162.875 136.835 163.045 ;
        RECT 136.560 162.735 136.835 162.875 ;
        RECT 137.005 162.535 137.195 163.895 ;
        RECT 137.375 163.530 137.885 164.065 ;
        RECT 138.105 163.255 138.350 163.860 ;
        RECT 138.795 163.325 139.180 163.895 ;
        RECT 139.350 163.605 139.675 164.065 ;
        RECT 140.195 163.435 140.475 163.895 ;
        RECT 137.395 163.085 138.625 163.255 ;
        RECT 136.185 162.365 137.195 162.535 ;
        RECT 137.365 162.520 138.115 162.710 ;
        RECT 135.845 162.025 136.970 162.195 ;
        RECT 137.365 161.855 137.535 162.520 ;
        RECT 138.285 162.275 138.625 163.085 ;
        RECT 135.505 161.685 137.535 161.855 ;
        RECT 137.705 161.515 137.875 162.275 ;
        RECT 138.110 161.865 138.625 162.275 ;
        RECT 138.795 162.655 139.075 163.325 ;
        RECT 139.350 163.265 140.475 163.435 ;
        RECT 139.350 163.155 139.800 163.265 ;
        RECT 139.245 162.825 139.800 163.155 ;
        RECT 140.665 163.095 141.065 163.895 ;
        RECT 141.465 163.605 141.735 164.065 ;
        RECT 141.905 163.435 142.190 163.895 ;
        RECT 138.795 161.685 139.180 162.655 ;
        RECT 139.350 162.365 139.800 162.825 ;
        RECT 139.970 162.535 141.065 163.095 ;
        RECT 139.350 162.145 140.475 162.365 ;
        RECT 139.350 161.515 139.675 161.975 ;
        RECT 140.195 161.685 140.475 162.145 ;
        RECT 140.665 161.685 141.065 162.535 ;
        RECT 141.235 163.265 142.190 163.435 ;
        RECT 142.565 163.515 142.735 163.895 ;
        RECT 142.915 163.685 143.245 164.065 ;
        RECT 142.565 163.345 143.230 163.515 ;
        RECT 143.425 163.390 143.685 163.895 ;
        RECT 141.235 162.365 141.445 163.265 ;
        RECT 141.615 162.535 142.305 163.095 ;
        RECT 142.495 162.795 142.825 163.165 ;
        RECT 143.060 163.090 143.230 163.345 ;
        RECT 143.060 162.760 143.345 163.090 ;
        RECT 143.060 162.615 143.230 162.760 ;
        RECT 142.565 162.445 143.230 162.615 ;
        RECT 143.515 162.590 143.685 163.390 ;
        RECT 143.945 163.515 144.115 163.895 ;
        RECT 144.330 163.685 144.660 164.065 ;
        RECT 143.945 163.345 144.660 163.515 ;
        RECT 143.855 162.795 144.210 163.165 ;
        RECT 144.490 163.155 144.660 163.345 ;
        RECT 144.830 163.320 145.085 163.895 ;
        RECT 144.490 162.825 144.745 163.155 ;
        RECT 144.490 162.615 144.660 162.825 ;
        RECT 141.235 162.145 142.190 162.365 ;
        RECT 141.465 161.515 141.735 161.975 ;
        RECT 141.905 161.685 142.190 162.145 ;
        RECT 142.565 161.685 142.735 162.445 ;
        RECT 142.915 161.515 143.245 162.275 ;
        RECT 143.415 161.685 143.685 162.590 ;
        RECT 143.945 162.445 144.660 162.615 ;
        RECT 144.915 162.590 145.085 163.320 ;
        RECT 145.260 163.225 145.520 164.065 ;
        RECT 145.695 163.315 146.905 164.065 ;
        RECT 143.945 161.685 144.115 162.445 ;
        RECT 144.330 161.515 144.660 162.275 ;
        RECT 144.830 161.685 145.085 162.590 ;
        RECT 145.260 161.515 145.520 162.665 ;
        RECT 145.695 162.605 146.215 163.145 ;
        RECT 146.385 162.775 146.905 163.315 ;
        RECT 145.695 161.515 146.905 162.605 ;
        RECT 17.270 161.345 146.990 161.515 ;
        RECT 17.355 160.255 18.565 161.345 ;
        RECT 18.735 160.910 24.080 161.345 ;
        RECT 24.255 160.910 29.600 161.345 ;
        RECT 17.355 159.545 17.875 160.085 ;
        RECT 18.045 159.715 18.565 160.255 ;
        RECT 17.355 158.795 18.565 159.545 ;
        RECT 20.320 159.340 20.660 160.170 ;
        RECT 22.140 159.660 22.490 160.910 ;
        RECT 25.840 159.340 26.180 160.170 ;
        RECT 27.660 159.660 28.010 160.910 ;
        RECT 30.235 160.180 30.525 161.345 ;
        RECT 30.695 160.255 33.285 161.345 ;
        RECT 30.695 159.565 31.905 160.085 ;
        RECT 32.075 159.735 33.285 160.255 ;
        RECT 33.950 160.555 34.485 161.175 ;
        RECT 18.735 158.795 24.080 159.340 ;
        RECT 24.255 158.795 29.600 159.340 ;
        RECT 30.235 158.795 30.525 159.520 ;
        RECT 30.695 158.795 33.285 159.565 ;
        RECT 33.950 159.535 34.265 160.555 ;
        RECT 34.655 160.545 34.985 161.345 ;
        RECT 35.470 160.375 35.860 160.550 ;
        RECT 34.435 160.205 35.860 160.375 ;
        RECT 36.215 160.475 36.490 161.175 ;
        RECT 36.660 160.800 36.915 161.345 ;
        RECT 37.085 160.835 37.565 161.175 ;
        RECT 37.740 160.790 38.345 161.345 ;
        RECT 37.730 160.690 38.345 160.790 ;
        RECT 37.730 160.665 37.915 160.690 ;
        RECT 34.435 159.705 34.605 160.205 ;
        RECT 33.950 158.965 34.565 159.535 ;
        RECT 34.855 159.475 35.120 160.035 ;
        RECT 35.290 159.305 35.460 160.205 ;
        RECT 35.630 159.475 35.985 160.035 ;
        RECT 36.215 159.445 36.385 160.475 ;
        RECT 36.660 160.345 37.415 160.595 ;
        RECT 37.585 160.420 37.915 160.665 ;
        RECT 36.660 160.310 37.430 160.345 ;
        RECT 36.660 160.300 37.445 160.310 ;
        RECT 36.555 160.285 37.450 160.300 ;
        RECT 36.555 160.270 37.470 160.285 ;
        RECT 36.555 160.260 37.490 160.270 ;
        RECT 36.555 160.250 37.515 160.260 ;
        RECT 36.555 160.220 37.585 160.250 ;
        RECT 36.555 160.190 37.605 160.220 ;
        RECT 36.555 160.160 37.625 160.190 ;
        RECT 36.555 160.135 37.655 160.160 ;
        RECT 36.555 160.100 37.690 160.135 ;
        RECT 36.555 160.095 37.720 160.100 ;
        RECT 36.555 159.700 36.785 160.095 ;
        RECT 37.330 160.090 37.720 160.095 ;
        RECT 37.355 160.080 37.720 160.090 ;
        RECT 37.370 160.075 37.720 160.080 ;
        RECT 37.385 160.070 37.720 160.075 ;
        RECT 38.085 160.070 38.345 160.520 ;
        RECT 38.525 160.375 38.855 161.175 ;
        RECT 39.025 160.545 39.255 161.345 ;
        RECT 39.425 160.375 39.755 161.175 ;
        RECT 38.525 160.205 39.755 160.375 ;
        RECT 39.925 160.205 40.180 161.345 ;
        RECT 40.365 160.625 40.695 161.345 ;
        RECT 37.385 160.065 38.345 160.070 ;
        RECT 37.395 160.055 38.345 160.065 ;
        RECT 37.405 160.050 38.345 160.055 ;
        RECT 37.415 160.040 38.345 160.050 ;
        RECT 37.420 160.030 38.345 160.040 ;
        RECT 37.425 160.025 38.345 160.030 ;
        RECT 37.435 160.010 38.345 160.025 ;
        RECT 37.440 159.995 38.345 160.010 ;
        RECT 37.450 159.970 38.345 159.995 ;
        RECT 36.955 159.500 37.285 159.925 ;
        RECT 34.735 158.795 34.950 159.305 ;
        RECT 35.180 158.975 35.460 159.305 ;
        RECT 35.640 158.795 35.880 159.305 ;
        RECT 36.215 158.965 36.475 159.445 ;
        RECT 36.645 158.795 36.895 159.335 ;
        RECT 37.065 159.015 37.285 159.500 ;
        RECT 37.455 159.900 38.345 159.970 ;
        RECT 37.455 159.175 37.625 159.900 ;
        RECT 37.795 159.345 38.345 159.730 ;
        RECT 38.515 159.705 38.825 160.035 ;
        RECT 38.525 159.305 38.855 159.535 ;
        RECT 39.030 159.475 39.405 160.035 ;
        RECT 39.575 159.305 39.755 160.205 ;
        RECT 39.940 159.455 40.160 160.035 ;
        RECT 40.355 159.985 40.585 160.325 ;
        RECT 40.875 159.985 41.090 161.100 ;
        RECT 41.285 160.400 41.615 161.175 ;
        RECT 41.785 160.570 42.495 161.345 ;
        RECT 41.285 160.185 42.435 160.400 ;
        RECT 40.355 159.785 40.685 159.985 ;
        RECT 40.875 159.805 41.325 159.985 ;
        RECT 40.995 159.785 41.325 159.805 ;
        RECT 41.495 159.785 41.965 160.015 ;
        RECT 42.150 159.615 42.435 160.185 ;
        RECT 42.665 159.740 42.945 161.175 ;
        RECT 43.115 160.255 46.625 161.345 ;
        RECT 46.795 160.790 47.400 161.345 ;
        RECT 47.575 160.835 48.055 161.175 ;
        RECT 48.225 160.800 48.480 161.345 ;
        RECT 46.795 160.690 47.410 160.790 ;
        RECT 47.225 160.665 47.410 160.690 ;
        RECT 37.455 159.005 38.345 159.175 ;
        RECT 38.525 158.965 39.755 159.305 ;
        RECT 40.355 159.425 41.535 159.615 ;
        RECT 39.925 158.795 40.180 159.285 ;
        RECT 40.355 158.965 40.695 159.425 ;
        RECT 41.205 159.345 41.535 159.425 ;
        RECT 41.725 159.425 42.435 159.615 ;
        RECT 41.725 159.285 42.025 159.425 ;
        RECT 41.710 159.275 42.025 159.285 ;
        RECT 41.700 159.265 42.025 159.275 ;
        RECT 41.690 159.260 42.025 159.265 ;
        RECT 40.865 158.795 41.035 159.255 ;
        RECT 41.685 159.250 42.025 159.260 ;
        RECT 41.680 159.245 42.025 159.250 ;
        RECT 41.675 159.235 42.025 159.245 ;
        RECT 41.670 159.230 42.025 159.235 ;
        RECT 41.665 158.965 42.025 159.230 ;
        RECT 42.265 158.795 42.435 159.255 ;
        RECT 42.605 158.965 42.945 159.740 ;
        RECT 43.115 159.565 44.765 160.085 ;
        RECT 44.935 159.735 46.625 160.255 ;
        RECT 46.795 160.070 47.055 160.520 ;
        RECT 47.225 160.420 47.555 160.665 ;
        RECT 47.725 160.345 48.480 160.595 ;
        RECT 48.650 160.475 48.925 161.175 ;
        RECT 49.095 160.910 54.440 161.345 ;
        RECT 47.710 160.310 48.480 160.345 ;
        RECT 47.695 160.300 48.480 160.310 ;
        RECT 47.690 160.285 48.585 160.300 ;
        RECT 47.670 160.270 48.585 160.285 ;
        RECT 47.650 160.260 48.585 160.270 ;
        RECT 47.625 160.250 48.585 160.260 ;
        RECT 47.555 160.220 48.585 160.250 ;
        RECT 47.535 160.190 48.585 160.220 ;
        RECT 47.515 160.160 48.585 160.190 ;
        RECT 47.485 160.135 48.585 160.160 ;
        RECT 47.450 160.100 48.585 160.135 ;
        RECT 47.420 160.095 48.585 160.100 ;
        RECT 47.420 160.090 47.810 160.095 ;
        RECT 47.420 160.080 47.785 160.090 ;
        RECT 47.420 160.075 47.770 160.080 ;
        RECT 47.420 160.070 47.755 160.075 ;
        RECT 46.795 160.065 47.755 160.070 ;
        RECT 46.795 160.055 47.745 160.065 ;
        RECT 46.795 160.050 47.735 160.055 ;
        RECT 46.795 160.040 47.725 160.050 ;
        RECT 46.795 160.030 47.720 160.040 ;
        RECT 46.795 160.025 47.715 160.030 ;
        RECT 46.795 160.010 47.705 160.025 ;
        RECT 46.795 159.995 47.700 160.010 ;
        RECT 46.795 159.970 47.690 159.995 ;
        RECT 46.795 159.900 47.685 159.970 ;
        RECT 43.115 158.795 46.625 159.565 ;
        RECT 46.795 159.345 47.345 159.730 ;
        RECT 47.515 159.175 47.685 159.900 ;
        RECT 46.795 159.005 47.685 159.175 ;
        RECT 47.855 159.500 48.185 159.925 ;
        RECT 48.355 159.700 48.585 160.095 ;
        RECT 47.855 159.015 48.075 159.500 ;
        RECT 48.755 159.445 48.925 160.475 ;
        RECT 48.245 158.795 48.495 159.335 ;
        RECT 48.665 158.965 48.925 159.445 ;
        RECT 50.680 159.340 51.020 160.170 ;
        RECT 52.500 159.660 52.850 160.910 ;
        RECT 54.625 160.375 54.955 161.160 ;
        RECT 54.625 160.205 55.305 160.375 ;
        RECT 55.485 160.205 55.815 161.345 ;
        RECT 54.615 159.785 54.965 160.035 ;
        RECT 55.135 159.605 55.305 160.205 ;
        RECT 55.995 160.180 56.285 161.345 ;
        RECT 56.455 160.790 57.060 161.345 ;
        RECT 57.235 160.835 57.715 161.175 ;
        RECT 57.885 160.800 58.140 161.345 ;
        RECT 56.455 160.690 57.070 160.790 ;
        RECT 56.885 160.665 57.070 160.690 ;
        RECT 56.455 160.070 56.715 160.520 ;
        RECT 56.885 160.420 57.215 160.665 ;
        RECT 57.385 160.345 58.140 160.595 ;
        RECT 58.310 160.475 58.585 161.175 ;
        RECT 58.845 160.675 59.015 161.175 ;
        RECT 59.185 160.845 59.515 161.345 ;
        RECT 58.845 160.505 59.510 160.675 ;
        RECT 57.370 160.310 58.140 160.345 ;
        RECT 57.355 160.300 58.140 160.310 ;
        RECT 57.350 160.285 58.245 160.300 ;
        RECT 57.330 160.270 58.245 160.285 ;
        RECT 57.310 160.260 58.245 160.270 ;
        RECT 57.285 160.250 58.245 160.260 ;
        RECT 57.215 160.220 58.245 160.250 ;
        RECT 57.195 160.190 58.245 160.220 ;
        RECT 57.175 160.160 58.245 160.190 ;
        RECT 57.145 160.135 58.245 160.160 ;
        RECT 57.110 160.100 58.245 160.135 ;
        RECT 57.080 160.095 58.245 160.100 ;
        RECT 57.080 160.090 57.470 160.095 ;
        RECT 57.080 160.080 57.445 160.090 ;
        RECT 57.080 160.075 57.430 160.080 ;
        RECT 57.080 160.070 57.415 160.075 ;
        RECT 56.455 160.065 57.415 160.070 ;
        RECT 56.455 160.055 57.405 160.065 ;
        RECT 56.455 160.050 57.395 160.055 ;
        RECT 56.455 160.040 57.385 160.050 ;
        RECT 55.475 159.785 55.825 160.035 ;
        RECT 56.455 160.030 57.380 160.040 ;
        RECT 56.455 160.025 57.375 160.030 ;
        RECT 56.455 160.010 57.365 160.025 ;
        RECT 56.455 159.995 57.360 160.010 ;
        RECT 56.455 159.970 57.350 159.995 ;
        RECT 56.455 159.900 57.345 159.970 ;
        RECT 49.095 158.795 54.440 159.340 ;
        RECT 54.635 158.795 54.875 159.605 ;
        RECT 55.045 158.965 55.375 159.605 ;
        RECT 55.545 158.795 55.815 159.605 ;
        RECT 55.995 158.795 56.285 159.520 ;
        RECT 56.455 159.345 57.005 159.730 ;
        RECT 57.175 159.175 57.345 159.900 ;
        RECT 56.455 159.005 57.345 159.175 ;
        RECT 57.515 159.500 57.845 159.925 ;
        RECT 58.015 159.700 58.245 160.095 ;
        RECT 57.515 159.015 57.735 159.500 ;
        RECT 58.415 159.445 58.585 160.475 ;
        RECT 58.760 159.685 59.110 160.335 ;
        RECT 59.280 159.515 59.510 160.505 ;
        RECT 57.905 158.795 58.155 159.335 ;
        RECT 58.325 158.965 58.585 159.445 ;
        RECT 58.845 159.345 59.510 159.515 ;
        RECT 58.845 159.055 59.015 159.345 ;
        RECT 59.185 158.795 59.515 159.175 ;
        RECT 59.685 159.055 59.870 161.175 ;
        RECT 60.110 160.885 60.375 161.345 ;
        RECT 60.545 160.750 60.795 161.175 ;
        RECT 61.005 160.900 62.110 161.070 ;
        RECT 60.490 160.620 60.795 160.750 ;
        RECT 60.040 159.425 60.320 160.375 ;
        RECT 60.490 159.515 60.660 160.620 ;
        RECT 60.830 159.835 61.070 160.430 ;
        RECT 61.240 160.365 61.770 160.730 ;
        RECT 61.240 159.665 61.410 160.365 ;
        RECT 61.940 160.285 62.110 160.900 ;
        RECT 62.280 160.545 62.450 161.345 ;
        RECT 62.620 160.845 62.870 161.175 ;
        RECT 63.095 160.875 63.980 161.045 ;
        RECT 61.940 160.195 62.450 160.285 ;
        RECT 60.490 159.385 60.715 159.515 ;
        RECT 60.885 159.445 61.410 159.665 ;
        RECT 61.580 160.025 62.450 160.195 ;
        RECT 60.125 158.795 60.375 159.255 ;
        RECT 60.545 159.245 60.715 159.385 ;
        RECT 61.580 159.245 61.750 160.025 ;
        RECT 62.280 159.955 62.450 160.025 ;
        RECT 61.960 159.775 62.160 159.805 ;
        RECT 62.620 159.775 62.790 160.845 ;
        RECT 62.960 159.955 63.150 160.675 ;
        RECT 61.960 159.475 62.790 159.775 ;
        RECT 63.320 159.745 63.640 160.705 ;
        RECT 60.545 159.075 60.880 159.245 ;
        RECT 61.075 159.075 61.750 159.245 ;
        RECT 62.070 158.795 62.440 159.295 ;
        RECT 62.620 159.245 62.790 159.475 ;
        RECT 63.175 159.415 63.640 159.745 ;
        RECT 63.810 160.035 63.980 160.875 ;
        RECT 64.160 160.845 64.475 161.345 ;
        RECT 64.705 160.615 65.045 161.175 ;
        RECT 64.150 160.240 65.045 160.615 ;
        RECT 65.215 160.335 65.385 161.345 ;
        RECT 64.855 160.035 65.045 160.240 ;
        RECT 65.555 160.285 65.885 161.130 ;
        RECT 65.555 160.205 65.945 160.285 ;
        RECT 65.730 160.155 65.945 160.205 ;
        RECT 63.810 159.705 64.685 160.035 ;
        RECT 64.855 159.705 65.605 160.035 ;
        RECT 63.810 159.245 63.980 159.705 ;
        RECT 64.855 159.535 65.055 159.705 ;
        RECT 65.775 159.575 65.945 160.155 ;
        RECT 65.720 159.535 65.945 159.575 ;
        RECT 62.620 159.075 63.025 159.245 ;
        RECT 63.195 159.075 63.980 159.245 ;
        RECT 64.255 158.795 64.465 159.325 ;
        RECT 64.725 159.010 65.055 159.535 ;
        RECT 65.565 159.450 65.945 159.535 ;
        RECT 65.225 158.795 65.395 159.405 ;
        RECT 65.565 159.015 65.895 159.450 ;
        RECT 66.125 158.975 66.385 161.165 ;
        RECT 66.555 160.615 66.895 161.345 ;
        RECT 67.075 160.435 67.345 161.165 ;
        RECT 66.575 160.215 67.345 160.435 ;
        RECT 67.525 160.455 67.755 161.165 ;
        RECT 67.925 160.635 68.255 161.345 ;
        RECT 68.425 160.455 68.685 161.165 ;
        RECT 67.525 160.215 68.685 160.455 ;
        RECT 66.575 159.545 66.865 160.215 ;
        RECT 68.875 160.205 69.135 161.345 ;
        RECT 69.305 160.195 69.635 161.175 ;
        RECT 69.805 160.205 70.085 161.345 ;
        RECT 70.715 160.205 71.100 161.175 ;
        RECT 71.270 160.885 71.595 161.345 ;
        RECT 72.115 160.715 72.395 161.175 ;
        RECT 71.270 160.495 72.395 160.715 ;
        RECT 67.045 159.725 67.510 160.035 ;
        RECT 67.690 159.725 68.215 160.035 ;
        RECT 66.575 159.345 67.805 159.545 ;
        RECT 66.645 158.795 67.315 159.165 ;
        RECT 67.495 158.975 67.805 159.345 ;
        RECT 67.985 159.085 68.215 159.725 ;
        RECT 68.395 159.705 68.695 160.035 ;
        RECT 68.895 159.785 69.230 160.035 ;
        RECT 69.400 159.595 69.570 160.195 ;
        RECT 69.740 159.765 70.075 160.035 ;
        RECT 68.395 158.795 68.685 159.525 ;
        RECT 68.875 158.965 69.570 159.595 ;
        RECT 69.775 158.795 70.085 159.595 ;
        RECT 70.715 159.535 70.995 160.205 ;
        RECT 71.270 160.035 71.720 160.495 ;
        RECT 72.585 160.325 72.985 161.175 ;
        RECT 73.385 160.885 73.655 161.345 ;
        RECT 73.825 160.715 74.110 161.175 ;
        RECT 71.165 159.705 71.720 160.035 ;
        RECT 71.890 159.765 72.985 160.325 ;
        RECT 71.270 159.595 71.720 159.705 ;
        RECT 70.715 158.965 71.100 159.535 ;
        RECT 71.270 159.425 72.395 159.595 ;
        RECT 71.270 158.795 71.595 159.255 ;
        RECT 72.115 158.965 72.395 159.425 ;
        RECT 72.585 158.965 72.985 159.765 ;
        RECT 73.155 160.495 74.110 160.715 ;
        RECT 74.485 160.675 74.655 161.175 ;
        RECT 74.825 160.845 75.155 161.345 ;
        RECT 74.485 160.505 75.150 160.675 ;
        RECT 73.155 159.595 73.365 160.495 ;
        RECT 73.535 159.765 74.225 160.325 ;
        RECT 74.400 159.685 74.750 160.335 ;
        RECT 73.155 159.425 74.110 159.595 ;
        RECT 74.920 159.515 75.150 160.505 ;
        RECT 73.385 158.795 73.655 159.255 ;
        RECT 73.825 158.965 74.110 159.425 ;
        RECT 74.485 159.345 75.150 159.515 ;
        RECT 74.485 159.055 74.655 159.345 ;
        RECT 74.825 158.795 75.155 159.175 ;
        RECT 75.325 159.055 75.510 161.175 ;
        RECT 75.750 160.885 76.015 161.345 ;
        RECT 76.185 160.750 76.435 161.175 ;
        RECT 76.645 160.900 77.750 161.070 ;
        RECT 76.130 160.620 76.435 160.750 ;
        RECT 75.680 159.425 75.960 160.375 ;
        RECT 76.130 159.515 76.300 160.620 ;
        RECT 76.470 159.835 76.710 160.430 ;
        RECT 76.880 160.365 77.410 160.730 ;
        RECT 76.880 159.665 77.050 160.365 ;
        RECT 77.580 160.285 77.750 160.900 ;
        RECT 77.920 160.545 78.090 161.345 ;
        RECT 78.260 160.845 78.510 161.175 ;
        RECT 78.735 160.875 79.620 161.045 ;
        RECT 77.580 160.195 78.090 160.285 ;
        RECT 76.130 159.385 76.355 159.515 ;
        RECT 76.525 159.445 77.050 159.665 ;
        RECT 77.220 160.025 78.090 160.195 ;
        RECT 75.765 158.795 76.015 159.255 ;
        RECT 76.185 159.245 76.355 159.385 ;
        RECT 77.220 159.245 77.390 160.025 ;
        RECT 77.920 159.955 78.090 160.025 ;
        RECT 77.600 159.775 77.800 159.805 ;
        RECT 78.260 159.775 78.430 160.845 ;
        RECT 78.600 159.955 78.790 160.675 ;
        RECT 77.600 159.475 78.430 159.775 ;
        RECT 78.960 159.745 79.280 160.705 ;
        RECT 76.185 159.075 76.520 159.245 ;
        RECT 76.715 159.075 77.390 159.245 ;
        RECT 77.710 158.795 78.080 159.295 ;
        RECT 78.260 159.245 78.430 159.475 ;
        RECT 78.815 159.415 79.280 159.745 ;
        RECT 79.450 160.035 79.620 160.875 ;
        RECT 79.800 160.845 80.115 161.345 ;
        RECT 80.345 160.615 80.685 161.175 ;
        RECT 79.790 160.240 80.685 160.615 ;
        RECT 80.855 160.335 81.025 161.345 ;
        RECT 80.495 160.035 80.685 160.240 ;
        RECT 81.195 160.285 81.525 161.130 ;
        RECT 81.195 160.205 81.585 160.285 ;
        RECT 81.370 160.155 81.585 160.205 ;
        RECT 81.755 160.180 82.045 161.345 ;
        RECT 82.225 160.375 82.555 161.160 ;
        RECT 82.225 160.205 82.905 160.375 ;
        RECT 83.085 160.205 83.415 161.345 ;
        RECT 83.595 160.255 85.265 161.345 ;
        RECT 79.450 159.705 80.325 160.035 ;
        RECT 80.495 159.705 81.245 160.035 ;
        RECT 79.450 159.245 79.620 159.705 ;
        RECT 80.495 159.535 80.695 159.705 ;
        RECT 81.415 159.575 81.585 160.155 ;
        RECT 82.215 159.785 82.565 160.035 ;
        RECT 82.735 159.605 82.905 160.205 ;
        RECT 83.075 159.785 83.425 160.035 ;
        RECT 81.360 159.535 81.585 159.575 ;
        RECT 78.260 159.075 78.665 159.245 ;
        RECT 78.835 159.075 79.620 159.245 ;
        RECT 79.895 158.795 80.105 159.325 ;
        RECT 80.365 159.010 80.695 159.535 ;
        RECT 81.205 159.450 81.585 159.535 ;
        RECT 80.865 158.795 81.035 159.405 ;
        RECT 81.205 159.015 81.535 159.450 ;
        RECT 81.755 158.795 82.045 159.520 ;
        RECT 82.235 158.795 82.475 159.605 ;
        RECT 82.645 158.965 82.975 159.605 ;
        RECT 83.145 158.795 83.415 159.605 ;
        RECT 83.595 159.565 84.345 160.085 ;
        RECT 84.515 159.735 85.265 160.255 ;
        RECT 85.445 160.395 85.720 161.165 ;
        RECT 85.890 160.735 86.220 161.165 ;
        RECT 86.390 160.905 86.585 161.345 ;
        RECT 86.765 160.735 87.095 161.165 ;
        RECT 85.890 160.565 87.095 160.735 ;
        RECT 85.445 160.205 86.030 160.395 ;
        RECT 86.200 160.235 87.095 160.565 ;
        RECT 83.595 158.795 85.265 159.565 ;
        RECT 85.445 159.385 85.685 160.035 ;
        RECT 85.855 159.535 86.030 160.205 ;
        RECT 87.735 160.140 88.025 161.345 ;
        RECT 88.195 160.205 88.470 161.175 ;
        RECT 88.680 160.545 88.960 161.345 ;
        RECT 89.130 160.835 90.325 161.125 ;
        RECT 90.585 160.675 90.755 161.175 ;
        RECT 90.925 160.845 91.255 161.345 ;
        RECT 89.140 160.495 90.305 160.665 ;
        RECT 90.585 160.505 91.250 160.675 ;
        RECT 89.140 160.375 89.310 160.495 ;
        RECT 88.640 160.205 89.310 160.375 ;
        RECT 86.200 159.705 86.615 160.035 ;
        RECT 86.795 159.705 87.090 160.035 ;
        RECT 85.855 159.355 86.185 159.535 ;
        RECT 85.460 158.795 85.790 159.185 ;
        RECT 85.960 158.975 86.185 159.355 ;
        RECT 86.385 159.085 86.615 159.705 ;
        RECT 86.795 158.795 87.095 159.525 ;
        RECT 87.735 158.795 88.025 159.625 ;
        RECT 88.195 159.470 88.365 160.205 ;
        RECT 88.640 160.035 88.810 160.205 ;
        RECT 89.580 160.035 89.805 160.325 ;
        RECT 89.975 160.205 90.305 160.495 ;
        RECT 88.535 159.705 88.810 160.035 ;
        RECT 88.980 159.705 89.805 160.035 ;
        RECT 89.975 159.705 90.325 160.035 ;
        RECT 88.640 159.535 88.810 159.705 ;
        RECT 90.500 159.685 90.850 160.335 ;
        RECT 88.195 159.125 88.470 159.470 ;
        RECT 88.640 159.365 90.305 159.535 ;
        RECT 91.020 159.515 91.250 160.505 ;
        RECT 88.660 158.795 89.040 159.195 ;
        RECT 89.210 159.015 89.380 159.365 ;
        RECT 89.550 158.795 89.880 159.195 ;
        RECT 90.050 159.015 90.305 159.365 ;
        RECT 90.585 159.345 91.250 159.515 ;
        RECT 90.585 159.055 90.755 159.345 ;
        RECT 90.925 158.795 91.255 159.175 ;
        RECT 91.425 159.055 91.610 161.175 ;
        RECT 91.850 160.885 92.115 161.345 ;
        RECT 92.285 160.750 92.535 161.175 ;
        RECT 92.745 160.900 93.850 161.070 ;
        RECT 92.230 160.620 92.535 160.750 ;
        RECT 91.780 159.425 92.060 160.375 ;
        RECT 92.230 159.515 92.400 160.620 ;
        RECT 92.570 159.835 92.810 160.430 ;
        RECT 92.980 160.365 93.510 160.730 ;
        RECT 92.980 159.665 93.150 160.365 ;
        RECT 93.680 160.285 93.850 160.900 ;
        RECT 94.020 160.545 94.190 161.345 ;
        RECT 94.360 160.845 94.610 161.175 ;
        RECT 94.835 160.875 95.720 161.045 ;
        RECT 93.680 160.195 94.190 160.285 ;
        RECT 92.230 159.385 92.455 159.515 ;
        RECT 92.625 159.445 93.150 159.665 ;
        RECT 93.320 160.025 94.190 160.195 ;
        RECT 91.865 158.795 92.115 159.255 ;
        RECT 92.285 159.245 92.455 159.385 ;
        RECT 93.320 159.245 93.490 160.025 ;
        RECT 94.020 159.955 94.190 160.025 ;
        RECT 93.700 159.775 93.900 159.805 ;
        RECT 94.360 159.775 94.530 160.845 ;
        RECT 94.700 159.955 94.890 160.675 ;
        RECT 93.700 159.475 94.530 159.775 ;
        RECT 95.060 159.745 95.380 160.705 ;
        RECT 92.285 159.075 92.620 159.245 ;
        RECT 92.815 159.075 93.490 159.245 ;
        RECT 93.810 158.795 94.180 159.295 ;
        RECT 94.360 159.245 94.530 159.475 ;
        RECT 94.915 159.415 95.380 159.745 ;
        RECT 95.550 160.035 95.720 160.875 ;
        RECT 95.900 160.845 96.215 161.345 ;
        RECT 96.445 160.615 96.785 161.175 ;
        RECT 95.890 160.240 96.785 160.615 ;
        RECT 96.955 160.335 97.125 161.345 ;
        RECT 96.595 160.035 96.785 160.240 ;
        RECT 97.295 160.285 97.625 161.130 ;
        RECT 98.835 160.285 99.165 161.130 ;
        RECT 99.335 160.335 99.505 161.345 ;
        RECT 99.675 160.615 100.015 161.175 ;
        RECT 100.245 160.845 100.560 161.345 ;
        RECT 100.740 160.875 101.625 161.045 ;
        RECT 97.295 160.205 97.685 160.285 ;
        RECT 97.470 160.155 97.685 160.205 ;
        RECT 95.550 159.705 96.425 160.035 ;
        RECT 96.595 159.705 97.345 160.035 ;
        RECT 95.550 159.245 95.720 159.705 ;
        RECT 96.595 159.535 96.795 159.705 ;
        RECT 97.515 159.575 97.685 160.155 ;
        RECT 97.460 159.535 97.685 159.575 ;
        RECT 94.360 159.075 94.765 159.245 ;
        RECT 94.935 159.075 95.720 159.245 ;
        RECT 95.995 158.795 96.205 159.325 ;
        RECT 96.465 159.010 96.795 159.535 ;
        RECT 97.305 159.450 97.685 159.535 ;
        RECT 98.775 160.205 99.165 160.285 ;
        RECT 99.675 160.240 100.570 160.615 ;
        RECT 98.775 160.155 98.990 160.205 ;
        RECT 98.775 159.575 98.945 160.155 ;
        RECT 99.675 160.035 99.865 160.240 ;
        RECT 100.740 160.035 100.910 160.875 ;
        RECT 101.850 160.845 102.100 161.175 ;
        RECT 99.115 159.705 99.865 160.035 ;
        RECT 100.035 159.705 100.910 160.035 ;
        RECT 98.775 159.535 99.000 159.575 ;
        RECT 99.665 159.535 99.865 159.705 ;
        RECT 98.775 159.450 99.155 159.535 ;
        RECT 96.965 158.795 97.135 159.405 ;
        RECT 97.305 159.015 97.635 159.450 ;
        RECT 98.825 159.015 99.155 159.450 ;
        RECT 99.325 158.795 99.495 159.405 ;
        RECT 99.665 159.010 99.995 159.535 ;
        RECT 100.255 158.795 100.465 159.325 ;
        RECT 100.740 159.245 100.910 159.705 ;
        RECT 101.080 159.745 101.400 160.705 ;
        RECT 101.570 159.955 101.760 160.675 ;
        RECT 101.930 159.775 102.100 160.845 ;
        RECT 102.270 160.545 102.440 161.345 ;
        RECT 102.610 160.900 103.715 161.070 ;
        RECT 102.610 160.285 102.780 160.900 ;
        RECT 103.925 160.750 104.175 161.175 ;
        RECT 104.345 160.885 104.610 161.345 ;
        RECT 102.950 160.365 103.480 160.730 ;
        RECT 103.925 160.620 104.230 160.750 ;
        RECT 102.270 160.195 102.780 160.285 ;
        RECT 102.270 160.025 103.140 160.195 ;
        RECT 102.270 159.955 102.440 160.025 ;
        RECT 102.560 159.775 102.760 159.805 ;
        RECT 101.080 159.415 101.545 159.745 ;
        RECT 101.930 159.475 102.760 159.775 ;
        RECT 101.930 159.245 102.100 159.475 ;
        RECT 100.740 159.075 101.525 159.245 ;
        RECT 101.695 159.075 102.100 159.245 ;
        RECT 102.280 158.795 102.650 159.295 ;
        RECT 102.970 159.245 103.140 160.025 ;
        RECT 103.310 159.665 103.480 160.365 ;
        RECT 103.650 159.835 103.890 160.430 ;
        RECT 103.310 159.445 103.835 159.665 ;
        RECT 104.060 159.515 104.230 160.620 ;
        RECT 104.005 159.385 104.230 159.515 ;
        RECT 104.400 159.425 104.680 160.375 ;
        RECT 104.005 159.245 104.175 159.385 ;
        RECT 102.970 159.075 103.645 159.245 ;
        RECT 103.840 159.075 104.175 159.245 ;
        RECT 104.345 158.795 104.595 159.255 ;
        RECT 104.850 159.055 105.035 161.175 ;
        RECT 105.205 160.845 105.535 161.345 ;
        RECT 105.705 160.675 105.875 161.175 ;
        RECT 105.210 160.505 105.875 160.675 ;
        RECT 105.210 159.515 105.440 160.505 ;
        RECT 105.610 159.685 105.960 160.335 ;
        RECT 106.135 160.255 107.345 161.345 ;
        RECT 106.135 159.545 106.655 160.085 ;
        RECT 106.825 159.715 107.345 160.255 ;
        RECT 107.515 160.180 107.805 161.345 ;
        RECT 107.980 160.205 108.315 161.175 ;
        RECT 108.485 160.205 108.655 161.345 ;
        RECT 108.825 161.005 110.855 161.175 ;
        RECT 105.210 159.345 105.875 159.515 ;
        RECT 105.205 158.795 105.535 159.175 ;
        RECT 105.705 159.055 105.875 159.345 ;
        RECT 106.135 158.795 107.345 159.545 ;
        RECT 107.980 159.535 108.150 160.205 ;
        RECT 108.825 160.035 108.995 161.005 ;
        RECT 108.320 159.705 108.575 160.035 ;
        RECT 108.800 159.705 108.995 160.035 ;
        RECT 109.165 160.665 110.290 160.835 ;
        RECT 108.405 159.535 108.575 159.705 ;
        RECT 109.165 159.535 109.335 160.665 ;
        RECT 107.515 158.795 107.805 159.520 ;
        RECT 107.980 158.965 108.235 159.535 ;
        RECT 108.405 159.365 109.335 159.535 ;
        RECT 109.505 160.325 110.515 160.495 ;
        RECT 109.505 159.525 109.675 160.325 ;
        RECT 109.880 159.985 110.155 160.125 ;
        RECT 109.875 159.815 110.155 159.985 ;
        RECT 109.160 159.330 109.335 159.365 ;
        RECT 108.405 158.795 108.735 159.195 ;
        RECT 109.160 158.965 109.690 159.330 ;
        RECT 109.880 158.965 110.155 159.815 ;
        RECT 110.325 158.965 110.515 160.325 ;
        RECT 110.685 160.340 110.855 161.005 ;
        RECT 111.025 160.585 111.195 161.345 ;
        RECT 111.430 160.585 111.945 160.995 ;
        RECT 110.685 160.150 111.435 160.340 ;
        RECT 111.605 159.775 111.945 160.585 ;
        RECT 112.125 160.375 112.455 161.160 ;
        RECT 112.125 160.205 112.805 160.375 ;
        RECT 112.985 160.205 113.315 161.345 ;
        RECT 113.495 160.910 118.840 161.345 ;
        RECT 112.115 159.785 112.465 160.035 ;
        RECT 110.715 159.605 111.945 159.775 ;
        RECT 112.635 159.605 112.805 160.205 ;
        RECT 112.975 159.785 113.325 160.035 ;
        RECT 110.695 158.795 111.205 159.330 ;
        RECT 111.425 159.000 111.670 159.605 ;
        RECT 112.135 158.795 112.375 159.605 ;
        RECT 112.545 158.965 112.875 159.605 ;
        RECT 113.045 158.795 113.315 159.605 ;
        RECT 115.080 159.340 115.420 160.170 ;
        RECT 116.900 159.660 117.250 160.910 ;
        RECT 119.015 160.205 119.295 161.345 ;
        RECT 119.465 160.195 119.795 161.175 ;
        RECT 119.965 160.205 120.225 161.345 ;
        RECT 120.395 160.255 122.065 161.345 ;
        RECT 119.025 159.765 119.360 160.035 ;
        RECT 119.530 159.595 119.700 160.195 ;
        RECT 119.870 159.785 120.205 160.035 ;
        RECT 113.495 158.795 118.840 159.340 ;
        RECT 119.015 158.795 119.325 159.595 ;
        RECT 119.530 158.965 120.225 159.595 ;
        RECT 120.395 159.565 121.145 160.085 ;
        RECT 121.315 159.735 122.065 160.255 ;
        RECT 122.735 160.205 122.965 161.345 ;
        RECT 123.135 160.195 123.465 161.175 ;
        RECT 123.635 160.205 123.845 161.345 ;
        RECT 125.295 160.705 125.625 161.135 ;
        RECT 125.170 160.535 125.625 160.705 ;
        RECT 125.805 160.705 126.055 161.125 ;
        RECT 126.285 160.875 126.615 161.345 ;
        RECT 126.845 160.705 127.095 161.125 ;
        RECT 125.805 160.535 127.095 160.705 ;
        RECT 122.715 159.785 123.045 160.035 ;
        RECT 120.395 158.795 122.065 159.565 ;
        RECT 122.735 158.795 122.965 159.615 ;
        RECT 123.215 159.595 123.465 160.195 ;
        RECT 123.135 158.965 123.465 159.595 ;
        RECT 123.635 158.795 123.845 159.615 ;
        RECT 125.170 159.535 125.340 160.535 ;
        RECT 125.510 159.705 125.755 160.365 ;
        RECT 125.970 159.705 126.235 160.365 ;
        RECT 126.430 159.705 126.715 160.365 ;
        RECT 126.890 160.035 127.105 160.365 ;
        RECT 127.285 160.205 127.535 161.345 ;
        RECT 127.705 160.285 128.035 161.135 ;
        RECT 126.890 159.705 127.195 160.035 ;
        RECT 127.365 159.705 127.675 160.035 ;
        RECT 127.365 159.535 127.535 159.705 ;
        RECT 125.170 159.365 127.535 159.535 ;
        RECT 127.845 159.520 128.035 160.285 ;
        RECT 128.215 160.205 128.475 161.345 ;
        RECT 128.645 160.195 128.975 161.175 ;
        RECT 129.145 160.205 129.425 161.345 ;
        RECT 129.595 160.255 133.105 161.345 ;
        RECT 128.235 159.785 128.570 160.035 ;
        RECT 128.740 159.645 128.910 160.195 ;
        RECT 129.080 159.765 129.415 160.035 ;
        RECT 128.735 159.595 128.910 159.645 ;
        RECT 125.325 158.795 125.655 159.195 ;
        RECT 125.825 159.025 126.155 159.365 ;
        RECT 127.205 158.795 127.535 159.195 ;
        RECT 127.705 159.010 128.035 159.520 ;
        RECT 128.215 158.965 128.910 159.595 ;
        RECT 129.115 158.795 129.425 159.595 ;
        RECT 129.595 159.565 131.245 160.085 ;
        RECT 131.415 159.735 133.105 160.255 ;
        RECT 133.275 160.180 133.565 161.345 ;
        RECT 133.825 160.675 133.995 161.175 ;
        RECT 134.165 160.845 134.495 161.345 ;
        RECT 133.825 160.505 134.490 160.675 ;
        RECT 133.740 159.685 134.090 160.335 ;
        RECT 129.595 158.795 133.105 159.565 ;
        RECT 133.275 158.795 133.565 159.520 ;
        RECT 134.260 159.515 134.490 160.505 ;
        RECT 133.825 159.345 134.490 159.515 ;
        RECT 133.825 159.055 133.995 159.345 ;
        RECT 134.165 158.795 134.495 159.175 ;
        RECT 134.665 159.055 134.850 161.175 ;
        RECT 135.090 160.885 135.355 161.345 ;
        RECT 135.525 160.750 135.775 161.175 ;
        RECT 135.985 160.900 137.090 161.070 ;
        RECT 135.470 160.620 135.775 160.750 ;
        RECT 135.020 159.425 135.300 160.375 ;
        RECT 135.470 159.515 135.640 160.620 ;
        RECT 135.810 159.835 136.050 160.430 ;
        RECT 136.220 160.365 136.750 160.730 ;
        RECT 136.220 159.665 136.390 160.365 ;
        RECT 136.920 160.285 137.090 160.900 ;
        RECT 137.260 160.545 137.430 161.345 ;
        RECT 137.600 160.845 137.850 161.175 ;
        RECT 138.075 160.875 138.960 161.045 ;
        RECT 136.920 160.195 137.430 160.285 ;
        RECT 135.470 159.385 135.695 159.515 ;
        RECT 135.865 159.445 136.390 159.665 ;
        RECT 136.560 160.025 137.430 160.195 ;
        RECT 135.105 158.795 135.355 159.255 ;
        RECT 135.525 159.245 135.695 159.385 ;
        RECT 136.560 159.245 136.730 160.025 ;
        RECT 137.260 159.955 137.430 160.025 ;
        RECT 136.940 159.775 137.140 159.805 ;
        RECT 137.600 159.775 137.770 160.845 ;
        RECT 137.940 159.955 138.130 160.675 ;
        RECT 136.940 159.475 137.770 159.775 ;
        RECT 138.300 159.745 138.620 160.705 ;
        RECT 135.525 159.075 135.860 159.245 ;
        RECT 136.055 159.075 136.730 159.245 ;
        RECT 137.050 158.795 137.420 159.295 ;
        RECT 137.600 159.245 137.770 159.475 ;
        RECT 138.155 159.415 138.620 159.745 ;
        RECT 138.790 160.035 138.960 160.875 ;
        RECT 139.140 160.845 139.455 161.345 ;
        RECT 139.685 160.615 140.025 161.175 ;
        RECT 139.130 160.240 140.025 160.615 ;
        RECT 140.195 160.335 140.365 161.345 ;
        RECT 139.835 160.035 140.025 160.240 ;
        RECT 140.535 160.285 140.865 161.130 ;
        RECT 140.535 160.205 140.925 160.285 ;
        RECT 140.710 160.155 140.925 160.205 ;
        RECT 138.790 159.705 139.665 160.035 ;
        RECT 139.835 159.705 140.585 160.035 ;
        RECT 138.790 159.245 138.960 159.705 ;
        RECT 139.835 159.535 140.035 159.705 ;
        RECT 140.755 159.575 140.925 160.155 ;
        RECT 140.700 159.535 140.925 159.575 ;
        RECT 137.600 159.075 138.005 159.245 ;
        RECT 138.175 159.075 138.960 159.245 ;
        RECT 139.235 158.795 139.445 159.325 ;
        RECT 139.705 159.010 140.035 159.535 ;
        RECT 140.545 159.450 140.925 159.535 ;
        RECT 141.100 160.205 141.435 161.175 ;
        RECT 141.605 160.205 141.775 161.345 ;
        RECT 141.945 161.005 143.975 161.175 ;
        RECT 141.100 159.535 141.270 160.205 ;
        RECT 141.945 160.035 142.115 161.005 ;
        RECT 141.440 159.705 141.695 160.035 ;
        RECT 141.920 159.705 142.115 160.035 ;
        RECT 142.285 160.665 143.410 160.835 ;
        RECT 141.525 159.535 141.695 159.705 ;
        RECT 142.285 159.535 142.455 160.665 ;
        RECT 140.205 158.795 140.375 159.405 ;
        RECT 140.545 159.015 140.875 159.450 ;
        RECT 141.100 158.965 141.355 159.535 ;
        RECT 141.525 159.365 142.455 159.535 ;
        RECT 142.625 160.325 143.635 160.495 ;
        RECT 142.625 159.525 142.795 160.325 ;
        RECT 142.280 159.330 142.455 159.365 ;
        RECT 141.525 158.795 141.855 159.195 ;
        RECT 142.280 158.965 142.810 159.330 ;
        RECT 143.000 159.305 143.275 160.125 ;
        RECT 142.995 159.135 143.275 159.305 ;
        RECT 143.000 158.965 143.275 159.135 ;
        RECT 143.445 158.965 143.635 160.325 ;
        RECT 143.805 160.340 143.975 161.005 ;
        RECT 144.145 160.585 144.315 161.345 ;
        RECT 144.550 160.585 145.065 160.995 ;
        RECT 143.805 160.150 144.555 160.340 ;
        RECT 144.725 159.775 145.065 160.585 ;
        RECT 143.835 159.605 145.065 159.775 ;
        RECT 145.695 160.255 146.905 161.345 ;
        RECT 145.695 159.715 146.215 160.255 ;
        RECT 143.815 158.795 144.325 159.330 ;
        RECT 144.545 159.000 144.790 159.605 ;
        RECT 146.385 159.545 146.905 160.085 ;
        RECT 145.695 158.795 146.905 159.545 ;
        RECT 17.270 158.625 146.990 158.795 ;
        RECT 17.355 157.875 18.565 158.625 ;
        RECT 18.735 158.080 24.080 158.625 ;
        RECT 24.255 158.080 29.600 158.625 ;
        RECT 17.355 157.335 17.875 157.875 ;
        RECT 18.045 157.165 18.565 157.705 ;
        RECT 20.320 157.250 20.660 158.080 ;
        RECT 17.355 156.075 18.565 157.165 ;
        RECT 22.140 156.510 22.490 157.760 ;
        RECT 25.840 157.250 26.180 158.080 ;
        RECT 30.695 157.825 31.390 158.455 ;
        RECT 31.595 157.825 31.905 158.625 ;
        RECT 32.075 158.245 32.965 158.415 ;
        RECT 31.215 157.775 31.390 157.825 ;
        RECT 27.660 156.510 28.010 157.760 ;
        RECT 30.715 157.385 31.050 157.635 ;
        RECT 31.220 157.225 31.390 157.775 ;
        RECT 32.075 157.690 32.625 158.075 ;
        RECT 31.560 157.385 31.895 157.655 ;
        RECT 32.795 157.520 32.965 158.245 ;
        RECT 32.075 157.450 32.965 157.520 ;
        RECT 33.135 157.945 33.355 158.405 ;
        RECT 33.525 158.085 33.775 158.625 ;
        RECT 33.945 157.975 34.205 158.455 ;
        RECT 33.135 157.920 33.385 157.945 ;
        RECT 33.135 157.495 33.465 157.920 ;
        RECT 32.075 157.425 32.970 157.450 ;
        RECT 32.075 157.410 32.980 157.425 ;
        RECT 32.075 157.395 32.985 157.410 ;
        RECT 32.075 157.390 32.995 157.395 ;
        RECT 32.075 157.380 33.000 157.390 ;
        RECT 32.075 157.370 33.005 157.380 ;
        RECT 32.075 157.365 33.015 157.370 ;
        RECT 32.075 157.355 33.025 157.365 ;
        RECT 32.075 157.350 33.035 157.355 ;
        RECT 18.735 156.075 24.080 156.510 ;
        RECT 24.255 156.075 29.600 156.510 ;
        RECT 30.695 156.075 30.955 157.215 ;
        RECT 31.125 156.245 31.455 157.225 ;
        RECT 31.625 156.075 31.905 157.215 ;
        RECT 32.075 156.900 32.335 157.350 ;
        RECT 32.700 157.345 33.035 157.350 ;
        RECT 32.700 157.340 33.050 157.345 ;
        RECT 32.700 157.330 33.065 157.340 ;
        RECT 32.700 157.325 33.090 157.330 ;
        RECT 33.635 157.325 33.865 157.720 ;
        RECT 32.700 157.320 33.865 157.325 ;
        RECT 32.730 157.285 33.865 157.320 ;
        RECT 32.765 157.260 33.865 157.285 ;
        RECT 32.795 157.230 33.865 157.260 ;
        RECT 32.815 157.200 33.865 157.230 ;
        RECT 32.835 157.170 33.865 157.200 ;
        RECT 32.905 157.160 33.865 157.170 ;
        RECT 32.930 157.150 33.865 157.160 ;
        RECT 32.950 157.135 33.865 157.150 ;
        RECT 32.970 157.120 33.865 157.135 ;
        RECT 32.975 157.110 33.760 157.120 ;
        RECT 32.990 157.075 33.760 157.110 ;
        RECT 32.505 156.755 32.835 157.000 ;
        RECT 33.005 156.825 33.760 157.075 ;
        RECT 34.035 156.945 34.205 157.975 ;
        RECT 34.465 158.075 34.635 158.365 ;
        RECT 34.805 158.245 35.135 158.625 ;
        RECT 34.465 157.905 35.130 158.075 ;
        RECT 34.380 157.085 34.730 157.735 ;
        RECT 32.505 156.730 32.690 156.755 ;
        RECT 32.075 156.630 32.690 156.730 ;
        RECT 32.075 156.075 32.680 156.630 ;
        RECT 32.855 156.245 33.335 156.585 ;
        RECT 33.505 156.075 33.760 156.620 ;
        RECT 33.930 156.245 34.205 156.945 ;
        RECT 34.900 156.915 35.130 157.905 ;
        RECT 34.465 156.745 35.130 156.915 ;
        RECT 34.465 156.245 34.635 156.745 ;
        RECT 34.805 156.075 35.135 156.575 ;
        RECT 35.305 156.245 35.490 158.365 ;
        RECT 35.745 158.165 35.995 158.625 ;
        RECT 36.165 158.175 36.500 158.345 ;
        RECT 36.695 158.175 37.370 158.345 ;
        RECT 36.165 158.035 36.335 158.175 ;
        RECT 35.660 157.045 35.940 157.995 ;
        RECT 36.110 157.905 36.335 158.035 ;
        RECT 36.110 156.800 36.280 157.905 ;
        RECT 36.505 157.755 37.030 157.975 ;
        RECT 36.450 156.990 36.690 157.585 ;
        RECT 36.860 157.055 37.030 157.755 ;
        RECT 37.200 157.395 37.370 158.175 ;
        RECT 37.690 158.125 38.060 158.625 ;
        RECT 38.240 158.175 38.645 158.345 ;
        RECT 38.815 158.175 39.600 158.345 ;
        RECT 38.240 157.945 38.410 158.175 ;
        RECT 37.580 157.645 38.410 157.945 ;
        RECT 38.795 157.675 39.260 158.005 ;
        RECT 37.580 157.615 37.780 157.645 ;
        RECT 37.900 157.395 38.070 157.465 ;
        RECT 37.200 157.225 38.070 157.395 ;
        RECT 37.560 157.135 38.070 157.225 ;
        RECT 36.110 156.670 36.415 156.800 ;
        RECT 36.860 156.690 37.390 157.055 ;
        RECT 35.730 156.075 35.995 156.535 ;
        RECT 36.165 156.245 36.415 156.670 ;
        RECT 37.560 156.520 37.730 157.135 ;
        RECT 36.625 156.350 37.730 156.520 ;
        RECT 37.900 156.075 38.070 156.875 ;
        RECT 38.240 156.575 38.410 157.645 ;
        RECT 38.580 156.745 38.770 157.465 ;
        RECT 38.940 156.715 39.260 157.675 ;
        RECT 39.430 157.715 39.600 158.175 ;
        RECT 39.875 158.095 40.085 158.625 ;
        RECT 40.345 157.885 40.675 158.410 ;
        RECT 40.845 158.015 41.015 158.625 ;
        RECT 41.185 157.970 41.515 158.405 ;
        RECT 41.185 157.885 41.565 157.970 ;
        RECT 40.475 157.715 40.675 157.885 ;
        RECT 41.340 157.845 41.565 157.885 ;
        RECT 39.430 157.385 40.305 157.715 ;
        RECT 40.475 157.385 41.225 157.715 ;
        RECT 38.240 156.245 38.490 156.575 ;
        RECT 39.430 156.545 39.600 157.385 ;
        RECT 40.475 157.180 40.665 157.385 ;
        RECT 41.395 157.265 41.565 157.845 ;
        RECT 41.735 157.875 42.945 158.625 ;
        RECT 43.115 157.900 43.405 158.625 ;
        RECT 41.735 157.335 42.255 157.875 ;
        RECT 43.575 157.855 45.245 158.625 ;
        RECT 41.350 157.215 41.565 157.265 ;
        RECT 39.770 156.805 40.665 157.180 ;
        RECT 41.175 157.135 41.565 157.215 ;
        RECT 42.425 157.165 42.945 157.705 ;
        RECT 43.575 157.335 44.325 157.855 ;
        RECT 38.715 156.375 39.600 156.545 ;
        RECT 39.780 156.075 40.095 156.575 ;
        RECT 40.325 156.245 40.665 156.805 ;
        RECT 40.835 156.075 41.005 157.085 ;
        RECT 41.175 156.290 41.505 157.135 ;
        RECT 41.735 156.075 42.945 157.165 ;
        RECT 43.115 156.075 43.405 157.240 ;
        RECT 44.495 157.165 45.245 157.685 ;
        RECT 43.575 156.075 45.245 157.165 ;
        RECT 45.415 156.245 45.695 158.345 ;
        RECT 45.925 158.165 46.095 158.625 ;
        RECT 46.365 158.235 47.615 158.415 ;
        RECT 46.750 157.995 47.115 158.065 ;
        RECT 45.865 157.815 47.115 157.995 ;
        RECT 47.285 158.015 47.615 158.235 ;
        RECT 47.785 158.185 47.955 158.625 ;
        RECT 48.125 158.015 48.465 158.430 ;
        RECT 47.285 157.845 48.465 158.015 ;
        RECT 48.635 157.875 49.845 158.625 ;
        RECT 50.105 157.975 50.275 158.455 ;
        RECT 50.445 158.145 50.775 158.625 ;
        RECT 51.000 158.205 52.535 158.455 ;
        RECT 51.000 157.975 51.170 158.205 ;
        RECT 45.865 157.215 46.140 157.815 ;
        RECT 46.310 157.385 46.665 157.635 ;
        RECT 46.860 157.605 47.325 157.635 ;
        RECT 46.855 157.435 47.325 157.605 ;
        RECT 46.860 157.385 47.325 157.435 ;
        RECT 47.495 157.385 47.825 157.635 ;
        RECT 48.000 157.435 48.465 157.635 ;
        RECT 47.645 157.265 47.825 157.385 ;
        RECT 48.635 157.335 49.155 157.875 ;
        RECT 50.105 157.805 51.170 157.975 ;
        RECT 45.865 157.005 47.475 157.215 ;
        RECT 47.645 157.095 47.975 157.265 ;
        RECT 47.065 156.905 47.475 157.005 ;
        RECT 45.885 156.075 46.670 156.835 ;
        RECT 47.065 156.245 47.450 156.905 ;
        RECT 47.775 156.305 47.975 157.095 ;
        RECT 48.145 156.075 48.465 157.255 ;
        RECT 49.325 157.165 49.845 157.705 ;
        RECT 51.350 157.635 51.630 158.035 ;
        RECT 50.020 157.425 50.370 157.635 ;
        RECT 50.540 157.435 50.985 157.635 ;
        RECT 51.155 157.435 51.630 157.635 ;
        RECT 51.900 157.635 52.185 158.035 ;
        RECT 52.365 157.975 52.535 158.205 ;
        RECT 52.705 158.145 53.035 158.625 ;
        RECT 53.250 158.125 53.505 158.455 ;
        RECT 53.320 158.045 53.505 158.125 ;
        RECT 52.365 157.805 53.165 157.975 ;
        RECT 51.900 157.435 52.230 157.635 ;
        RECT 52.400 157.435 52.765 157.635 ;
        RECT 52.995 157.255 53.165 157.805 ;
        RECT 48.635 156.075 49.845 157.165 ;
        RECT 50.105 157.085 53.165 157.255 ;
        RECT 50.105 156.245 50.275 157.085 ;
        RECT 53.335 156.925 53.505 158.045 ;
        RECT 53.705 157.895 54.005 158.625 ;
        RECT 54.185 157.715 54.415 158.335 ;
        RECT 54.615 158.065 54.840 158.445 ;
        RECT 55.010 158.235 55.340 158.625 ;
        RECT 54.615 157.885 54.945 158.065 ;
        RECT 53.710 157.385 54.005 157.715 ;
        RECT 54.185 157.385 54.600 157.715 ;
        RECT 54.770 157.215 54.945 157.885 ;
        RECT 55.115 157.385 55.355 158.035 ;
        RECT 56.545 157.975 56.715 158.455 ;
        RECT 56.885 158.145 57.215 158.625 ;
        RECT 57.440 158.205 58.975 158.455 ;
        RECT 57.440 157.975 57.610 158.205 ;
        RECT 56.545 157.805 57.610 157.975 ;
        RECT 57.790 157.635 58.070 158.035 ;
        RECT 56.460 157.425 56.810 157.635 ;
        RECT 56.980 157.435 57.425 157.635 ;
        RECT 57.595 157.435 58.070 157.635 ;
        RECT 58.340 157.635 58.625 158.035 ;
        RECT 58.805 157.975 58.975 158.205 ;
        RECT 59.145 158.145 59.475 158.625 ;
        RECT 59.690 158.125 59.945 158.455 ;
        RECT 59.760 158.045 59.945 158.125 ;
        RECT 58.805 157.805 59.605 157.975 ;
        RECT 58.340 157.435 58.670 157.635 ;
        RECT 58.840 157.605 59.205 157.635 ;
        RECT 58.840 157.435 59.215 157.605 ;
        RECT 59.435 157.255 59.605 157.805 ;
        RECT 53.295 156.915 53.505 156.925 ;
        RECT 50.445 156.415 50.775 156.915 ;
        RECT 50.945 156.675 52.580 156.915 ;
        RECT 50.945 156.585 51.175 156.675 ;
        RECT 51.285 156.415 51.615 156.455 ;
        RECT 50.445 156.245 51.615 156.415 ;
        RECT 51.805 156.075 52.160 156.495 ;
        RECT 52.330 156.245 52.580 156.675 ;
        RECT 52.750 156.075 53.080 156.835 ;
        RECT 53.250 156.245 53.505 156.915 ;
        RECT 53.705 156.855 54.600 157.185 ;
        RECT 54.770 157.025 55.355 157.215 ;
        RECT 53.705 156.685 54.910 156.855 ;
        RECT 53.705 156.255 54.035 156.685 ;
        RECT 54.215 156.075 54.410 156.515 ;
        RECT 54.580 156.255 54.910 156.685 ;
        RECT 55.080 156.255 55.355 157.025 ;
        RECT 56.545 157.085 59.605 157.255 ;
        RECT 56.545 156.245 56.715 157.085 ;
        RECT 59.775 156.925 59.945 158.045 ;
        RECT 61.060 157.860 61.515 158.625 ;
        RECT 61.790 158.245 63.090 158.455 ;
        RECT 63.345 158.265 63.675 158.625 ;
        RECT 62.920 158.095 63.090 158.245 ;
        RECT 63.845 158.125 64.105 158.455 ;
        RECT 61.990 157.635 62.210 158.035 ;
        RECT 61.055 157.435 61.545 157.635 ;
        RECT 61.735 157.425 62.210 157.635 ;
        RECT 62.455 157.635 62.665 158.035 ;
        RECT 62.920 157.970 63.675 158.095 ;
        RECT 62.920 157.925 63.765 157.970 ;
        RECT 63.495 157.805 63.765 157.925 ;
        RECT 62.455 157.425 62.785 157.635 ;
        RECT 62.955 157.365 63.365 157.670 ;
        RECT 59.735 156.915 59.945 156.925 ;
        RECT 56.885 156.415 57.215 156.915 ;
        RECT 57.385 156.675 59.020 156.915 ;
        RECT 57.385 156.585 57.615 156.675 ;
        RECT 57.725 156.415 58.055 156.455 ;
        RECT 56.885 156.245 58.055 156.415 ;
        RECT 58.245 156.075 58.600 156.495 ;
        RECT 58.770 156.245 59.020 156.675 ;
        RECT 59.190 156.075 59.520 156.835 ;
        RECT 59.690 156.245 59.945 156.915 ;
        RECT 61.060 157.195 62.235 157.255 ;
        RECT 63.595 157.230 63.765 157.805 ;
        RECT 63.565 157.195 63.765 157.230 ;
        RECT 61.060 157.085 63.765 157.195 ;
        RECT 61.060 156.465 61.315 157.085 ;
        RECT 61.905 157.025 63.705 157.085 ;
        RECT 61.905 156.995 62.235 157.025 ;
        RECT 63.935 156.925 64.105 158.125 ;
        RECT 61.565 156.825 61.750 156.915 ;
        RECT 62.340 156.825 63.175 156.835 ;
        RECT 61.565 156.625 63.175 156.825 ;
        RECT 61.565 156.585 61.795 156.625 ;
        RECT 61.060 156.245 61.395 156.465 ;
        RECT 62.400 156.075 62.755 156.455 ;
        RECT 62.925 156.245 63.175 156.625 ;
        RECT 63.425 156.075 63.675 156.855 ;
        RECT 63.845 156.245 64.105 156.925 ;
        RECT 64.310 157.885 64.925 158.455 ;
        RECT 65.095 158.115 65.310 158.625 ;
        RECT 65.540 158.115 65.820 158.445 ;
        RECT 66.000 158.115 66.240 158.625 ;
        RECT 64.310 156.865 64.625 157.885 ;
        RECT 64.795 157.215 64.965 157.715 ;
        RECT 65.215 157.385 65.480 157.945 ;
        RECT 65.650 157.215 65.820 158.115 ;
        RECT 65.990 157.385 66.345 157.945 ;
        RECT 66.575 157.855 68.245 158.625 ;
        RECT 68.875 157.900 69.165 158.625 ;
        RECT 69.885 158.075 70.055 158.365 ;
        RECT 70.225 158.245 70.555 158.625 ;
        RECT 69.885 157.905 70.550 158.075 ;
        RECT 66.575 157.335 67.325 157.855 ;
        RECT 64.795 157.045 66.220 157.215 ;
        RECT 67.495 157.165 68.245 157.685 ;
        RECT 64.310 156.245 64.845 156.865 ;
        RECT 65.015 156.075 65.345 156.875 ;
        RECT 65.830 156.870 66.220 157.045 ;
        RECT 66.575 156.075 68.245 157.165 ;
        RECT 68.875 156.075 69.165 157.240 ;
        RECT 69.800 157.085 70.150 157.735 ;
        RECT 70.320 156.915 70.550 157.905 ;
        RECT 69.885 156.745 70.550 156.915 ;
        RECT 69.885 156.245 70.055 156.745 ;
        RECT 70.225 156.075 70.555 156.575 ;
        RECT 70.725 156.245 70.910 158.365 ;
        RECT 71.165 158.165 71.415 158.625 ;
        RECT 71.585 158.175 71.920 158.345 ;
        RECT 72.115 158.175 72.790 158.345 ;
        RECT 71.585 158.035 71.755 158.175 ;
        RECT 71.080 157.045 71.360 157.995 ;
        RECT 71.530 157.905 71.755 158.035 ;
        RECT 71.530 156.800 71.700 157.905 ;
        RECT 71.925 157.755 72.450 157.975 ;
        RECT 71.870 156.990 72.110 157.585 ;
        RECT 72.280 157.055 72.450 157.755 ;
        RECT 72.620 157.395 72.790 158.175 ;
        RECT 73.110 158.125 73.480 158.625 ;
        RECT 73.660 158.175 74.065 158.345 ;
        RECT 74.235 158.175 75.020 158.345 ;
        RECT 73.660 157.945 73.830 158.175 ;
        RECT 73.000 157.645 73.830 157.945 ;
        RECT 74.215 157.675 74.680 158.005 ;
        RECT 73.000 157.615 73.200 157.645 ;
        RECT 73.320 157.395 73.490 157.465 ;
        RECT 72.620 157.225 73.490 157.395 ;
        RECT 72.980 157.135 73.490 157.225 ;
        RECT 71.530 156.670 71.835 156.800 ;
        RECT 72.280 156.690 72.810 157.055 ;
        RECT 71.150 156.075 71.415 156.535 ;
        RECT 71.585 156.245 71.835 156.670 ;
        RECT 72.980 156.520 73.150 157.135 ;
        RECT 72.045 156.350 73.150 156.520 ;
        RECT 73.320 156.075 73.490 156.875 ;
        RECT 73.660 156.575 73.830 157.645 ;
        RECT 74.000 156.745 74.190 157.465 ;
        RECT 74.360 156.715 74.680 157.675 ;
        RECT 74.850 157.715 75.020 158.175 ;
        RECT 75.295 158.095 75.505 158.625 ;
        RECT 75.765 157.885 76.095 158.410 ;
        RECT 76.265 158.015 76.435 158.625 ;
        RECT 76.605 157.970 76.935 158.405 ;
        RECT 76.605 157.885 76.985 157.970 ;
        RECT 75.895 157.715 76.095 157.885 ;
        RECT 76.760 157.845 76.985 157.885 ;
        RECT 74.850 157.385 75.725 157.715 ;
        RECT 75.895 157.385 76.645 157.715 ;
        RECT 73.660 156.245 73.910 156.575 ;
        RECT 74.850 156.545 75.020 157.385 ;
        RECT 75.895 157.180 76.085 157.385 ;
        RECT 76.815 157.265 76.985 157.845 ;
        RECT 77.155 157.855 79.745 158.625 ;
        RECT 80.375 158.115 80.680 158.625 ;
        RECT 77.155 157.335 78.365 157.855 ;
        RECT 76.770 157.215 76.985 157.265 ;
        RECT 75.190 156.805 76.085 157.180 ;
        RECT 76.595 157.135 76.985 157.215 ;
        RECT 78.535 157.165 79.745 157.685 ;
        RECT 80.375 157.385 80.690 157.945 ;
        RECT 80.860 157.635 81.110 158.445 ;
        RECT 81.280 158.100 81.540 158.625 ;
        RECT 81.720 157.635 81.970 158.445 ;
        RECT 82.140 158.065 82.400 158.625 ;
        RECT 82.570 157.975 82.830 158.430 ;
        RECT 83.000 158.145 83.260 158.625 ;
        RECT 83.430 157.975 83.690 158.430 ;
        RECT 83.860 158.145 84.120 158.625 ;
        RECT 84.290 157.975 84.550 158.430 ;
        RECT 84.720 158.145 84.965 158.625 ;
        RECT 85.135 157.975 85.410 158.430 ;
        RECT 85.580 158.145 85.825 158.625 ;
        RECT 85.995 157.975 86.255 158.430 ;
        RECT 86.435 158.145 86.685 158.625 ;
        RECT 86.855 157.975 87.115 158.430 ;
        RECT 87.295 158.145 87.545 158.625 ;
        RECT 87.715 157.975 87.975 158.430 ;
        RECT 88.155 158.145 88.415 158.625 ;
        RECT 88.585 157.975 88.845 158.430 ;
        RECT 89.015 158.145 89.315 158.625 ;
        RECT 89.690 157.995 89.975 158.455 ;
        RECT 90.145 158.165 90.415 158.625 ;
        RECT 82.570 157.805 89.315 157.975 ;
        RECT 89.690 157.825 90.645 157.995 ;
        RECT 80.860 157.385 87.980 157.635 ;
        RECT 74.135 156.375 75.020 156.545 ;
        RECT 75.200 156.075 75.515 156.575 ;
        RECT 75.745 156.245 76.085 156.805 ;
        RECT 76.255 156.075 76.425 157.085 ;
        RECT 76.595 156.290 76.925 157.135 ;
        RECT 77.155 156.075 79.745 157.165 ;
        RECT 80.385 156.075 80.680 156.885 ;
        RECT 80.860 156.245 81.105 157.385 ;
        RECT 81.280 156.075 81.540 156.885 ;
        RECT 81.720 156.250 81.970 157.385 ;
        RECT 88.150 157.215 89.315 157.805 ;
        RECT 82.570 156.990 89.315 157.215 ;
        RECT 89.575 157.095 90.265 157.655 ;
        RECT 82.570 156.975 87.975 156.990 ;
        RECT 82.140 156.080 82.400 156.875 ;
        RECT 82.570 156.250 82.830 156.975 ;
        RECT 83.000 156.080 83.260 156.805 ;
        RECT 83.430 156.250 83.690 156.975 ;
        RECT 83.860 156.080 84.120 156.805 ;
        RECT 84.290 156.250 84.550 156.975 ;
        RECT 84.720 156.080 84.980 156.805 ;
        RECT 85.150 156.250 85.410 156.975 ;
        RECT 85.580 156.080 85.825 156.805 ;
        RECT 85.995 156.250 86.255 156.975 ;
        RECT 86.440 156.080 86.685 156.805 ;
        RECT 86.855 156.250 87.115 156.975 ;
        RECT 87.300 156.080 87.545 156.805 ;
        RECT 87.715 156.250 87.975 156.975 ;
        RECT 88.160 156.080 88.415 156.805 ;
        RECT 88.585 156.250 88.875 156.990 ;
        RECT 90.435 156.925 90.645 157.825 ;
        RECT 82.140 156.075 88.415 156.080 ;
        RECT 89.045 156.075 89.315 156.820 ;
        RECT 89.690 156.705 90.645 156.925 ;
        RECT 90.815 157.655 91.215 158.455 ;
        RECT 91.405 157.995 91.685 158.455 ;
        RECT 92.205 158.165 92.530 158.625 ;
        RECT 91.405 157.825 92.530 157.995 ;
        RECT 92.700 157.885 93.085 158.455 ;
        RECT 92.080 157.715 92.530 157.825 ;
        RECT 90.815 157.095 91.910 157.655 ;
        RECT 92.080 157.385 92.635 157.715 ;
        RECT 89.690 156.245 89.975 156.705 ;
        RECT 90.145 156.075 90.415 156.535 ;
        RECT 90.815 156.245 91.215 157.095 ;
        RECT 92.080 156.925 92.530 157.385 ;
        RECT 92.805 157.215 93.085 157.885 ;
        RECT 93.255 157.875 94.465 158.625 ;
        RECT 94.635 157.900 94.925 158.625 ;
        RECT 95.100 157.885 95.355 158.455 ;
        RECT 95.525 158.225 95.855 158.625 ;
        RECT 96.280 158.090 96.810 158.455 ;
        RECT 96.280 158.055 96.455 158.090 ;
        RECT 95.525 157.885 96.455 158.055 ;
        RECT 93.255 157.335 93.775 157.875 ;
        RECT 91.405 156.705 92.530 156.925 ;
        RECT 91.405 156.245 91.685 156.705 ;
        RECT 92.205 156.075 92.530 156.535 ;
        RECT 92.700 156.245 93.085 157.215 ;
        RECT 93.945 157.165 94.465 157.705 ;
        RECT 93.255 156.075 94.465 157.165 ;
        RECT 94.635 156.075 94.925 157.240 ;
        RECT 95.100 157.215 95.270 157.885 ;
        RECT 95.525 157.715 95.695 157.885 ;
        RECT 95.440 157.385 95.695 157.715 ;
        RECT 95.920 157.385 96.115 157.715 ;
        RECT 95.100 156.245 95.435 157.215 ;
        RECT 95.605 156.075 95.775 157.215 ;
        RECT 95.945 156.415 96.115 157.385 ;
        RECT 96.285 156.755 96.455 157.885 ;
        RECT 96.625 157.095 96.795 157.895 ;
        RECT 97.000 157.605 97.275 158.455 ;
        RECT 96.995 157.435 97.275 157.605 ;
        RECT 97.000 157.295 97.275 157.435 ;
        RECT 97.445 157.095 97.635 158.455 ;
        RECT 97.815 158.090 98.325 158.625 ;
        RECT 98.545 157.815 98.790 158.420 ;
        RECT 99.240 157.885 99.495 158.455 ;
        RECT 99.665 158.225 99.995 158.625 ;
        RECT 100.420 158.090 100.950 158.455 ;
        RECT 100.420 158.055 100.595 158.090 ;
        RECT 99.665 157.885 100.595 158.055 ;
        RECT 97.835 157.645 99.065 157.815 ;
        RECT 96.625 156.925 97.635 157.095 ;
        RECT 97.805 157.080 98.555 157.270 ;
        RECT 96.285 156.585 97.410 156.755 ;
        RECT 97.805 156.415 97.975 157.080 ;
        RECT 98.725 156.835 99.065 157.645 ;
        RECT 95.945 156.245 97.975 156.415 ;
        RECT 98.145 156.075 98.315 156.835 ;
        RECT 98.550 156.425 99.065 156.835 ;
        RECT 99.240 157.215 99.410 157.885 ;
        RECT 99.665 157.715 99.835 157.885 ;
        RECT 99.580 157.385 99.835 157.715 ;
        RECT 100.060 157.385 100.255 157.715 ;
        RECT 99.240 156.245 99.575 157.215 ;
        RECT 99.745 156.075 99.915 157.215 ;
        RECT 100.085 156.415 100.255 157.385 ;
        RECT 100.425 156.755 100.595 157.885 ;
        RECT 100.765 157.095 100.935 157.895 ;
        RECT 101.140 157.605 101.415 158.455 ;
        RECT 101.135 157.435 101.415 157.605 ;
        RECT 101.140 157.295 101.415 157.435 ;
        RECT 101.585 157.095 101.775 158.455 ;
        RECT 101.955 158.090 102.465 158.625 ;
        RECT 102.685 157.815 102.930 158.420 ;
        RECT 101.975 157.645 103.205 157.815 ;
        RECT 103.435 157.805 103.645 158.625 ;
        RECT 103.815 157.825 104.145 158.455 ;
        RECT 100.765 156.925 101.775 157.095 ;
        RECT 101.945 157.080 102.695 157.270 ;
        RECT 100.425 156.585 101.550 156.755 ;
        RECT 101.945 156.415 102.115 157.080 ;
        RECT 102.865 156.835 103.205 157.645 ;
        RECT 103.815 157.225 104.065 157.825 ;
        RECT 104.315 157.805 104.545 158.625 ;
        RECT 104.760 157.885 105.015 158.455 ;
        RECT 105.185 158.225 105.515 158.625 ;
        RECT 105.940 158.090 106.470 158.455 ;
        RECT 105.940 158.055 106.115 158.090 ;
        RECT 105.185 157.885 106.115 158.055 ;
        RECT 104.235 157.385 104.565 157.635 ;
        RECT 100.085 156.245 102.115 156.415 ;
        RECT 102.285 156.075 102.455 156.835 ;
        RECT 102.690 156.425 103.205 156.835 ;
        RECT 103.435 156.075 103.645 157.215 ;
        RECT 103.815 156.245 104.145 157.225 ;
        RECT 104.760 157.215 104.930 157.885 ;
        RECT 105.185 157.715 105.355 157.885 ;
        RECT 105.100 157.385 105.355 157.715 ;
        RECT 105.580 157.385 105.775 157.715 ;
        RECT 104.315 156.075 104.545 157.215 ;
        RECT 104.760 156.245 105.095 157.215 ;
        RECT 105.265 156.075 105.435 157.215 ;
        RECT 105.605 156.415 105.775 157.385 ;
        RECT 105.945 156.755 106.115 157.885 ;
        RECT 106.285 157.095 106.455 157.895 ;
        RECT 106.660 157.605 106.935 158.455 ;
        RECT 106.655 157.435 106.935 157.605 ;
        RECT 106.660 157.295 106.935 157.435 ;
        RECT 107.105 157.095 107.295 158.455 ;
        RECT 107.475 158.090 107.985 158.625 ;
        RECT 108.205 157.815 108.450 158.420 ;
        RECT 108.895 157.855 110.565 158.625 ;
        RECT 110.850 157.995 111.135 158.455 ;
        RECT 111.305 158.165 111.575 158.625 ;
        RECT 107.495 157.645 108.725 157.815 ;
        RECT 106.285 156.925 107.295 157.095 ;
        RECT 107.465 157.080 108.215 157.270 ;
        RECT 105.945 156.585 107.070 156.755 ;
        RECT 107.465 156.415 107.635 157.080 ;
        RECT 108.385 156.835 108.725 157.645 ;
        RECT 108.895 157.335 109.645 157.855 ;
        RECT 110.850 157.825 111.805 157.995 ;
        RECT 109.815 157.165 110.565 157.685 ;
        RECT 105.605 156.245 107.635 156.415 ;
        RECT 107.805 156.075 107.975 156.835 ;
        RECT 108.210 156.425 108.725 156.835 ;
        RECT 108.895 156.075 110.565 157.165 ;
        RECT 110.735 157.095 111.425 157.655 ;
        RECT 111.595 156.925 111.805 157.825 ;
        RECT 110.850 156.705 111.805 156.925 ;
        RECT 111.975 157.655 112.375 158.455 ;
        RECT 112.565 157.995 112.845 158.455 ;
        RECT 113.365 158.165 113.690 158.625 ;
        RECT 112.565 157.825 113.690 157.995 ;
        RECT 113.860 157.885 114.245 158.455 ;
        RECT 114.420 158.095 114.710 158.445 ;
        RECT 114.905 158.265 115.235 158.625 ;
        RECT 115.405 158.095 115.635 158.400 ;
        RECT 114.420 157.925 115.635 158.095 ;
        RECT 113.240 157.715 113.690 157.825 ;
        RECT 111.975 157.095 113.070 157.655 ;
        RECT 113.240 157.385 113.795 157.715 ;
        RECT 110.850 156.245 111.135 156.705 ;
        RECT 111.305 156.075 111.575 156.535 ;
        RECT 111.975 156.245 112.375 157.095 ;
        RECT 113.240 156.925 113.690 157.385 ;
        RECT 113.965 157.215 114.245 157.885 ;
        RECT 115.825 157.755 115.995 158.320 ;
        RECT 114.480 157.605 114.740 157.715 ;
        RECT 114.475 157.435 114.740 157.605 ;
        RECT 114.480 157.385 114.740 157.435 ;
        RECT 114.920 157.385 115.305 157.715 ;
        RECT 115.475 157.585 115.995 157.755 ;
        RECT 116.345 157.755 116.515 158.320 ;
        RECT 116.705 158.095 116.935 158.400 ;
        RECT 117.105 158.265 117.435 158.625 ;
        RECT 117.630 158.095 117.920 158.445 ;
        RECT 116.705 157.925 117.920 158.095 ;
        RECT 118.100 158.095 118.390 158.445 ;
        RECT 118.585 158.265 118.915 158.625 ;
        RECT 119.085 158.095 119.315 158.400 ;
        RECT 118.100 157.925 119.315 158.095 ;
        RECT 119.505 157.755 119.675 158.320 ;
        RECT 120.395 157.900 120.685 158.625 ;
        RECT 121.645 158.225 121.975 158.625 ;
        RECT 122.145 158.055 122.475 158.395 ;
        RECT 123.525 158.225 123.855 158.625 ;
        RECT 116.345 157.585 116.865 157.755 ;
        RECT 112.565 156.705 113.690 156.925 ;
        RECT 112.565 156.245 112.845 156.705 ;
        RECT 113.365 156.075 113.690 156.535 ;
        RECT 113.860 156.245 114.245 157.215 ;
        RECT 114.420 156.075 114.740 157.215 ;
        RECT 114.920 156.335 115.115 157.385 ;
        RECT 115.475 157.205 115.645 157.585 ;
        RECT 115.295 156.925 115.645 157.205 ;
        RECT 115.835 157.055 116.080 157.415 ;
        RECT 116.260 157.055 116.505 157.415 ;
        RECT 116.695 157.205 116.865 157.585 ;
        RECT 117.035 157.385 117.420 157.715 ;
        RECT 117.600 157.605 117.860 157.715 ;
        RECT 118.160 157.605 118.420 157.715 ;
        RECT 117.600 157.435 117.865 157.605 ;
        RECT 118.155 157.435 118.420 157.605 ;
        RECT 117.600 157.385 117.860 157.435 ;
        RECT 118.160 157.385 118.420 157.435 ;
        RECT 118.600 157.385 118.985 157.715 ;
        RECT 119.155 157.585 119.675 157.755 ;
        RECT 121.490 157.885 123.855 158.055 ;
        RECT 124.025 157.900 124.355 158.410 ;
        RECT 116.695 156.925 117.045 157.205 ;
        RECT 115.295 156.245 115.625 156.925 ;
        RECT 115.825 156.075 116.080 156.875 ;
        RECT 116.260 156.075 116.515 156.875 ;
        RECT 116.715 156.245 117.045 156.925 ;
        RECT 117.225 156.335 117.420 157.385 ;
        RECT 117.600 156.075 117.920 157.215 ;
        RECT 118.100 156.075 118.420 157.215 ;
        RECT 118.600 156.335 118.795 157.385 ;
        RECT 119.155 157.205 119.325 157.585 ;
        RECT 118.975 156.925 119.325 157.205 ;
        RECT 119.515 157.055 119.760 157.415 ;
        RECT 118.975 156.245 119.305 156.925 ;
        RECT 119.505 156.075 119.760 156.875 ;
        RECT 120.395 156.075 120.685 157.240 ;
        RECT 121.490 156.885 121.660 157.885 ;
        RECT 123.685 157.715 123.855 157.885 ;
        RECT 121.830 157.055 122.075 157.715 ;
        RECT 122.290 157.055 122.555 157.715 ;
        RECT 122.750 157.055 123.035 157.715 ;
        RECT 123.210 157.385 123.515 157.715 ;
        RECT 123.685 157.385 123.995 157.715 ;
        RECT 123.210 157.055 123.425 157.385 ;
        RECT 121.490 156.715 121.945 156.885 ;
        RECT 121.615 156.285 121.945 156.715 ;
        RECT 122.125 156.715 123.415 156.885 ;
        RECT 122.125 156.295 122.375 156.715 ;
        RECT 122.605 156.075 122.935 156.545 ;
        RECT 123.165 156.295 123.415 156.715 ;
        RECT 123.605 156.075 123.855 157.215 ;
        RECT 124.165 157.135 124.355 157.900 ;
        RECT 124.535 157.825 124.845 158.625 ;
        RECT 125.050 157.825 125.745 158.455 ;
        RECT 127.000 158.115 127.240 158.625 ;
        RECT 127.420 158.115 127.700 158.445 ;
        RECT 127.930 158.115 128.145 158.625 ;
        RECT 124.545 157.385 124.880 157.655 ;
        RECT 125.050 157.225 125.220 157.825 ;
        RECT 125.390 157.385 125.725 157.635 ;
        RECT 126.895 157.385 127.250 157.945 ;
        RECT 124.025 156.285 124.355 157.135 ;
        RECT 124.535 156.075 124.815 157.215 ;
        RECT 124.985 156.245 125.315 157.225 ;
        RECT 127.420 157.215 127.590 158.115 ;
        RECT 127.760 157.385 128.025 157.945 ;
        RECT 128.315 157.885 128.930 158.455 ;
        RECT 128.275 157.215 128.445 157.715 ;
        RECT 125.485 156.075 125.745 157.215 ;
        RECT 127.020 157.045 128.445 157.215 ;
        RECT 127.020 156.870 127.410 157.045 ;
        RECT 127.895 156.075 128.225 156.875 ;
        RECT 128.615 156.865 128.930 157.885 ;
        RECT 129.140 157.860 129.595 158.625 ;
        RECT 129.870 158.245 131.170 158.455 ;
        RECT 131.425 158.265 131.755 158.625 ;
        RECT 131.000 158.095 131.170 158.245 ;
        RECT 131.925 158.125 132.185 158.455 ;
        RECT 131.955 158.115 132.185 158.125 ;
        RECT 130.070 157.635 130.290 158.035 ;
        RECT 129.135 157.435 129.625 157.635 ;
        RECT 129.815 157.425 130.290 157.635 ;
        RECT 130.535 157.635 130.745 158.035 ;
        RECT 131.000 157.970 131.755 158.095 ;
        RECT 131.000 157.925 131.845 157.970 ;
        RECT 131.575 157.805 131.845 157.925 ;
        RECT 130.535 157.425 130.865 157.635 ;
        RECT 131.035 157.365 131.445 157.670 ;
        RECT 128.395 156.245 128.930 156.865 ;
        RECT 129.140 157.195 130.315 157.255 ;
        RECT 131.675 157.230 131.845 157.805 ;
        RECT 131.645 157.195 131.845 157.230 ;
        RECT 129.140 157.085 131.845 157.195 ;
        RECT 129.140 156.465 129.395 157.085 ;
        RECT 129.985 157.025 131.785 157.085 ;
        RECT 129.985 156.995 130.315 157.025 ;
        RECT 132.015 156.925 132.185 158.115 ;
        RECT 132.355 157.855 134.025 158.625 ;
        RECT 134.285 158.075 134.455 158.365 ;
        RECT 134.625 158.245 134.955 158.625 ;
        RECT 134.285 157.905 134.950 158.075 ;
        RECT 132.355 157.335 133.105 157.855 ;
        RECT 133.275 157.165 134.025 157.685 ;
        RECT 129.645 156.825 129.830 156.915 ;
        RECT 130.420 156.825 131.255 156.835 ;
        RECT 129.645 156.625 131.255 156.825 ;
        RECT 129.645 156.585 129.875 156.625 ;
        RECT 129.140 156.245 129.475 156.465 ;
        RECT 130.480 156.075 130.835 156.455 ;
        RECT 131.005 156.245 131.255 156.625 ;
        RECT 131.505 156.075 131.755 156.855 ;
        RECT 131.925 156.245 132.185 156.925 ;
        RECT 132.355 156.075 134.025 157.165 ;
        RECT 134.200 157.085 134.550 157.735 ;
        RECT 134.720 156.915 134.950 157.905 ;
        RECT 134.285 156.745 134.950 156.915 ;
        RECT 134.285 156.245 134.455 156.745 ;
        RECT 134.625 156.075 134.955 156.575 ;
        RECT 135.125 156.245 135.310 158.365 ;
        RECT 135.565 158.165 135.815 158.625 ;
        RECT 135.985 158.175 136.320 158.345 ;
        RECT 136.515 158.175 137.190 158.345 ;
        RECT 135.985 158.035 136.155 158.175 ;
        RECT 135.480 157.045 135.760 157.995 ;
        RECT 135.930 157.905 136.155 158.035 ;
        RECT 135.930 156.800 136.100 157.905 ;
        RECT 136.325 157.755 136.850 157.975 ;
        RECT 136.270 156.990 136.510 157.585 ;
        RECT 136.680 157.055 136.850 157.755 ;
        RECT 137.020 157.395 137.190 158.175 ;
        RECT 137.510 158.125 137.880 158.625 ;
        RECT 138.060 158.175 138.465 158.345 ;
        RECT 138.635 158.175 139.420 158.345 ;
        RECT 138.060 157.945 138.230 158.175 ;
        RECT 137.400 157.645 138.230 157.945 ;
        RECT 138.615 157.675 139.080 158.005 ;
        RECT 137.400 157.615 137.600 157.645 ;
        RECT 137.720 157.395 137.890 157.465 ;
        RECT 137.020 157.225 137.890 157.395 ;
        RECT 137.380 157.135 137.890 157.225 ;
        RECT 135.930 156.670 136.235 156.800 ;
        RECT 136.680 156.690 137.210 157.055 ;
        RECT 135.550 156.075 135.815 156.535 ;
        RECT 135.985 156.245 136.235 156.670 ;
        RECT 137.380 156.520 137.550 157.135 ;
        RECT 136.445 156.350 137.550 156.520 ;
        RECT 137.720 156.075 137.890 156.875 ;
        RECT 138.060 156.575 138.230 157.645 ;
        RECT 138.400 156.745 138.590 157.465 ;
        RECT 138.760 156.715 139.080 157.675 ;
        RECT 139.250 157.715 139.420 158.175 ;
        RECT 139.695 158.095 139.905 158.625 ;
        RECT 140.165 157.885 140.495 158.410 ;
        RECT 140.665 158.015 140.835 158.625 ;
        RECT 141.005 157.970 141.335 158.405 ;
        RECT 141.005 157.885 141.385 157.970 ;
        RECT 140.295 157.715 140.495 157.885 ;
        RECT 141.160 157.845 141.385 157.885 ;
        RECT 139.250 157.385 140.125 157.715 ;
        RECT 140.295 157.385 141.045 157.715 ;
        RECT 138.060 156.245 138.310 156.575 ;
        RECT 139.250 156.545 139.420 157.385 ;
        RECT 140.295 157.180 140.485 157.385 ;
        RECT 141.215 157.265 141.385 157.845 ;
        RECT 141.170 157.215 141.385 157.265 ;
        RECT 139.590 156.805 140.485 157.180 ;
        RECT 140.995 157.135 141.385 157.215 ;
        RECT 141.560 157.885 141.815 158.455 ;
        RECT 141.985 158.225 142.315 158.625 ;
        RECT 142.740 158.090 143.270 158.455 ;
        RECT 142.740 158.055 142.915 158.090 ;
        RECT 141.985 157.885 142.915 158.055 ;
        RECT 141.560 157.215 141.730 157.885 ;
        RECT 141.985 157.715 142.155 157.885 ;
        RECT 141.900 157.385 142.155 157.715 ;
        RECT 142.380 157.385 142.575 157.715 ;
        RECT 138.535 156.375 139.420 156.545 ;
        RECT 139.600 156.075 139.915 156.575 ;
        RECT 140.145 156.245 140.485 156.805 ;
        RECT 140.655 156.075 140.825 157.085 ;
        RECT 140.995 156.290 141.325 157.135 ;
        RECT 141.560 156.245 141.895 157.215 ;
        RECT 142.065 156.075 142.235 157.215 ;
        RECT 142.405 156.415 142.575 157.385 ;
        RECT 142.745 156.755 142.915 157.885 ;
        RECT 143.085 157.095 143.255 157.895 ;
        RECT 143.460 157.605 143.735 158.455 ;
        RECT 143.455 157.435 143.735 157.605 ;
        RECT 143.460 157.295 143.735 157.435 ;
        RECT 143.905 157.095 144.095 158.455 ;
        RECT 144.275 158.090 144.785 158.625 ;
        RECT 145.005 157.815 145.250 158.420 ;
        RECT 145.695 157.875 146.905 158.625 ;
        RECT 144.295 157.645 145.525 157.815 ;
        RECT 143.085 156.925 144.095 157.095 ;
        RECT 144.265 157.080 145.015 157.270 ;
        RECT 142.745 156.585 143.870 156.755 ;
        RECT 144.265 156.415 144.435 157.080 ;
        RECT 145.185 156.835 145.525 157.645 ;
        RECT 142.405 156.245 144.435 156.415 ;
        RECT 144.605 156.075 144.775 156.835 ;
        RECT 145.010 156.425 145.525 156.835 ;
        RECT 145.695 157.165 146.215 157.705 ;
        RECT 146.385 157.335 146.905 157.875 ;
        RECT 145.695 156.075 146.905 157.165 ;
        RECT 17.270 155.905 146.990 156.075 ;
        RECT 17.355 154.815 18.565 155.905 ;
        RECT 18.735 155.470 24.080 155.905 ;
        RECT 24.255 155.470 29.600 155.905 ;
        RECT 17.355 154.105 17.875 154.645 ;
        RECT 18.045 154.275 18.565 154.815 ;
        RECT 17.355 153.355 18.565 154.105 ;
        RECT 20.320 153.900 20.660 154.730 ;
        RECT 22.140 154.220 22.490 155.470 ;
        RECT 25.840 153.900 26.180 154.730 ;
        RECT 27.660 154.220 28.010 155.470 ;
        RECT 30.235 154.740 30.525 155.905 ;
        RECT 31.215 154.845 31.545 155.690 ;
        RECT 31.715 154.895 31.885 155.905 ;
        RECT 32.055 155.175 32.395 155.735 ;
        RECT 32.625 155.405 32.940 155.905 ;
        RECT 33.120 155.435 34.005 155.605 ;
        RECT 31.155 154.765 31.545 154.845 ;
        RECT 32.055 154.800 32.950 155.175 ;
        RECT 31.155 154.715 31.370 154.765 ;
        RECT 31.155 154.135 31.325 154.715 ;
        RECT 32.055 154.595 32.245 154.800 ;
        RECT 33.120 154.595 33.290 155.435 ;
        RECT 34.230 155.405 34.480 155.735 ;
        RECT 31.495 154.265 32.245 154.595 ;
        RECT 32.415 154.265 33.290 154.595 ;
        RECT 31.155 154.095 31.380 154.135 ;
        RECT 32.045 154.095 32.245 154.265 ;
        RECT 18.735 153.355 24.080 153.900 ;
        RECT 24.255 153.355 29.600 153.900 ;
        RECT 30.235 153.355 30.525 154.080 ;
        RECT 31.155 154.010 31.535 154.095 ;
        RECT 31.205 153.575 31.535 154.010 ;
        RECT 31.705 153.355 31.875 153.965 ;
        RECT 32.045 153.570 32.375 154.095 ;
        RECT 32.635 153.355 32.845 153.885 ;
        RECT 33.120 153.805 33.290 154.265 ;
        RECT 33.460 154.305 33.780 155.265 ;
        RECT 33.950 154.515 34.140 155.235 ;
        RECT 34.310 154.335 34.480 155.405 ;
        RECT 34.650 155.105 34.820 155.905 ;
        RECT 34.990 155.460 36.095 155.630 ;
        RECT 34.990 154.845 35.160 155.460 ;
        RECT 36.305 155.310 36.555 155.735 ;
        RECT 36.725 155.445 36.990 155.905 ;
        RECT 35.330 154.925 35.860 155.290 ;
        RECT 36.305 155.180 36.610 155.310 ;
        RECT 34.650 154.755 35.160 154.845 ;
        RECT 34.650 154.585 35.520 154.755 ;
        RECT 34.650 154.515 34.820 154.585 ;
        RECT 34.940 154.335 35.140 154.365 ;
        RECT 33.460 153.975 33.925 154.305 ;
        RECT 34.310 154.035 35.140 154.335 ;
        RECT 34.310 153.805 34.480 154.035 ;
        RECT 33.120 153.635 33.905 153.805 ;
        RECT 34.075 153.635 34.480 153.805 ;
        RECT 34.660 153.355 35.030 153.855 ;
        RECT 35.350 153.805 35.520 154.585 ;
        RECT 35.690 154.225 35.860 154.925 ;
        RECT 36.030 154.395 36.270 154.990 ;
        RECT 35.690 154.005 36.215 154.225 ;
        RECT 36.440 154.075 36.610 155.180 ;
        RECT 36.385 153.945 36.610 154.075 ;
        RECT 36.780 153.985 37.060 154.935 ;
        RECT 36.385 153.805 36.555 153.945 ;
        RECT 35.350 153.635 36.025 153.805 ;
        RECT 36.220 153.635 36.555 153.805 ;
        RECT 36.725 153.355 36.975 153.815 ;
        RECT 37.230 153.615 37.415 155.735 ;
        RECT 37.585 155.405 37.915 155.905 ;
        RECT 38.085 155.235 38.255 155.735 ;
        RECT 37.590 155.065 38.255 155.235 ;
        RECT 37.590 154.075 37.820 155.065 ;
        RECT 37.990 154.245 38.340 154.895 ;
        RECT 38.525 154.845 38.855 155.695 ;
        RECT 38.525 154.080 38.715 154.845 ;
        RECT 39.025 154.765 39.275 155.905 ;
        RECT 39.465 155.265 39.715 155.685 ;
        RECT 39.945 155.435 40.275 155.905 ;
        RECT 40.505 155.265 40.755 155.685 ;
        RECT 39.465 155.095 40.755 155.265 ;
        RECT 40.935 155.265 41.265 155.695 ;
        RECT 40.935 155.095 41.390 155.265 ;
        RECT 39.455 154.595 39.670 154.925 ;
        RECT 38.885 154.265 39.195 154.595 ;
        RECT 39.365 154.265 39.670 154.595 ;
        RECT 39.845 154.265 40.130 154.925 ;
        RECT 40.325 154.265 40.590 154.925 ;
        RECT 40.805 154.265 41.050 154.925 ;
        RECT 39.025 154.095 39.195 154.265 ;
        RECT 41.220 154.095 41.390 155.095 ;
        RECT 42.235 154.955 42.525 155.725 ;
        RECT 43.095 155.365 43.355 155.725 ;
        RECT 43.525 155.535 43.855 155.905 ;
        RECT 44.025 155.365 44.285 155.725 ;
        RECT 43.095 155.135 44.285 155.365 ;
        RECT 44.475 155.185 44.805 155.905 ;
        RECT 44.975 154.955 45.240 155.725 ;
        RECT 42.235 154.775 44.730 154.955 ;
        RECT 42.205 154.265 42.475 154.595 ;
        RECT 42.655 154.265 43.090 154.595 ;
        RECT 43.270 154.265 43.845 154.595 ;
        RECT 44.025 154.265 44.305 154.595 ;
        RECT 37.590 153.905 38.255 154.075 ;
        RECT 37.585 153.355 37.915 153.735 ;
        RECT 38.085 153.615 38.255 153.905 ;
        RECT 38.525 153.570 38.855 154.080 ;
        RECT 39.025 153.925 41.390 154.095 ;
        RECT 44.505 154.085 44.730 154.775 ;
        RECT 39.025 153.355 39.355 153.755 ;
        RECT 40.405 153.585 40.735 153.925 ;
        RECT 42.245 153.895 44.730 154.085 ;
        RECT 40.905 153.355 41.235 153.755 ;
        RECT 42.245 153.535 42.470 153.895 ;
        RECT 42.650 153.355 42.980 153.725 ;
        RECT 43.160 153.535 43.415 153.895 ;
        RECT 43.980 153.355 44.725 153.725 ;
        RECT 44.905 153.535 45.240 154.955 ;
        RECT 45.435 155.015 45.695 155.725 ;
        RECT 45.865 155.195 46.195 155.905 ;
        RECT 46.365 155.015 46.595 155.725 ;
        RECT 45.435 154.775 46.595 155.015 ;
        RECT 46.775 154.995 47.045 155.725 ;
        RECT 47.225 155.175 47.565 155.905 ;
        RECT 46.775 154.775 47.545 154.995 ;
        RECT 45.425 154.265 45.725 154.595 ;
        RECT 45.905 154.285 46.430 154.595 ;
        RECT 46.610 154.285 47.075 154.595 ;
        RECT 45.435 153.355 45.725 154.085 ;
        RECT 45.905 153.645 46.135 154.285 ;
        RECT 47.255 154.105 47.545 154.775 ;
        RECT 46.315 153.905 47.545 154.105 ;
        RECT 46.315 153.535 46.625 153.905 ;
        RECT 46.805 153.355 47.475 153.725 ;
        RECT 47.735 153.535 47.995 155.725 ;
        RECT 48.175 155.470 53.520 155.905 ;
        RECT 49.760 153.900 50.100 154.730 ;
        RECT 51.580 154.220 51.930 155.470 ;
        RECT 53.695 154.815 55.365 155.905 ;
        RECT 53.695 154.125 54.445 154.645 ;
        RECT 54.615 154.295 55.365 154.815 ;
        RECT 55.995 154.740 56.285 155.905 ;
        RECT 57.575 155.235 57.855 155.905 ;
        RECT 58.025 155.015 58.325 155.565 ;
        RECT 58.525 155.185 58.855 155.905 ;
        RECT 59.045 155.185 59.505 155.735 ;
        RECT 59.675 155.395 59.935 155.905 ;
        RECT 57.390 154.595 57.655 154.955 ;
        RECT 58.025 154.845 58.965 155.015 ;
        RECT 58.795 154.595 58.965 154.845 ;
        RECT 57.390 154.345 58.065 154.595 ;
        RECT 58.285 154.345 58.625 154.595 ;
        RECT 58.795 154.265 59.085 154.595 ;
        RECT 58.795 154.175 58.965 154.265 ;
        RECT 48.175 153.355 53.520 153.900 ;
        RECT 53.695 153.355 55.365 154.125 ;
        RECT 55.995 153.355 56.285 154.080 ;
        RECT 57.575 153.985 58.965 154.175 ;
        RECT 57.575 153.625 57.905 153.985 ;
        RECT 59.255 153.815 59.505 155.185 ;
        RECT 59.675 154.345 60.015 155.225 ;
        RECT 60.185 154.515 60.355 155.735 ;
        RECT 60.595 155.400 61.210 155.905 ;
        RECT 60.595 154.865 60.845 155.230 ;
        RECT 61.015 155.225 61.210 155.400 ;
        RECT 61.380 155.395 61.855 155.735 ;
        RECT 62.025 155.360 62.240 155.905 ;
        RECT 61.015 155.035 61.345 155.225 ;
        RECT 61.565 154.865 62.280 155.160 ;
        RECT 62.450 155.035 62.725 155.735 ;
        RECT 60.595 154.695 62.385 154.865 ;
        RECT 60.185 154.265 60.980 154.515 ;
        RECT 60.185 154.175 60.435 154.265 ;
        RECT 58.525 153.355 58.775 153.815 ;
        RECT 58.945 153.525 59.505 153.815 ;
        RECT 59.675 153.355 59.935 154.175 ;
        RECT 60.105 153.755 60.435 154.175 ;
        RECT 61.150 153.840 61.405 154.695 ;
        RECT 60.615 153.575 61.405 153.840 ;
        RECT 61.575 153.995 61.985 154.515 ;
        RECT 62.155 154.265 62.385 154.695 ;
        RECT 62.555 154.005 62.725 155.035 ;
        RECT 61.575 153.575 61.775 153.995 ;
        RECT 61.965 153.355 62.295 153.815 ;
        RECT 62.465 153.525 62.725 154.005 ;
        RECT 62.930 155.115 63.465 155.735 ;
        RECT 62.930 154.095 63.245 155.115 ;
        RECT 63.635 155.105 63.965 155.905 ;
        RECT 65.195 155.470 70.540 155.905 ;
        RECT 70.715 155.470 76.060 155.905 ;
        RECT 64.450 154.935 64.840 155.110 ;
        RECT 63.415 154.765 64.840 154.935 ;
        RECT 63.415 154.265 63.585 154.765 ;
        RECT 62.930 153.525 63.545 154.095 ;
        RECT 63.835 154.035 64.100 154.595 ;
        RECT 64.270 153.865 64.440 154.765 ;
        RECT 64.610 154.035 64.965 154.595 ;
        RECT 66.780 153.900 67.120 154.730 ;
        RECT 68.600 154.220 68.950 155.470 ;
        RECT 72.300 153.900 72.640 154.730 ;
        RECT 74.120 154.220 74.470 155.470 ;
        RECT 76.730 155.115 77.265 155.735 ;
        RECT 76.730 154.095 77.045 155.115 ;
        RECT 77.435 155.105 77.765 155.905 ;
        RECT 78.250 154.935 78.640 155.110 ;
        RECT 77.215 154.765 78.640 154.935 ;
        RECT 79.055 154.765 79.265 155.905 ;
        RECT 77.215 154.265 77.385 154.765 ;
        RECT 63.715 153.355 63.930 153.865 ;
        RECT 64.160 153.535 64.440 153.865 ;
        RECT 64.620 153.355 64.860 153.865 ;
        RECT 65.195 153.355 70.540 153.900 ;
        RECT 70.715 153.355 76.060 153.900 ;
        RECT 76.730 153.525 77.345 154.095 ;
        RECT 77.635 154.035 77.900 154.595 ;
        RECT 78.070 153.865 78.240 154.765 ;
        RECT 79.435 154.755 79.765 155.735 ;
        RECT 79.935 154.765 80.165 155.905 ;
        RECT 80.375 154.815 81.585 155.905 ;
        RECT 78.410 154.035 78.765 154.595 ;
        RECT 77.515 153.355 77.730 153.865 ;
        RECT 77.960 153.535 78.240 153.865 ;
        RECT 78.420 153.355 78.660 153.865 ;
        RECT 79.055 153.355 79.265 154.175 ;
        RECT 79.435 154.155 79.685 154.755 ;
        RECT 79.855 154.345 80.185 154.595 ;
        RECT 79.435 153.525 79.765 154.155 ;
        RECT 79.935 153.355 80.165 154.175 ;
        RECT 80.375 154.105 80.895 154.645 ;
        RECT 81.065 154.275 81.585 154.815 ;
        RECT 81.755 154.740 82.045 155.905 ;
        RECT 82.215 154.815 85.725 155.905 ;
        RECT 85.895 154.815 87.105 155.905 ;
        RECT 87.335 154.845 87.665 155.690 ;
        RECT 87.835 154.895 88.005 155.905 ;
        RECT 88.175 155.175 88.515 155.735 ;
        RECT 88.745 155.405 89.060 155.905 ;
        RECT 89.240 155.435 90.125 155.605 ;
        RECT 82.215 154.125 83.865 154.645 ;
        RECT 84.035 154.295 85.725 154.815 ;
        RECT 80.375 153.355 81.585 154.105 ;
        RECT 81.755 153.355 82.045 154.080 ;
        RECT 82.215 153.355 85.725 154.125 ;
        RECT 85.895 154.105 86.415 154.645 ;
        RECT 86.585 154.275 87.105 154.815 ;
        RECT 87.275 154.765 87.665 154.845 ;
        RECT 88.175 154.800 89.070 155.175 ;
        RECT 87.275 154.715 87.490 154.765 ;
        RECT 87.275 154.135 87.445 154.715 ;
        RECT 88.175 154.595 88.365 154.800 ;
        RECT 89.240 154.595 89.410 155.435 ;
        RECT 90.350 155.405 90.600 155.735 ;
        RECT 87.615 154.265 88.365 154.595 ;
        RECT 88.535 154.265 89.410 154.595 ;
        RECT 85.895 153.355 87.105 154.105 ;
        RECT 87.275 154.095 87.500 154.135 ;
        RECT 88.165 154.095 88.365 154.265 ;
        RECT 87.275 154.010 87.655 154.095 ;
        RECT 87.325 153.575 87.655 154.010 ;
        RECT 87.825 153.355 87.995 153.965 ;
        RECT 88.165 153.570 88.495 154.095 ;
        RECT 88.755 153.355 88.965 153.885 ;
        RECT 89.240 153.805 89.410 154.265 ;
        RECT 89.580 154.305 89.900 155.265 ;
        RECT 90.070 154.515 90.260 155.235 ;
        RECT 90.430 154.335 90.600 155.405 ;
        RECT 90.770 155.105 90.940 155.905 ;
        RECT 91.110 155.460 92.215 155.630 ;
        RECT 91.110 154.845 91.280 155.460 ;
        RECT 92.425 155.310 92.675 155.735 ;
        RECT 92.845 155.445 93.110 155.905 ;
        RECT 91.450 154.925 91.980 155.290 ;
        RECT 92.425 155.180 92.730 155.310 ;
        RECT 90.770 154.755 91.280 154.845 ;
        RECT 90.770 154.585 91.640 154.755 ;
        RECT 90.770 154.515 90.940 154.585 ;
        RECT 91.060 154.335 91.260 154.365 ;
        RECT 89.580 153.975 90.045 154.305 ;
        RECT 90.430 154.035 91.260 154.335 ;
        RECT 90.430 153.805 90.600 154.035 ;
        RECT 89.240 153.635 90.025 153.805 ;
        RECT 90.195 153.635 90.600 153.805 ;
        RECT 90.780 153.355 91.150 153.855 ;
        RECT 91.470 153.805 91.640 154.585 ;
        RECT 91.810 154.225 91.980 154.925 ;
        RECT 92.150 154.395 92.390 154.990 ;
        RECT 91.810 154.005 92.335 154.225 ;
        RECT 92.560 154.075 92.730 155.180 ;
        RECT 92.505 153.945 92.730 154.075 ;
        RECT 92.900 153.985 93.180 154.935 ;
        RECT 92.505 153.805 92.675 153.945 ;
        RECT 91.470 153.635 92.145 153.805 ;
        RECT 92.340 153.635 92.675 153.805 ;
        RECT 92.845 153.355 93.095 153.815 ;
        RECT 93.350 153.615 93.535 155.735 ;
        RECT 93.705 155.405 94.035 155.905 ;
        RECT 94.205 155.235 94.375 155.735 ;
        RECT 93.710 155.065 94.375 155.235 ;
        RECT 94.725 155.235 94.895 155.735 ;
        RECT 95.065 155.405 95.395 155.905 ;
        RECT 94.725 155.065 95.390 155.235 ;
        RECT 93.710 154.075 93.940 155.065 ;
        RECT 94.110 154.245 94.460 154.895 ;
        RECT 94.640 154.245 94.990 154.895 ;
        RECT 95.160 154.075 95.390 155.065 ;
        RECT 93.710 153.905 94.375 154.075 ;
        RECT 93.705 153.355 94.035 153.735 ;
        RECT 94.205 153.615 94.375 153.905 ;
        RECT 94.725 153.905 95.390 154.075 ;
        RECT 94.725 153.615 94.895 153.905 ;
        RECT 95.065 153.355 95.395 153.735 ;
        RECT 95.565 153.615 95.750 155.735 ;
        RECT 95.990 155.445 96.255 155.905 ;
        RECT 96.425 155.310 96.675 155.735 ;
        RECT 96.885 155.460 97.990 155.630 ;
        RECT 96.370 155.180 96.675 155.310 ;
        RECT 95.920 153.985 96.200 154.935 ;
        RECT 96.370 154.075 96.540 155.180 ;
        RECT 96.710 154.395 96.950 154.990 ;
        RECT 97.120 154.925 97.650 155.290 ;
        RECT 97.120 154.225 97.290 154.925 ;
        RECT 97.820 154.845 97.990 155.460 ;
        RECT 98.160 155.105 98.330 155.905 ;
        RECT 98.500 155.405 98.750 155.735 ;
        RECT 98.975 155.435 99.860 155.605 ;
        RECT 97.820 154.755 98.330 154.845 ;
        RECT 96.370 153.945 96.595 154.075 ;
        RECT 96.765 154.005 97.290 154.225 ;
        RECT 97.460 154.585 98.330 154.755 ;
        RECT 96.005 153.355 96.255 153.815 ;
        RECT 96.425 153.805 96.595 153.945 ;
        RECT 97.460 153.805 97.630 154.585 ;
        RECT 98.160 154.515 98.330 154.585 ;
        RECT 97.840 154.335 98.040 154.365 ;
        RECT 98.500 154.335 98.670 155.405 ;
        RECT 98.840 154.515 99.030 155.235 ;
        RECT 97.840 154.035 98.670 154.335 ;
        RECT 99.200 154.305 99.520 155.265 ;
        RECT 96.425 153.635 96.760 153.805 ;
        RECT 96.955 153.635 97.630 153.805 ;
        RECT 97.950 153.355 98.320 153.855 ;
        RECT 98.500 153.805 98.670 154.035 ;
        RECT 99.055 153.975 99.520 154.305 ;
        RECT 99.690 154.595 99.860 155.435 ;
        RECT 100.040 155.405 100.355 155.905 ;
        RECT 100.585 155.175 100.925 155.735 ;
        RECT 100.030 154.800 100.925 155.175 ;
        RECT 101.095 154.895 101.265 155.905 ;
        RECT 100.735 154.595 100.925 154.800 ;
        RECT 101.435 154.845 101.765 155.690 ;
        RECT 103.030 155.275 103.315 155.735 ;
        RECT 103.485 155.445 103.755 155.905 ;
        RECT 103.030 155.055 103.985 155.275 ;
        RECT 101.435 154.765 101.825 154.845 ;
        RECT 101.610 154.715 101.825 154.765 ;
        RECT 99.690 154.265 100.565 154.595 ;
        RECT 100.735 154.265 101.485 154.595 ;
        RECT 99.690 153.805 99.860 154.265 ;
        RECT 100.735 154.095 100.935 154.265 ;
        RECT 101.655 154.135 101.825 154.715 ;
        RECT 102.915 154.325 103.605 154.885 ;
        RECT 103.775 154.155 103.985 155.055 ;
        RECT 101.600 154.095 101.825 154.135 ;
        RECT 98.500 153.635 98.905 153.805 ;
        RECT 99.075 153.635 99.860 153.805 ;
        RECT 100.135 153.355 100.345 153.885 ;
        RECT 100.605 153.570 100.935 154.095 ;
        RECT 101.445 154.010 101.825 154.095 ;
        RECT 101.105 153.355 101.275 153.965 ;
        RECT 101.445 153.575 101.775 154.010 ;
        RECT 103.030 153.985 103.985 154.155 ;
        RECT 104.155 154.885 104.555 155.735 ;
        RECT 104.745 155.275 105.025 155.735 ;
        RECT 105.545 155.445 105.870 155.905 ;
        RECT 104.745 155.055 105.870 155.275 ;
        RECT 104.155 154.325 105.250 154.885 ;
        RECT 105.420 154.595 105.870 155.055 ;
        RECT 106.040 154.765 106.425 155.735 ;
        RECT 103.030 153.525 103.315 153.985 ;
        RECT 103.485 153.355 103.755 153.815 ;
        RECT 104.155 153.525 104.555 154.325 ;
        RECT 105.420 154.265 105.975 154.595 ;
        RECT 105.420 154.155 105.870 154.265 ;
        RECT 104.745 153.985 105.870 154.155 ;
        RECT 106.145 154.095 106.425 154.765 ;
        RECT 107.515 154.740 107.805 155.905 ;
        RECT 108.035 154.845 108.365 155.690 ;
        RECT 108.535 154.895 108.705 155.905 ;
        RECT 108.875 155.175 109.215 155.735 ;
        RECT 109.445 155.405 109.760 155.905 ;
        RECT 109.940 155.435 110.825 155.605 ;
        RECT 107.975 154.765 108.365 154.845 ;
        RECT 108.875 154.800 109.770 155.175 ;
        RECT 104.745 153.525 105.025 153.985 ;
        RECT 105.545 153.355 105.870 153.815 ;
        RECT 106.040 153.525 106.425 154.095 ;
        RECT 107.975 154.715 108.190 154.765 ;
        RECT 107.975 154.135 108.145 154.715 ;
        RECT 108.875 154.595 109.065 154.800 ;
        RECT 109.940 154.595 110.110 155.435 ;
        RECT 111.050 155.405 111.300 155.735 ;
        RECT 108.315 154.265 109.065 154.595 ;
        RECT 109.235 154.265 110.110 154.595 ;
        RECT 107.975 154.095 108.200 154.135 ;
        RECT 108.865 154.095 109.065 154.265 ;
        RECT 107.515 153.355 107.805 154.080 ;
        RECT 107.975 154.010 108.355 154.095 ;
        RECT 108.025 153.575 108.355 154.010 ;
        RECT 108.525 153.355 108.695 153.965 ;
        RECT 108.865 153.570 109.195 154.095 ;
        RECT 109.455 153.355 109.665 153.885 ;
        RECT 109.940 153.805 110.110 154.265 ;
        RECT 110.280 154.305 110.600 155.265 ;
        RECT 110.770 154.515 110.960 155.235 ;
        RECT 111.130 154.335 111.300 155.405 ;
        RECT 111.470 155.105 111.640 155.905 ;
        RECT 111.810 155.460 112.915 155.630 ;
        RECT 111.810 154.845 111.980 155.460 ;
        RECT 113.125 155.310 113.375 155.735 ;
        RECT 113.545 155.445 113.810 155.905 ;
        RECT 112.150 154.925 112.680 155.290 ;
        RECT 113.125 155.180 113.430 155.310 ;
        RECT 111.470 154.755 111.980 154.845 ;
        RECT 111.470 154.585 112.340 154.755 ;
        RECT 111.470 154.515 111.640 154.585 ;
        RECT 111.760 154.335 111.960 154.365 ;
        RECT 110.280 153.975 110.745 154.305 ;
        RECT 111.130 154.035 111.960 154.335 ;
        RECT 111.130 153.805 111.300 154.035 ;
        RECT 109.940 153.635 110.725 153.805 ;
        RECT 110.895 153.635 111.300 153.805 ;
        RECT 111.480 153.355 111.850 153.855 ;
        RECT 112.170 153.805 112.340 154.585 ;
        RECT 112.510 154.225 112.680 154.925 ;
        RECT 112.850 154.395 113.090 154.990 ;
        RECT 112.510 154.005 113.035 154.225 ;
        RECT 113.260 154.075 113.430 155.180 ;
        RECT 113.205 153.945 113.430 154.075 ;
        RECT 113.600 153.985 113.880 154.935 ;
        RECT 113.205 153.805 113.375 153.945 ;
        RECT 112.170 153.635 112.845 153.805 ;
        RECT 113.040 153.635 113.375 153.805 ;
        RECT 113.545 153.355 113.795 153.815 ;
        RECT 114.050 153.615 114.235 155.735 ;
        RECT 114.405 155.405 114.735 155.905 ;
        RECT 114.905 155.235 115.075 155.735 ;
        RECT 114.410 155.065 115.075 155.235 ;
        RECT 114.410 154.075 114.640 155.065 ;
        RECT 114.810 154.245 115.160 154.895 ;
        RECT 115.340 154.765 115.675 155.735 ;
        RECT 115.845 154.765 116.015 155.905 ;
        RECT 116.185 155.565 118.215 155.735 ;
        RECT 115.340 154.095 115.510 154.765 ;
        RECT 116.185 154.595 116.355 155.565 ;
        RECT 115.680 154.265 115.935 154.595 ;
        RECT 116.160 154.265 116.355 154.595 ;
        RECT 116.525 155.225 117.650 155.395 ;
        RECT 115.765 154.095 115.935 154.265 ;
        RECT 116.525 154.095 116.695 155.225 ;
        RECT 114.410 153.905 115.075 154.075 ;
        RECT 114.405 153.355 114.735 153.735 ;
        RECT 114.905 153.615 115.075 153.905 ;
        RECT 115.340 153.525 115.595 154.095 ;
        RECT 115.765 153.925 116.695 154.095 ;
        RECT 116.865 154.885 117.875 155.055 ;
        RECT 116.865 154.085 117.035 154.885 ;
        RECT 116.520 153.890 116.695 153.925 ;
        RECT 115.765 153.355 116.095 153.755 ;
        RECT 116.520 153.525 117.050 153.890 ;
        RECT 117.240 153.865 117.515 154.685 ;
        RECT 117.235 153.695 117.515 153.865 ;
        RECT 117.240 153.525 117.515 153.695 ;
        RECT 117.685 153.525 117.875 154.885 ;
        RECT 118.045 154.900 118.215 155.565 ;
        RECT 118.385 155.145 118.555 155.905 ;
        RECT 118.790 155.145 119.305 155.555 ;
        RECT 118.045 154.710 118.795 154.900 ;
        RECT 118.965 154.335 119.305 155.145 ;
        RECT 119.590 155.275 119.875 155.735 ;
        RECT 120.045 155.445 120.315 155.905 ;
        RECT 119.590 155.055 120.545 155.275 ;
        RECT 118.075 154.165 119.305 154.335 ;
        RECT 119.475 154.325 120.165 154.885 ;
        RECT 118.055 153.355 118.565 153.890 ;
        RECT 118.785 153.560 119.030 154.165 ;
        RECT 120.335 154.155 120.545 155.055 ;
        RECT 119.590 153.985 120.545 154.155 ;
        RECT 120.715 154.885 121.115 155.735 ;
        RECT 121.305 155.275 121.585 155.735 ;
        RECT 122.105 155.445 122.430 155.905 ;
        RECT 121.305 155.055 122.430 155.275 ;
        RECT 120.715 154.325 121.810 154.885 ;
        RECT 121.980 154.595 122.430 155.055 ;
        RECT 122.600 154.765 122.985 155.735 ;
        RECT 123.160 155.105 123.415 155.905 ;
        RECT 123.615 155.055 123.945 155.735 ;
        RECT 119.590 153.525 119.875 153.985 ;
        RECT 120.045 153.355 120.315 153.815 ;
        RECT 120.715 153.525 121.115 154.325 ;
        RECT 121.980 154.265 122.535 154.595 ;
        RECT 121.980 154.155 122.430 154.265 ;
        RECT 121.305 153.985 122.430 154.155 ;
        RECT 122.705 154.095 122.985 154.765 ;
        RECT 123.160 154.565 123.405 154.925 ;
        RECT 123.595 154.775 123.945 155.055 ;
        RECT 123.595 154.395 123.765 154.775 ;
        RECT 124.125 154.595 124.320 155.645 ;
        RECT 124.500 154.765 124.820 155.905 ;
        RECT 125.000 154.765 125.335 155.735 ;
        RECT 125.505 154.765 125.675 155.905 ;
        RECT 125.845 155.565 127.875 155.735 ;
        RECT 121.305 153.525 121.585 153.985 ;
        RECT 122.105 153.355 122.430 153.815 ;
        RECT 122.600 153.525 122.985 154.095 ;
        RECT 123.245 154.225 123.765 154.395 ;
        RECT 123.935 154.265 124.320 154.595 ;
        RECT 124.500 154.545 124.760 154.595 ;
        RECT 124.500 154.375 124.765 154.545 ;
        RECT 124.500 154.265 124.760 154.375 ;
        RECT 123.245 153.660 123.415 154.225 ;
        RECT 125.000 154.095 125.170 154.765 ;
        RECT 125.845 154.595 126.015 155.565 ;
        RECT 125.340 154.265 125.595 154.595 ;
        RECT 125.820 154.265 126.015 154.595 ;
        RECT 126.185 155.225 127.310 155.395 ;
        RECT 125.425 154.095 125.595 154.265 ;
        RECT 126.185 154.095 126.355 155.225 ;
        RECT 123.605 153.885 124.820 154.055 ;
        RECT 123.605 153.580 123.835 153.885 ;
        RECT 124.005 153.355 124.335 153.715 ;
        RECT 124.530 153.535 124.820 153.885 ;
        RECT 125.000 153.525 125.255 154.095 ;
        RECT 125.425 153.925 126.355 154.095 ;
        RECT 126.525 154.885 127.535 155.055 ;
        RECT 126.525 154.085 126.695 154.885 ;
        RECT 126.180 153.890 126.355 153.925 ;
        RECT 125.425 153.355 125.755 153.755 ;
        RECT 126.180 153.525 126.710 153.890 ;
        RECT 126.900 153.865 127.175 154.685 ;
        RECT 126.895 153.695 127.175 153.865 ;
        RECT 126.900 153.525 127.175 153.695 ;
        RECT 127.345 153.525 127.535 154.885 ;
        RECT 127.705 154.900 127.875 155.565 ;
        RECT 128.045 155.145 128.215 155.905 ;
        RECT 128.450 155.145 128.965 155.555 ;
        RECT 127.705 154.710 128.455 154.900 ;
        RECT 128.625 154.335 128.965 155.145 ;
        RECT 127.735 154.165 128.965 154.335 ;
        RECT 129.135 154.765 129.520 155.735 ;
        RECT 129.690 155.445 130.015 155.905 ;
        RECT 130.535 155.275 130.815 155.735 ;
        RECT 129.690 155.055 130.815 155.275 ;
        RECT 127.715 153.355 128.225 153.890 ;
        RECT 128.445 153.560 128.690 154.165 ;
        RECT 129.135 154.095 129.415 154.765 ;
        RECT 129.690 154.595 130.140 155.055 ;
        RECT 131.005 154.885 131.405 155.735 ;
        RECT 131.805 155.445 132.075 155.905 ;
        RECT 132.245 155.275 132.530 155.735 ;
        RECT 129.585 154.265 130.140 154.595 ;
        RECT 130.310 154.325 131.405 154.885 ;
        RECT 129.690 154.155 130.140 154.265 ;
        RECT 129.135 153.525 129.520 154.095 ;
        RECT 129.690 153.985 130.815 154.155 ;
        RECT 129.690 153.355 130.015 153.815 ;
        RECT 130.535 153.525 130.815 153.985 ;
        RECT 131.005 153.525 131.405 154.325 ;
        RECT 131.575 155.055 132.530 155.275 ;
        RECT 131.575 154.155 131.785 155.055 ;
        RECT 131.955 154.325 132.645 154.885 ;
        RECT 133.275 154.740 133.565 155.905 ;
        RECT 134.285 155.235 134.455 155.735 ;
        RECT 134.625 155.405 134.955 155.905 ;
        RECT 134.285 155.065 134.950 155.235 ;
        RECT 134.200 154.245 134.550 154.895 ;
        RECT 131.575 153.985 132.530 154.155 ;
        RECT 131.805 153.355 132.075 153.815 ;
        RECT 132.245 153.525 132.530 153.985 ;
        RECT 133.275 153.355 133.565 154.080 ;
        RECT 134.720 154.075 134.950 155.065 ;
        RECT 134.285 153.905 134.950 154.075 ;
        RECT 134.285 153.615 134.455 153.905 ;
        RECT 134.625 153.355 134.955 153.735 ;
        RECT 135.125 153.615 135.310 155.735 ;
        RECT 135.550 155.445 135.815 155.905 ;
        RECT 135.985 155.310 136.235 155.735 ;
        RECT 136.445 155.460 137.550 155.630 ;
        RECT 135.930 155.180 136.235 155.310 ;
        RECT 135.480 153.985 135.760 154.935 ;
        RECT 135.930 154.075 136.100 155.180 ;
        RECT 136.270 154.395 136.510 154.990 ;
        RECT 136.680 154.925 137.210 155.290 ;
        RECT 136.680 154.225 136.850 154.925 ;
        RECT 137.380 154.845 137.550 155.460 ;
        RECT 137.720 155.105 137.890 155.905 ;
        RECT 138.060 155.405 138.310 155.735 ;
        RECT 138.535 155.435 139.420 155.605 ;
        RECT 137.380 154.755 137.890 154.845 ;
        RECT 135.930 153.945 136.155 154.075 ;
        RECT 136.325 154.005 136.850 154.225 ;
        RECT 137.020 154.585 137.890 154.755 ;
        RECT 135.565 153.355 135.815 153.815 ;
        RECT 135.985 153.805 136.155 153.945 ;
        RECT 137.020 153.805 137.190 154.585 ;
        RECT 137.720 154.515 137.890 154.585 ;
        RECT 137.400 154.335 137.600 154.365 ;
        RECT 138.060 154.335 138.230 155.405 ;
        RECT 138.400 154.515 138.590 155.235 ;
        RECT 137.400 154.035 138.230 154.335 ;
        RECT 138.760 154.305 139.080 155.265 ;
        RECT 135.985 153.635 136.320 153.805 ;
        RECT 136.515 153.635 137.190 153.805 ;
        RECT 137.510 153.355 137.880 153.855 ;
        RECT 138.060 153.805 138.230 154.035 ;
        RECT 138.615 153.975 139.080 154.305 ;
        RECT 139.250 154.595 139.420 155.435 ;
        RECT 139.600 155.405 139.915 155.905 ;
        RECT 140.145 155.175 140.485 155.735 ;
        RECT 139.590 154.800 140.485 155.175 ;
        RECT 140.655 154.895 140.825 155.905 ;
        RECT 140.295 154.595 140.485 154.800 ;
        RECT 140.995 154.845 141.325 155.690 ;
        RECT 142.130 155.275 142.415 155.735 ;
        RECT 142.585 155.445 142.855 155.905 ;
        RECT 142.130 155.055 143.085 155.275 ;
        RECT 140.995 154.765 141.385 154.845 ;
        RECT 141.170 154.715 141.385 154.765 ;
        RECT 139.250 154.265 140.125 154.595 ;
        RECT 140.295 154.265 141.045 154.595 ;
        RECT 139.250 153.805 139.420 154.265 ;
        RECT 140.295 154.095 140.495 154.265 ;
        RECT 141.215 154.135 141.385 154.715 ;
        RECT 142.015 154.325 142.705 154.885 ;
        RECT 142.875 154.155 143.085 155.055 ;
        RECT 141.160 154.095 141.385 154.135 ;
        RECT 138.060 153.635 138.465 153.805 ;
        RECT 138.635 153.635 139.420 153.805 ;
        RECT 139.695 153.355 139.905 153.885 ;
        RECT 140.165 153.570 140.495 154.095 ;
        RECT 141.005 154.010 141.385 154.095 ;
        RECT 140.665 153.355 140.835 153.965 ;
        RECT 141.005 153.575 141.335 154.010 ;
        RECT 142.130 153.985 143.085 154.155 ;
        RECT 143.255 154.885 143.655 155.735 ;
        RECT 143.845 155.275 144.125 155.735 ;
        RECT 144.645 155.445 144.970 155.905 ;
        RECT 143.845 155.055 144.970 155.275 ;
        RECT 143.255 154.325 144.350 154.885 ;
        RECT 144.520 154.595 144.970 155.055 ;
        RECT 145.140 154.765 145.525 155.735 ;
        RECT 142.130 153.525 142.415 153.985 ;
        RECT 142.585 153.355 142.855 153.815 ;
        RECT 143.255 153.525 143.655 154.325 ;
        RECT 144.520 154.265 145.075 154.595 ;
        RECT 144.520 154.155 144.970 154.265 ;
        RECT 143.845 153.985 144.970 154.155 ;
        RECT 145.245 154.095 145.525 154.765 ;
        RECT 145.695 154.815 146.905 155.905 ;
        RECT 145.695 154.275 146.215 154.815 ;
        RECT 146.385 154.105 146.905 154.645 ;
        RECT 143.845 153.525 144.125 153.985 ;
        RECT 144.645 153.355 144.970 153.815 ;
        RECT 145.140 153.525 145.525 154.095 ;
        RECT 145.695 153.355 146.905 154.105 ;
        RECT 17.270 153.185 146.990 153.355 ;
        RECT 17.355 152.435 18.565 153.185 ;
        RECT 18.735 152.640 24.080 153.185 ;
        RECT 24.255 152.640 29.600 153.185 ;
        RECT 17.355 151.895 17.875 152.435 ;
        RECT 18.045 151.725 18.565 152.265 ;
        RECT 20.320 151.810 20.660 152.640 ;
        RECT 17.355 150.635 18.565 151.725 ;
        RECT 22.140 151.070 22.490 152.320 ;
        RECT 25.840 151.810 26.180 152.640 ;
        RECT 29.775 152.415 31.445 153.185 ;
        RECT 32.080 152.680 32.415 153.185 ;
        RECT 32.585 152.615 32.825 152.990 ;
        RECT 33.105 152.855 33.275 153.000 ;
        RECT 33.105 152.660 33.480 152.855 ;
        RECT 33.840 152.690 34.235 153.185 ;
        RECT 27.660 151.070 28.010 152.320 ;
        RECT 29.775 151.895 30.525 152.415 ;
        RECT 30.695 151.725 31.445 152.245 ;
        RECT 18.735 150.635 24.080 151.070 ;
        RECT 24.255 150.635 29.600 151.070 ;
        RECT 29.775 150.635 31.445 151.725 ;
        RECT 32.135 151.655 32.435 152.505 ;
        RECT 32.605 152.465 32.825 152.615 ;
        RECT 32.605 152.135 33.140 152.465 ;
        RECT 33.310 152.325 33.480 152.660 ;
        RECT 34.405 152.495 34.645 153.015 ;
        RECT 32.605 151.485 32.840 152.135 ;
        RECT 33.310 151.965 34.295 152.325 ;
        RECT 32.165 151.255 32.840 151.485 ;
        RECT 33.010 151.945 34.295 151.965 ;
        RECT 33.010 151.795 33.870 151.945 ;
        RECT 32.165 150.825 32.335 151.255 ;
        RECT 32.505 150.635 32.835 151.085 ;
        RECT 33.010 150.850 33.295 151.795 ;
        RECT 34.470 151.690 34.645 152.495 ;
        RECT 35.775 152.455 36.065 153.185 ;
        RECT 35.765 151.945 36.065 152.275 ;
        RECT 36.245 152.255 36.475 152.895 ;
        RECT 36.655 152.635 36.965 153.005 ;
        RECT 37.145 152.815 37.815 153.185 ;
        RECT 36.655 152.435 37.885 152.635 ;
        RECT 36.245 151.945 36.770 152.255 ;
        RECT 36.950 151.945 37.415 152.255 ;
        RECT 37.595 151.765 37.885 152.435 ;
        RECT 33.470 151.315 34.165 151.625 ;
        RECT 33.475 150.635 34.160 151.105 ;
        RECT 34.340 150.905 34.645 151.690 ;
        RECT 35.775 151.525 36.935 151.765 ;
        RECT 35.775 150.815 36.035 151.525 ;
        RECT 36.205 150.635 36.535 151.345 ;
        RECT 36.705 150.815 36.935 151.525 ;
        RECT 37.115 151.545 37.885 151.765 ;
        RECT 37.115 150.815 37.385 151.545 ;
        RECT 37.565 150.635 37.905 151.365 ;
        RECT 38.075 150.815 38.335 153.005 ;
        RECT 38.515 152.465 38.855 152.975 ;
        RECT 38.515 151.065 38.775 152.465 ;
        RECT 39.025 152.385 39.295 153.185 ;
        RECT 38.950 151.945 39.280 152.195 ;
        RECT 39.475 151.945 39.755 152.915 ;
        RECT 39.935 151.945 40.235 152.915 ;
        RECT 40.415 151.945 40.765 152.910 ;
        RECT 40.985 152.685 41.480 153.015 ;
        RECT 38.965 151.775 39.280 151.945 ;
        RECT 40.985 151.775 41.155 152.685 ;
        RECT 38.965 151.605 41.155 151.775 ;
        RECT 38.515 150.805 38.855 151.065 ;
        RECT 39.025 150.635 39.355 151.435 ;
        RECT 39.820 150.805 40.070 151.605 ;
        RECT 40.255 150.635 40.585 151.355 ;
        RECT 40.805 150.805 41.055 151.605 ;
        RECT 41.325 151.195 41.565 152.505 ;
        RECT 41.735 152.435 42.945 153.185 ;
        RECT 43.115 152.460 43.405 153.185 ;
        RECT 43.575 152.640 48.920 153.185 ;
        RECT 49.095 152.640 54.440 153.185 ;
        RECT 41.735 151.895 42.255 152.435 ;
        RECT 42.425 151.725 42.945 152.265 ;
        RECT 45.160 151.810 45.500 152.640 ;
        RECT 41.225 150.635 41.560 151.015 ;
        RECT 41.735 150.635 42.945 151.725 ;
        RECT 43.115 150.635 43.405 151.800 ;
        RECT 46.980 151.070 47.330 152.320 ;
        RECT 50.680 151.810 51.020 152.640 ;
        RECT 54.615 152.385 55.310 153.015 ;
        RECT 55.515 152.385 55.825 153.185 ;
        RECT 52.500 151.070 52.850 152.320 ;
        RECT 54.635 151.945 54.970 152.195 ;
        RECT 55.140 151.785 55.310 152.385 ;
        RECT 56.455 152.365 56.715 153.185 ;
        RECT 56.885 152.365 57.215 152.785 ;
        RECT 57.395 152.700 58.185 152.965 ;
        RECT 56.965 152.275 57.215 152.365 ;
        RECT 55.480 151.945 55.815 152.215 ;
        RECT 43.575 150.635 48.920 151.070 ;
        RECT 49.095 150.635 54.440 151.070 ;
        RECT 54.615 150.635 54.875 151.775 ;
        RECT 55.045 150.805 55.375 151.785 ;
        RECT 55.545 150.635 55.825 151.775 ;
        RECT 56.455 151.315 56.795 152.195 ;
        RECT 56.965 152.025 57.760 152.275 ;
        RECT 56.455 150.635 56.715 151.145 ;
        RECT 56.965 150.805 57.135 152.025 ;
        RECT 57.930 151.845 58.185 152.700 ;
        RECT 58.355 152.545 58.555 152.965 ;
        RECT 58.745 152.725 59.075 153.185 ;
        RECT 58.355 152.025 58.765 152.545 ;
        RECT 59.245 152.535 59.505 153.015 ;
        RECT 58.935 151.845 59.165 152.275 ;
        RECT 57.375 151.675 59.165 151.845 ;
        RECT 57.375 151.310 57.625 151.675 ;
        RECT 57.795 151.315 58.125 151.505 ;
        RECT 58.345 151.380 59.060 151.675 ;
        RECT 59.335 151.505 59.505 152.535 ;
        RECT 60.225 152.635 60.395 152.925 ;
        RECT 60.565 152.805 60.895 153.185 ;
        RECT 60.225 152.465 60.890 152.635 ;
        RECT 60.140 151.645 60.490 152.295 ;
        RECT 57.795 151.140 57.990 151.315 ;
        RECT 57.375 150.635 57.990 151.140 ;
        RECT 58.160 150.805 58.635 151.145 ;
        RECT 58.805 150.635 59.020 151.180 ;
        RECT 59.230 150.805 59.505 151.505 ;
        RECT 60.660 151.475 60.890 152.465 ;
        RECT 60.225 151.305 60.890 151.475 ;
        RECT 60.225 150.805 60.395 151.305 ;
        RECT 60.565 150.635 60.895 151.135 ;
        RECT 61.065 150.805 61.250 152.925 ;
        RECT 61.505 152.725 61.755 153.185 ;
        RECT 61.925 152.735 62.260 152.905 ;
        RECT 62.455 152.735 63.130 152.905 ;
        RECT 61.925 152.595 62.095 152.735 ;
        RECT 61.420 151.605 61.700 152.555 ;
        RECT 61.870 152.465 62.095 152.595 ;
        RECT 61.870 151.360 62.040 152.465 ;
        RECT 62.265 152.315 62.790 152.535 ;
        RECT 62.210 151.550 62.450 152.145 ;
        RECT 62.620 151.615 62.790 152.315 ;
        RECT 62.960 151.955 63.130 152.735 ;
        RECT 63.450 152.685 63.820 153.185 ;
        RECT 64.000 152.735 64.405 152.905 ;
        RECT 64.575 152.735 65.360 152.905 ;
        RECT 64.000 152.505 64.170 152.735 ;
        RECT 63.340 152.205 64.170 152.505 ;
        RECT 64.555 152.235 65.020 152.565 ;
        RECT 63.340 152.175 63.540 152.205 ;
        RECT 63.660 151.955 63.830 152.025 ;
        RECT 62.960 151.785 63.830 151.955 ;
        RECT 63.320 151.695 63.830 151.785 ;
        RECT 61.870 151.230 62.175 151.360 ;
        RECT 62.620 151.250 63.150 151.615 ;
        RECT 61.490 150.635 61.755 151.095 ;
        RECT 61.925 150.805 62.175 151.230 ;
        RECT 63.320 151.080 63.490 151.695 ;
        RECT 62.385 150.910 63.490 151.080 ;
        RECT 63.660 150.635 63.830 151.435 ;
        RECT 64.000 151.135 64.170 152.205 ;
        RECT 64.340 151.305 64.530 152.025 ;
        RECT 64.700 151.275 65.020 152.235 ;
        RECT 65.190 152.275 65.360 152.735 ;
        RECT 65.635 152.655 65.845 153.185 ;
        RECT 66.105 152.445 66.435 152.970 ;
        RECT 66.605 152.575 66.775 153.185 ;
        RECT 66.945 152.530 67.275 152.965 ;
        RECT 66.945 152.445 67.325 152.530 ;
        RECT 66.235 152.275 66.435 152.445 ;
        RECT 67.100 152.405 67.325 152.445 ;
        RECT 65.190 151.945 66.065 152.275 ;
        RECT 66.235 151.945 66.985 152.275 ;
        RECT 64.000 150.805 64.250 151.135 ;
        RECT 65.190 151.105 65.360 151.945 ;
        RECT 66.235 151.740 66.425 151.945 ;
        RECT 67.155 151.825 67.325 152.405 ;
        RECT 67.495 152.435 68.705 153.185 ;
        RECT 68.875 152.460 69.165 153.185 ;
        RECT 67.495 151.895 68.015 152.435 ;
        RECT 69.335 152.415 71.925 153.185 ;
        RECT 67.110 151.775 67.325 151.825 ;
        RECT 65.530 151.365 66.425 151.740 ;
        RECT 66.935 151.695 67.325 151.775 ;
        RECT 68.185 151.725 68.705 152.265 ;
        RECT 69.335 151.895 70.545 152.415 ;
        RECT 72.095 152.385 72.405 153.185 ;
        RECT 72.610 152.385 73.305 153.015 ;
        RECT 64.475 150.935 65.360 151.105 ;
        RECT 65.540 150.635 65.855 151.135 ;
        RECT 66.085 150.805 66.425 151.365 ;
        RECT 66.595 150.635 66.765 151.645 ;
        RECT 66.935 150.850 67.265 151.695 ;
        RECT 67.495 150.635 68.705 151.725 ;
        RECT 68.875 150.635 69.165 151.800 ;
        RECT 70.715 151.725 71.925 152.245 ;
        RECT 72.105 151.945 72.440 152.215 ;
        RECT 72.610 151.825 72.780 152.385 ;
        RECT 73.475 152.240 73.815 153.015 ;
        RECT 73.985 152.725 74.155 153.185 ;
        RECT 74.395 152.750 74.755 153.015 ;
        RECT 74.395 152.745 74.750 152.750 ;
        RECT 74.395 152.735 74.745 152.745 ;
        RECT 74.395 152.730 74.740 152.735 ;
        RECT 74.395 152.720 74.735 152.730 ;
        RECT 75.385 152.725 75.555 153.185 ;
        RECT 74.395 152.715 74.730 152.720 ;
        RECT 74.395 152.705 74.720 152.715 ;
        RECT 74.395 152.695 74.710 152.705 ;
        RECT 74.395 152.555 74.695 152.695 ;
        RECT 73.985 152.365 74.695 152.555 ;
        RECT 74.885 152.555 75.215 152.635 ;
        RECT 75.725 152.555 76.065 153.015 ;
        RECT 74.885 152.365 76.065 152.555 ;
        RECT 76.700 152.445 76.955 153.015 ;
        RECT 77.125 152.785 77.455 153.185 ;
        RECT 77.880 152.650 78.410 153.015 ;
        RECT 78.600 152.845 78.875 153.015 ;
        RECT 78.595 152.675 78.875 152.845 ;
        RECT 77.880 152.615 78.055 152.650 ;
        RECT 77.125 152.445 78.055 152.615 ;
        RECT 72.950 151.945 73.285 152.195 ;
        RECT 72.610 151.785 72.785 151.825 ;
        RECT 69.335 150.635 71.925 151.725 ;
        RECT 72.095 150.635 72.375 151.775 ;
        RECT 72.545 150.805 72.875 151.785 ;
        RECT 73.045 150.635 73.305 151.775 ;
        RECT 73.475 150.805 73.755 152.240 ;
        RECT 73.985 151.795 74.270 152.365 ;
        RECT 74.455 151.965 74.925 152.195 ;
        RECT 75.095 152.175 75.425 152.195 ;
        RECT 75.095 151.995 75.545 152.175 ;
        RECT 75.735 151.995 76.065 152.195 ;
        RECT 73.985 151.580 75.135 151.795 ;
        RECT 73.925 150.635 74.635 151.410 ;
        RECT 74.805 150.805 75.135 151.580 ;
        RECT 75.330 150.880 75.545 151.995 ;
        RECT 75.835 151.655 76.065 151.995 ;
        RECT 76.700 151.775 76.870 152.445 ;
        RECT 77.125 152.275 77.295 152.445 ;
        RECT 77.040 151.945 77.295 152.275 ;
        RECT 77.520 151.945 77.715 152.275 ;
        RECT 75.725 150.635 76.055 151.355 ;
        RECT 76.700 150.805 77.035 151.775 ;
        RECT 77.205 150.635 77.375 151.775 ;
        RECT 77.545 150.975 77.715 151.945 ;
        RECT 77.885 151.315 78.055 152.445 ;
        RECT 78.225 151.655 78.395 152.455 ;
        RECT 78.600 151.855 78.875 152.675 ;
        RECT 79.045 151.655 79.235 153.015 ;
        RECT 79.415 152.650 79.925 153.185 ;
        RECT 80.145 152.375 80.390 152.980 ;
        RECT 81.465 152.670 81.635 153.185 ;
        RECT 81.805 152.530 82.135 152.965 ;
        RECT 82.305 152.575 82.475 153.185 ;
        RECT 81.755 152.445 82.135 152.530 ;
        RECT 82.645 152.445 82.975 152.970 ;
        RECT 83.235 152.655 83.445 153.185 ;
        RECT 83.720 152.735 84.505 152.905 ;
        RECT 84.675 152.735 85.080 152.905 ;
        RECT 81.755 152.405 81.980 152.445 ;
        RECT 79.435 152.205 80.665 152.375 ;
        RECT 78.225 151.485 79.235 151.655 ;
        RECT 79.405 151.640 80.155 151.830 ;
        RECT 77.885 151.145 79.010 151.315 ;
        RECT 79.405 150.975 79.575 151.640 ;
        RECT 80.325 151.395 80.665 152.205 ;
        RECT 81.755 151.825 81.925 152.405 ;
        RECT 82.645 152.275 82.845 152.445 ;
        RECT 83.720 152.275 83.890 152.735 ;
        RECT 82.095 151.945 82.845 152.275 ;
        RECT 83.015 151.945 83.890 152.275 ;
        RECT 81.755 151.775 81.970 151.825 ;
        RECT 81.755 151.695 82.145 151.775 ;
        RECT 77.545 150.805 79.575 150.975 ;
        RECT 79.745 150.635 79.915 151.395 ;
        RECT 80.150 150.985 80.665 151.395 ;
        RECT 81.475 150.635 81.645 151.550 ;
        RECT 81.815 150.850 82.145 151.695 ;
        RECT 82.655 151.740 82.845 151.945 ;
        RECT 82.315 150.635 82.485 151.645 ;
        RECT 82.655 151.365 83.550 151.740 ;
        RECT 82.655 150.805 82.995 151.365 ;
        RECT 83.225 150.635 83.540 151.135 ;
        RECT 83.720 151.105 83.890 151.945 ;
        RECT 84.060 152.235 84.525 152.565 ;
        RECT 84.910 152.505 85.080 152.735 ;
        RECT 85.260 152.685 85.630 153.185 ;
        RECT 85.950 152.735 86.625 152.905 ;
        RECT 86.820 152.735 87.155 152.905 ;
        RECT 84.060 151.275 84.380 152.235 ;
        RECT 84.910 152.205 85.740 152.505 ;
        RECT 84.550 151.305 84.740 152.025 ;
        RECT 84.910 151.135 85.080 152.205 ;
        RECT 85.540 152.175 85.740 152.205 ;
        RECT 85.250 151.955 85.420 152.025 ;
        RECT 85.950 151.955 86.120 152.735 ;
        RECT 86.985 152.595 87.155 152.735 ;
        RECT 87.325 152.725 87.575 153.185 ;
        RECT 85.250 151.785 86.120 151.955 ;
        RECT 86.290 152.315 86.815 152.535 ;
        RECT 86.985 152.465 87.210 152.595 ;
        RECT 85.250 151.695 85.760 151.785 ;
        RECT 83.720 150.935 84.605 151.105 ;
        RECT 84.830 150.805 85.080 151.135 ;
        RECT 85.250 150.635 85.420 151.435 ;
        RECT 85.590 151.080 85.760 151.695 ;
        RECT 86.290 151.615 86.460 152.315 ;
        RECT 85.930 151.250 86.460 151.615 ;
        RECT 86.630 151.550 86.870 152.145 ;
        RECT 87.040 151.360 87.210 152.465 ;
        RECT 87.380 151.605 87.660 152.555 ;
        RECT 86.905 151.230 87.210 151.360 ;
        RECT 85.590 150.910 86.695 151.080 ;
        RECT 86.905 150.805 87.155 151.230 ;
        RECT 87.325 150.635 87.590 151.095 ;
        RECT 87.830 150.805 88.015 152.925 ;
        RECT 88.185 152.805 88.515 153.185 ;
        RECT 88.685 152.635 88.855 152.925 ;
        RECT 88.190 152.465 88.855 152.635 ;
        RECT 88.190 151.475 88.420 152.465 ;
        RECT 89.115 152.415 91.705 153.185 ;
        RECT 88.590 151.645 88.940 152.295 ;
        RECT 89.115 151.895 90.325 152.415 ;
        RECT 90.495 151.725 91.705 152.245 ;
        RECT 88.190 151.305 88.855 151.475 ;
        RECT 88.185 150.635 88.515 151.135 ;
        RECT 88.685 150.805 88.855 151.305 ;
        RECT 89.115 150.635 91.705 151.725 ;
        RECT 91.875 152.240 92.215 153.015 ;
        RECT 92.385 152.725 92.555 153.185 ;
        RECT 92.795 152.750 93.155 153.015 ;
        RECT 92.795 152.745 93.150 152.750 ;
        RECT 92.795 152.735 93.145 152.745 ;
        RECT 92.795 152.730 93.140 152.735 ;
        RECT 92.795 152.720 93.135 152.730 ;
        RECT 93.785 152.725 93.955 153.185 ;
        RECT 92.795 152.715 93.130 152.720 ;
        RECT 92.795 152.705 93.120 152.715 ;
        RECT 92.795 152.695 93.110 152.705 ;
        RECT 92.795 152.555 93.095 152.695 ;
        RECT 92.385 152.365 93.095 152.555 ;
        RECT 93.285 152.555 93.615 152.635 ;
        RECT 94.125 152.555 94.465 153.015 ;
        RECT 93.285 152.365 94.465 152.555 ;
        RECT 94.635 152.460 94.925 153.185 ;
        RECT 95.095 152.445 95.480 153.015 ;
        RECT 95.650 152.725 95.975 153.185 ;
        RECT 96.495 152.555 96.775 153.015 ;
        RECT 91.875 150.805 92.155 152.240 ;
        RECT 92.385 151.795 92.670 152.365 ;
        RECT 92.855 151.965 93.325 152.195 ;
        RECT 93.495 152.175 93.825 152.195 ;
        RECT 93.495 151.995 93.945 152.175 ;
        RECT 94.135 151.995 94.465 152.195 ;
        RECT 92.385 151.580 93.535 151.795 ;
        RECT 92.325 150.635 93.035 151.410 ;
        RECT 93.205 150.805 93.535 151.580 ;
        RECT 93.730 150.880 93.945 151.995 ;
        RECT 94.235 151.655 94.465 151.995 ;
        RECT 94.125 150.635 94.455 151.355 ;
        RECT 94.635 150.635 94.925 151.800 ;
        RECT 95.095 151.775 95.375 152.445 ;
        RECT 95.650 152.385 96.775 152.555 ;
        RECT 95.650 152.275 96.100 152.385 ;
        RECT 95.545 151.945 96.100 152.275 ;
        RECT 96.965 152.215 97.365 153.015 ;
        RECT 97.765 152.725 98.035 153.185 ;
        RECT 98.205 152.555 98.490 153.015 ;
        RECT 95.095 150.805 95.480 151.775 ;
        RECT 95.650 151.485 96.100 151.945 ;
        RECT 96.270 151.655 97.365 152.215 ;
        RECT 95.650 151.265 96.775 151.485 ;
        RECT 95.650 150.635 95.975 151.095 ;
        RECT 96.495 150.805 96.775 151.265 ;
        RECT 96.965 150.805 97.365 151.655 ;
        RECT 97.535 152.385 98.490 152.555 ;
        RECT 98.775 152.435 99.985 153.185 ;
        RECT 100.270 152.555 100.555 153.015 ;
        RECT 100.725 152.725 100.995 153.185 ;
        RECT 97.535 151.485 97.745 152.385 ;
        RECT 97.915 151.655 98.605 152.215 ;
        RECT 98.775 151.895 99.295 152.435 ;
        RECT 100.270 152.385 101.225 152.555 ;
        RECT 99.465 151.725 99.985 152.265 ;
        RECT 97.535 151.265 98.490 151.485 ;
        RECT 97.765 150.635 98.035 151.095 ;
        RECT 98.205 150.805 98.490 151.265 ;
        RECT 98.775 150.635 99.985 151.725 ;
        RECT 100.155 151.655 100.845 152.215 ;
        RECT 101.015 151.485 101.225 152.385 ;
        RECT 100.270 151.265 101.225 151.485 ;
        RECT 101.395 152.215 101.795 153.015 ;
        RECT 101.985 152.555 102.265 153.015 ;
        RECT 102.785 152.725 103.110 153.185 ;
        RECT 101.985 152.385 103.110 152.555 ;
        RECT 103.280 152.445 103.665 153.015 ;
        RECT 102.660 152.275 103.110 152.385 ;
        RECT 101.395 151.655 102.490 152.215 ;
        RECT 102.660 151.945 103.215 152.275 ;
        RECT 100.270 150.805 100.555 151.265 ;
        RECT 100.725 150.635 100.995 151.095 ;
        RECT 101.395 150.805 101.795 151.655 ;
        RECT 102.660 151.485 103.110 151.945 ;
        RECT 103.385 151.775 103.665 152.445 ;
        RECT 101.985 151.265 103.110 151.485 ;
        RECT 101.985 150.805 102.265 151.265 ;
        RECT 102.785 150.635 103.110 151.095 ;
        RECT 103.280 150.805 103.665 151.775 ;
        RECT 103.835 152.240 104.175 153.015 ;
        RECT 104.345 152.725 104.515 153.185 ;
        RECT 104.755 152.750 105.115 153.015 ;
        RECT 104.755 152.745 105.110 152.750 ;
        RECT 104.755 152.735 105.105 152.745 ;
        RECT 104.755 152.730 105.100 152.735 ;
        RECT 104.755 152.720 105.095 152.730 ;
        RECT 105.745 152.725 105.915 153.185 ;
        RECT 104.755 152.715 105.090 152.720 ;
        RECT 104.755 152.705 105.080 152.715 ;
        RECT 104.755 152.695 105.070 152.705 ;
        RECT 104.755 152.555 105.055 152.695 ;
        RECT 104.345 152.365 105.055 152.555 ;
        RECT 105.245 152.555 105.575 152.635 ;
        RECT 106.085 152.555 106.425 153.015 ;
        RECT 106.595 152.640 111.940 153.185 ;
        RECT 105.245 152.365 106.425 152.555 ;
        RECT 103.835 150.805 104.115 152.240 ;
        RECT 104.345 151.795 104.630 152.365 ;
        RECT 104.815 151.965 105.285 152.195 ;
        RECT 105.455 152.175 105.785 152.195 ;
        RECT 105.455 151.995 105.905 152.175 ;
        RECT 106.095 151.995 106.425 152.195 ;
        RECT 104.345 151.580 105.495 151.795 ;
        RECT 104.285 150.635 104.995 151.410 ;
        RECT 105.165 150.805 105.495 151.580 ;
        RECT 105.690 150.880 105.905 151.995 ;
        RECT 106.195 151.655 106.425 151.995 ;
        RECT 108.180 151.810 108.520 152.640 ;
        RECT 112.205 152.635 112.375 152.925 ;
        RECT 112.545 152.805 112.875 153.185 ;
        RECT 112.205 152.465 112.870 152.635 ;
        RECT 106.085 150.635 106.415 151.355 ;
        RECT 110.000 151.070 110.350 152.320 ;
        RECT 112.120 151.645 112.470 152.295 ;
        RECT 112.640 151.475 112.870 152.465 ;
        RECT 112.205 151.305 112.870 151.475 ;
        RECT 106.595 150.635 111.940 151.070 ;
        RECT 112.205 150.805 112.375 151.305 ;
        RECT 112.545 150.635 112.875 151.135 ;
        RECT 113.045 150.805 113.230 152.925 ;
        RECT 113.485 152.725 113.735 153.185 ;
        RECT 113.905 152.735 114.240 152.905 ;
        RECT 114.435 152.735 115.110 152.905 ;
        RECT 113.905 152.595 114.075 152.735 ;
        RECT 113.400 151.605 113.680 152.555 ;
        RECT 113.850 152.465 114.075 152.595 ;
        RECT 113.850 151.360 114.020 152.465 ;
        RECT 114.245 152.315 114.770 152.535 ;
        RECT 114.190 151.550 114.430 152.145 ;
        RECT 114.600 151.615 114.770 152.315 ;
        RECT 114.940 151.955 115.110 152.735 ;
        RECT 115.430 152.685 115.800 153.185 ;
        RECT 115.980 152.735 116.385 152.905 ;
        RECT 116.555 152.735 117.340 152.905 ;
        RECT 115.980 152.505 116.150 152.735 ;
        RECT 115.320 152.205 116.150 152.505 ;
        RECT 116.535 152.235 117.000 152.565 ;
        RECT 115.320 152.175 115.520 152.205 ;
        RECT 115.640 151.955 115.810 152.025 ;
        RECT 114.940 151.785 115.810 151.955 ;
        RECT 115.300 151.695 115.810 151.785 ;
        RECT 113.850 151.230 114.155 151.360 ;
        RECT 114.600 151.250 115.130 151.615 ;
        RECT 113.470 150.635 113.735 151.095 ;
        RECT 113.905 150.805 114.155 151.230 ;
        RECT 115.300 151.080 115.470 151.695 ;
        RECT 114.365 150.910 115.470 151.080 ;
        RECT 115.640 150.635 115.810 151.435 ;
        RECT 115.980 151.135 116.150 152.205 ;
        RECT 116.320 151.305 116.510 152.025 ;
        RECT 116.680 151.275 117.000 152.235 ;
        RECT 117.170 152.275 117.340 152.735 ;
        RECT 117.615 152.655 117.825 153.185 ;
        RECT 118.085 152.445 118.415 152.970 ;
        RECT 118.585 152.575 118.755 153.185 ;
        RECT 118.925 152.530 119.255 152.965 ;
        RECT 118.925 152.445 119.305 152.530 ;
        RECT 120.395 152.460 120.685 153.185 ;
        RECT 118.215 152.275 118.415 152.445 ;
        RECT 119.080 152.405 119.305 152.445 ;
        RECT 120.860 152.420 121.315 153.185 ;
        RECT 121.590 152.805 122.890 153.015 ;
        RECT 123.145 152.825 123.475 153.185 ;
        RECT 122.720 152.655 122.890 152.805 ;
        RECT 123.645 152.685 123.905 153.015 ;
        RECT 123.675 152.675 123.905 152.685 ;
        RECT 117.170 151.945 118.045 152.275 ;
        RECT 118.215 151.945 118.965 152.275 ;
        RECT 115.980 150.805 116.230 151.135 ;
        RECT 117.170 151.105 117.340 151.945 ;
        RECT 118.215 151.740 118.405 151.945 ;
        RECT 119.135 151.825 119.305 152.405 ;
        RECT 121.790 152.195 122.010 152.595 ;
        RECT 120.855 151.995 121.345 152.195 ;
        RECT 121.535 151.985 122.010 152.195 ;
        RECT 122.255 152.195 122.465 152.595 ;
        RECT 122.720 152.530 123.475 152.655 ;
        RECT 122.720 152.485 123.565 152.530 ;
        RECT 123.295 152.365 123.565 152.485 ;
        RECT 122.255 151.985 122.585 152.195 ;
        RECT 122.755 151.925 123.165 152.230 ;
        RECT 119.090 151.775 119.305 151.825 ;
        RECT 117.510 151.365 118.405 151.740 ;
        RECT 118.915 151.695 119.305 151.775 ;
        RECT 116.455 150.935 117.340 151.105 ;
        RECT 117.520 150.635 117.835 151.135 ;
        RECT 118.065 150.805 118.405 151.365 ;
        RECT 118.575 150.635 118.745 151.645 ;
        RECT 118.915 150.850 119.245 151.695 ;
        RECT 120.395 150.635 120.685 151.800 ;
        RECT 120.860 151.755 122.035 151.815 ;
        RECT 123.395 151.790 123.565 152.365 ;
        RECT 123.365 151.755 123.565 151.790 ;
        RECT 120.860 151.645 123.565 151.755 ;
        RECT 120.860 151.025 121.115 151.645 ;
        RECT 121.705 151.585 123.505 151.645 ;
        RECT 121.705 151.555 122.035 151.585 ;
        RECT 123.735 151.485 123.905 152.675 ;
        RECT 124.165 152.635 124.335 152.925 ;
        RECT 124.505 152.805 124.835 153.185 ;
        RECT 124.165 152.465 124.830 152.635 ;
        RECT 124.080 151.645 124.430 152.295 ;
        RECT 121.365 151.385 121.550 151.475 ;
        RECT 122.140 151.385 122.975 151.395 ;
        RECT 121.365 151.185 122.975 151.385 ;
        RECT 121.365 151.145 121.595 151.185 ;
        RECT 120.860 150.805 121.195 151.025 ;
        RECT 122.200 150.635 122.555 151.015 ;
        RECT 122.725 150.805 122.975 151.185 ;
        RECT 123.225 150.635 123.475 151.415 ;
        RECT 123.645 150.805 123.905 151.485 ;
        RECT 124.600 151.475 124.830 152.465 ;
        RECT 124.165 151.305 124.830 151.475 ;
        RECT 124.165 150.805 124.335 151.305 ;
        RECT 124.505 150.635 124.835 151.135 ;
        RECT 125.005 150.805 125.190 152.925 ;
        RECT 125.445 152.725 125.695 153.185 ;
        RECT 125.865 152.735 126.200 152.905 ;
        RECT 126.395 152.735 127.070 152.905 ;
        RECT 125.865 152.595 126.035 152.735 ;
        RECT 125.360 151.605 125.640 152.555 ;
        RECT 125.810 152.465 126.035 152.595 ;
        RECT 125.810 151.360 125.980 152.465 ;
        RECT 126.205 152.315 126.730 152.535 ;
        RECT 126.150 151.550 126.390 152.145 ;
        RECT 126.560 151.615 126.730 152.315 ;
        RECT 126.900 151.955 127.070 152.735 ;
        RECT 127.390 152.685 127.760 153.185 ;
        RECT 127.940 152.735 128.345 152.905 ;
        RECT 128.515 152.735 129.300 152.905 ;
        RECT 127.940 152.505 128.110 152.735 ;
        RECT 127.280 152.205 128.110 152.505 ;
        RECT 128.495 152.235 128.960 152.565 ;
        RECT 127.280 152.175 127.480 152.205 ;
        RECT 127.600 151.955 127.770 152.025 ;
        RECT 126.900 151.785 127.770 151.955 ;
        RECT 127.260 151.695 127.770 151.785 ;
        RECT 125.810 151.230 126.115 151.360 ;
        RECT 126.560 151.250 127.090 151.615 ;
        RECT 125.430 150.635 125.695 151.095 ;
        RECT 125.865 150.805 126.115 151.230 ;
        RECT 127.260 151.080 127.430 151.695 ;
        RECT 126.325 150.910 127.430 151.080 ;
        RECT 127.600 150.635 127.770 151.435 ;
        RECT 127.940 151.135 128.110 152.205 ;
        RECT 128.280 151.305 128.470 152.025 ;
        RECT 128.640 151.275 128.960 152.235 ;
        RECT 129.130 152.275 129.300 152.735 ;
        RECT 129.575 152.655 129.785 153.185 ;
        RECT 130.045 152.445 130.375 152.970 ;
        RECT 130.545 152.575 130.715 153.185 ;
        RECT 130.885 152.530 131.215 152.965 ;
        RECT 131.435 152.640 136.780 153.185 ;
        RECT 130.885 152.445 131.265 152.530 ;
        RECT 130.175 152.275 130.375 152.445 ;
        RECT 131.040 152.405 131.265 152.445 ;
        RECT 129.130 151.945 130.005 152.275 ;
        RECT 130.175 151.945 130.925 152.275 ;
        RECT 127.940 150.805 128.190 151.135 ;
        RECT 129.130 151.105 129.300 151.945 ;
        RECT 130.175 151.740 130.365 151.945 ;
        RECT 131.095 151.825 131.265 152.405 ;
        RECT 131.050 151.775 131.265 151.825 ;
        RECT 133.020 151.810 133.360 152.640 ;
        RECT 137.505 152.635 137.675 153.015 ;
        RECT 137.855 152.805 138.185 153.185 ;
        RECT 137.505 152.465 138.170 152.635 ;
        RECT 138.365 152.510 138.625 153.015 ;
        RECT 129.470 151.365 130.365 151.740 ;
        RECT 130.875 151.695 131.265 151.775 ;
        RECT 128.415 150.935 129.300 151.105 ;
        RECT 129.480 150.635 129.795 151.135 ;
        RECT 130.025 150.805 130.365 151.365 ;
        RECT 130.535 150.635 130.705 151.645 ;
        RECT 130.875 150.850 131.205 151.695 ;
        RECT 134.840 151.070 135.190 152.320 ;
        RECT 137.435 151.915 137.765 152.285 ;
        RECT 138.000 152.210 138.170 152.465 ;
        RECT 138.000 151.880 138.285 152.210 ;
        RECT 138.000 151.735 138.170 151.880 ;
        RECT 137.505 151.565 138.170 151.735 ;
        RECT 138.455 151.710 138.625 152.510 ;
        RECT 131.435 150.635 136.780 151.070 ;
        RECT 137.505 150.805 137.675 151.565 ;
        RECT 137.855 150.635 138.185 151.395 ;
        RECT 138.355 150.805 138.625 151.710 ;
        RECT 138.795 152.510 139.055 153.015 ;
        RECT 139.235 152.805 139.565 153.185 ;
        RECT 139.745 152.635 139.915 153.015 ;
        RECT 138.795 151.710 138.965 152.510 ;
        RECT 139.250 152.465 139.915 152.635 ;
        RECT 140.265 152.635 140.435 153.015 ;
        RECT 140.650 152.805 140.980 153.185 ;
        RECT 140.265 152.465 140.980 152.635 ;
        RECT 139.250 152.210 139.420 152.465 ;
        RECT 139.135 151.880 139.420 152.210 ;
        RECT 139.655 151.915 139.985 152.285 ;
        RECT 140.175 151.915 140.530 152.285 ;
        RECT 140.810 152.275 140.980 152.465 ;
        RECT 141.150 152.440 141.405 153.015 ;
        RECT 140.810 151.945 141.065 152.275 ;
        RECT 139.250 151.735 139.420 151.880 ;
        RECT 140.810 151.735 140.980 151.945 ;
        RECT 138.795 150.805 139.065 151.710 ;
        RECT 139.250 151.565 139.915 151.735 ;
        RECT 139.235 150.635 139.565 151.395 ;
        RECT 139.745 150.805 139.915 151.565 ;
        RECT 140.265 151.565 140.980 151.735 ;
        RECT 141.235 151.710 141.405 152.440 ;
        RECT 141.580 152.345 141.840 153.185 ;
        RECT 142.130 152.555 142.415 153.015 ;
        RECT 142.585 152.725 142.855 153.185 ;
        RECT 142.130 152.385 143.085 152.555 ;
        RECT 140.265 150.805 140.435 151.565 ;
        RECT 140.650 150.635 140.980 151.395 ;
        RECT 141.150 150.805 141.405 151.710 ;
        RECT 141.580 150.635 141.840 151.785 ;
        RECT 142.015 151.655 142.705 152.215 ;
        RECT 142.875 151.485 143.085 152.385 ;
        RECT 142.130 151.265 143.085 151.485 ;
        RECT 143.255 152.215 143.655 153.015 ;
        RECT 143.845 152.555 144.125 153.015 ;
        RECT 144.645 152.725 144.970 153.185 ;
        RECT 143.845 152.385 144.970 152.555 ;
        RECT 145.140 152.445 145.525 153.015 ;
        RECT 144.520 152.275 144.970 152.385 ;
        RECT 143.255 151.655 144.350 152.215 ;
        RECT 144.520 151.945 145.075 152.275 ;
        RECT 142.130 150.805 142.415 151.265 ;
        RECT 142.585 150.635 142.855 151.095 ;
        RECT 143.255 150.805 143.655 151.655 ;
        RECT 144.520 151.485 144.970 151.945 ;
        RECT 145.245 151.775 145.525 152.445 ;
        RECT 145.695 152.435 146.905 153.185 ;
        RECT 143.845 151.265 144.970 151.485 ;
        RECT 143.845 150.805 144.125 151.265 ;
        RECT 144.645 150.635 144.970 151.095 ;
        RECT 145.140 150.805 145.525 151.775 ;
        RECT 145.695 151.725 146.215 152.265 ;
        RECT 146.385 151.895 146.905 152.435 ;
        RECT 145.695 150.635 146.905 151.725 ;
        RECT 17.270 150.465 146.990 150.635 ;
        RECT 17.355 149.375 18.565 150.465 ;
        RECT 18.735 150.030 24.080 150.465 ;
        RECT 24.255 150.030 29.600 150.465 ;
        RECT 17.355 148.665 17.875 149.205 ;
        RECT 18.045 148.835 18.565 149.375 ;
        RECT 17.355 147.915 18.565 148.665 ;
        RECT 20.320 148.460 20.660 149.290 ;
        RECT 22.140 148.780 22.490 150.030 ;
        RECT 25.840 148.460 26.180 149.290 ;
        RECT 27.660 148.780 28.010 150.030 ;
        RECT 30.235 149.300 30.525 150.465 ;
        RECT 30.695 149.375 32.365 150.465 ;
        RECT 32.535 149.955 32.795 150.465 ;
        RECT 30.695 148.685 31.445 149.205 ;
        RECT 31.615 148.855 32.365 149.375 ;
        RECT 32.535 148.905 32.875 149.785 ;
        RECT 33.045 149.075 33.215 150.295 ;
        RECT 33.455 149.960 34.070 150.465 ;
        RECT 33.455 149.425 33.705 149.790 ;
        RECT 33.875 149.785 34.070 149.960 ;
        RECT 34.240 149.955 34.715 150.295 ;
        RECT 34.885 149.920 35.100 150.465 ;
        RECT 33.875 149.595 34.205 149.785 ;
        RECT 34.425 149.425 35.140 149.720 ;
        RECT 35.310 149.595 35.585 150.295 ;
        RECT 35.845 149.795 36.015 150.295 ;
        RECT 36.185 149.965 36.515 150.465 ;
        RECT 35.845 149.625 36.510 149.795 ;
        RECT 33.455 149.255 35.245 149.425 ;
        RECT 33.045 148.825 33.840 149.075 ;
        RECT 33.045 148.735 33.295 148.825 ;
        RECT 18.735 147.915 24.080 148.460 ;
        RECT 24.255 147.915 29.600 148.460 ;
        RECT 30.235 147.915 30.525 148.640 ;
        RECT 30.695 147.915 32.365 148.685 ;
        RECT 32.535 147.915 32.795 148.735 ;
        RECT 32.965 148.315 33.295 148.735 ;
        RECT 34.010 148.400 34.265 149.255 ;
        RECT 33.475 148.135 34.265 148.400 ;
        RECT 34.435 148.555 34.845 149.075 ;
        RECT 35.015 148.825 35.245 149.255 ;
        RECT 35.415 148.565 35.585 149.595 ;
        RECT 35.760 148.805 36.110 149.455 ;
        RECT 36.280 148.635 36.510 149.625 ;
        RECT 34.435 148.135 34.635 148.555 ;
        RECT 34.825 147.915 35.155 148.375 ;
        RECT 35.325 148.085 35.585 148.565 ;
        RECT 35.845 148.465 36.510 148.635 ;
        RECT 35.845 148.175 36.015 148.465 ;
        RECT 36.185 147.915 36.515 148.295 ;
        RECT 36.685 148.175 36.870 150.295 ;
        RECT 37.110 150.005 37.375 150.465 ;
        RECT 37.545 149.870 37.795 150.295 ;
        RECT 38.005 150.020 39.110 150.190 ;
        RECT 37.490 149.740 37.795 149.870 ;
        RECT 37.040 148.545 37.320 149.495 ;
        RECT 37.490 148.635 37.660 149.740 ;
        RECT 37.830 148.955 38.070 149.550 ;
        RECT 38.240 149.485 38.770 149.850 ;
        RECT 38.240 148.785 38.410 149.485 ;
        RECT 38.940 149.405 39.110 150.020 ;
        RECT 39.280 149.665 39.450 150.465 ;
        RECT 39.620 149.965 39.870 150.295 ;
        RECT 40.095 149.995 40.980 150.165 ;
        RECT 38.940 149.315 39.450 149.405 ;
        RECT 37.490 148.505 37.715 148.635 ;
        RECT 37.885 148.565 38.410 148.785 ;
        RECT 38.580 149.145 39.450 149.315 ;
        RECT 37.125 147.915 37.375 148.375 ;
        RECT 37.545 148.365 37.715 148.505 ;
        RECT 38.580 148.365 38.750 149.145 ;
        RECT 39.280 149.075 39.450 149.145 ;
        RECT 38.960 148.895 39.160 148.925 ;
        RECT 39.620 148.895 39.790 149.965 ;
        RECT 39.960 149.075 40.150 149.795 ;
        RECT 38.960 148.595 39.790 148.895 ;
        RECT 40.320 148.865 40.640 149.825 ;
        RECT 37.545 148.195 37.880 148.365 ;
        RECT 38.075 148.195 38.750 148.365 ;
        RECT 39.070 147.915 39.440 148.415 ;
        RECT 39.620 148.365 39.790 148.595 ;
        RECT 40.175 148.535 40.640 148.865 ;
        RECT 40.810 149.155 40.980 149.995 ;
        RECT 41.160 149.965 41.475 150.465 ;
        RECT 41.705 149.735 42.045 150.295 ;
        RECT 41.150 149.360 42.045 149.735 ;
        RECT 42.215 149.455 42.385 150.465 ;
        RECT 41.855 149.155 42.045 149.360 ;
        RECT 42.555 149.405 42.885 150.250 ;
        RECT 42.555 149.325 42.945 149.405 ;
        RECT 43.115 149.375 44.325 150.465 ;
        RECT 44.745 149.735 45.040 150.465 ;
        RECT 45.210 149.565 45.470 150.290 ;
        RECT 45.640 149.735 45.900 150.465 ;
        RECT 46.070 149.565 46.330 150.290 ;
        RECT 46.500 149.735 46.760 150.465 ;
        RECT 46.930 149.565 47.190 150.290 ;
        RECT 47.360 149.735 47.620 150.465 ;
        RECT 47.790 149.565 48.050 150.290 ;
        RECT 42.730 149.275 42.945 149.325 ;
        RECT 40.810 148.825 41.685 149.155 ;
        RECT 41.855 148.825 42.605 149.155 ;
        RECT 40.810 148.365 40.980 148.825 ;
        RECT 41.855 148.655 42.055 148.825 ;
        RECT 42.775 148.695 42.945 149.275 ;
        RECT 42.720 148.655 42.945 148.695 ;
        RECT 39.620 148.195 40.025 148.365 ;
        RECT 40.195 148.195 40.980 148.365 ;
        RECT 41.255 147.915 41.465 148.445 ;
        RECT 41.725 148.130 42.055 148.655 ;
        RECT 42.565 148.570 42.945 148.655 ;
        RECT 43.115 148.665 43.635 149.205 ;
        RECT 43.805 148.835 44.325 149.375 ;
        RECT 44.740 149.325 48.050 149.565 ;
        RECT 48.220 149.355 48.480 150.465 ;
        RECT 44.740 148.735 45.710 149.325 ;
        RECT 48.650 149.155 48.900 150.290 ;
        RECT 49.080 149.355 49.375 150.465 ;
        RECT 49.555 149.375 52.145 150.465 ;
        RECT 45.880 148.905 48.900 149.155 ;
        RECT 42.225 147.915 42.395 148.525 ;
        RECT 42.565 148.135 42.895 148.570 ;
        RECT 43.115 147.915 44.325 148.665 ;
        RECT 44.740 148.565 48.050 148.735 ;
        RECT 44.740 147.915 45.040 148.395 ;
        RECT 45.210 148.110 45.470 148.565 ;
        RECT 45.640 147.915 45.900 148.395 ;
        RECT 46.070 148.110 46.330 148.565 ;
        RECT 46.500 147.915 46.760 148.395 ;
        RECT 46.930 148.110 47.190 148.565 ;
        RECT 47.360 147.915 47.620 148.395 ;
        RECT 47.790 148.110 48.050 148.565 ;
        RECT 48.220 147.915 48.480 148.440 ;
        RECT 48.650 148.095 48.900 148.905 ;
        RECT 49.070 148.545 49.385 149.155 ;
        RECT 49.555 148.685 50.765 149.205 ;
        RECT 50.935 148.855 52.145 149.375 ;
        RECT 52.785 149.405 53.115 150.255 ;
        RECT 49.080 147.915 49.325 148.375 ;
        RECT 49.555 147.915 52.145 148.685 ;
        RECT 52.785 148.640 52.975 149.405 ;
        RECT 53.285 149.325 53.535 150.465 ;
        RECT 53.725 149.825 53.975 150.245 ;
        RECT 54.205 149.995 54.535 150.465 ;
        RECT 54.765 149.825 55.015 150.245 ;
        RECT 53.725 149.655 55.015 149.825 ;
        RECT 55.195 149.825 55.525 150.255 ;
        RECT 55.195 149.655 55.650 149.825 ;
        RECT 53.715 149.155 53.930 149.485 ;
        RECT 53.145 148.825 53.455 149.155 ;
        RECT 53.625 148.825 53.930 149.155 ;
        RECT 54.105 148.825 54.390 149.485 ;
        RECT 54.585 148.825 54.850 149.485 ;
        RECT 55.065 148.825 55.310 149.485 ;
        RECT 53.285 148.655 53.455 148.825 ;
        RECT 55.480 148.655 55.650 149.655 ;
        RECT 55.995 149.300 56.285 150.465 ;
        RECT 56.455 149.375 57.665 150.465 ;
        RECT 52.785 148.130 53.115 148.640 ;
        RECT 53.285 148.485 55.650 148.655 ;
        RECT 56.455 148.665 56.975 149.205 ;
        RECT 57.145 148.835 57.665 149.375 ;
        RECT 57.845 149.355 58.140 150.465 ;
        RECT 58.320 149.155 58.570 150.290 ;
        RECT 58.740 149.355 59.000 150.465 ;
        RECT 59.170 149.565 59.430 150.290 ;
        RECT 59.600 149.735 59.860 150.465 ;
        RECT 60.030 149.565 60.290 150.290 ;
        RECT 60.460 149.735 60.720 150.465 ;
        RECT 60.890 149.565 61.150 150.290 ;
        RECT 61.320 149.735 61.580 150.465 ;
        RECT 61.750 149.565 62.010 150.290 ;
        RECT 62.180 149.735 62.475 150.465 ;
        RECT 62.950 149.665 63.250 150.465 ;
        RECT 59.170 149.325 62.480 149.565 ;
        RECT 63.420 149.495 63.750 150.295 ;
        RECT 63.920 149.665 64.090 150.465 ;
        RECT 64.260 149.495 64.590 150.295 ;
        RECT 64.760 149.665 64.930 150.465 ;
        RECT 65.100 149.495 65.430 150.295 ;
        RECT 65.600 149.665 65.770 150.465 ;
        RECT 65.940 149.495 66.270 150.295 ;
        RECT 66.440 149.665 66.695 150.465 ;
        RECT 67.035 149.595 67.310 150.295 ;
        RECT 67.480 149.920 67.735 150.465 ;
        RECT 67.905 149.955 68.385 150.295 ;
        RECT 68.560 149.910 69.165 150.465 ;
        RECT 68.550 149.810 69.165 149.910 ;
        RECT 68.550 149.785 68.735 149.810 ;
        RECT 53.285 147.915 53.615 148.315 ;
        RECT 54.665 148.145 54.995 148.485 ;
        RECT 55.165 147.915 55.495 148.315 ;
        RECT 55.995 147.915 56.285 148.640 ;
        RECT 56.455 147.915 57.665 148.665 ;
        RECT 57.835 148.545 58.150 149.155 ;
        RECT 58.320 148.905 61.340 149.155 ;
        RECT 57.895 147.915 58.140 148.375 ;
        RECT 58.320 148.095 58.570 148.905 ;
        RECT 61.510 148.735 62.480 149.325 ;
        RECT 59.170 148.565 62.480 148.735 ;
        RECT 62.895 149.325 66.865 149.495 ;
        RECT 62.895 148.735 63.215 149.325 ;
        RECT 63.415 148.905 66.270 149.155 ;
        RECT 66.520 148.735 66.865 149.325 ;
        RECT 58.740 147.915 59.000 148.440 ;
        RECT 59.170 148.110 59.430 148.565 ;
        RECT 59.600 147.915 59.860 148.395 ;
        RECT 60.030 148.110 60.290 148.565 ;
        RECT 60.460 147.915 60.720 148.395 ;
        RECT 60.890 148.110 61.150 148.565 ;
        RECT 61.320 147.915 61.580 148.395 ;
        RECT 61.750 148.110 62.010 148.565 ;
        RECT 62.895 148.545 66.865 148.735 ;
        RECT 67.035 148.565 67.205 149.595 ;
        RECT 67.480 149.465 68.235 149.715 ;
        RECT 68.405 149.540 68.735 149.785 ;
        RECT 67.480 149.430 68.250 149.465 ;
        RECT 67.480 149.420 68.265 149.430 ;
        RECT 67.375 149.405 68.270 149.420 ;
        RECT 67.375 149.390 68.290 149.405 ;
        RECT 67.375 149.380 68.310 149.390 ;
        RECT 67.375 149.370 68.335 149.380 ;
        RECT 67.375 149.340 68.405 149.370 ;
        RECT 67.375 149.310 68.425 149.340 ;
        RECT 67.375 149.280 68.445 149.310 ;
        RECT 67.375 149.255 68.475 149.280 ;
        RECT 67.375 149.220 68.510 149.255 ;
        RECT 67.375 149.215 68.540 149.220 ;
        RECT 67.375 148.820 67.605 149.215 ;
        RECT 68.150 149.210 68.540 149.215 ;
        RECT 68.175 149.200 68.540 149.210 ;
        RECT 68.190 149.195 68.540 149.200 ;
        RECT 68.205 149.190 68.540 149.195 ;
        RECT 68.905 149.190 69.165 149.640 ;
        RECT 69.340 149.325 69.660 150.465 ;
        RECT 68.205 149.185 69.165 149.190 ;
        RECT 68.215 149.175 69.165 149.185 ;
        RECT 68.225 149.170 69.165 149.175 ;
        RECT 68.235 149.160 69.165 149.170 ;
        RECT 68.240 149.150 69.165 149.160 ;
        RECT 69.840 149.155 70.035 150.205 ;
        RECT 70.215 149.615 70.545 150.295 ;
        RECT 70.745 149.665 71.000 150.465 ;
        RECT 71.265 149.795 71.435 150.295 ;
        RECT 71.605 149.965 71.935 150.465 ;
        RECT 71.265 149.625 71.930 149.795 ;
        RECT 70.215 149.335 70.565 149.615 ;
        RECT 68.245 149.145 69.165 149.150 ;
        RECT 68.255 149.130 69.165 149.145 ;
        RECT 68.260 149.115 69.165 149.130 ;
        RECT 68.270 149.090 69.165 149.115 ;
        RECT 69.400 149.105 69.660 149.155 ;
        RECT 67.775 148.620 68.105 149.045 ;
        RECT 62.180 147.915 62.480 148.395 ;
        RECT 62.945 147.915 63.250 148.375 ;
        RECT 63.420 148.085 63.750 148.545 ;
        RECT 63.920 147.915 64.090 148.375 ;
        RECT 64.260 148.085 64.590 148.545 ;
        RECT 64.760 147.915 64.930 148.375 ;
        RECT 65.100 148.085 65.430 148.545 ;
        RECT 65.600 147.915 65.770 148.375 ;
        RECT 65.940 148.085 66.270 148.545 ;
        RECT 66.440 147.915 66.695 148.375 ;
        RECT 67.035 148.085 67.295 148.565 ;
        RECT 67.465 147.915 67.715 148.455 ;
        RECT 67.885 148.135 68.105 148.620 ;
        RECT 68.275 149.020 69.165 149.090 ;
        RECT 68.275 148.295 68.445 149.020 ;
        RECT 69.395 148.935 69.660 149.105 ;
        RECT 68.615 148.465 69.165 148.850 ;
        RECT 69.400 148.825 69.660 148.935 ;
        RECT 69.840 148.825 70.225 149.155 ;
        RECT 70.395 148.955 70.565 149.335 ;
        RECT 70.755 149.125 71.000 149.485 ;
        RECT 70.395 148.785 70.915 148.955 ;
        RECT 71.180 148.805 71.530 149.455 ;
        RECT 70.745 148.765 70.915 148.785 ;
        RECT 69.340 148.445 70.555 148.615 ;
        RECT 68.275 148.125 69.165 148.295 ;
        RECT 69.340 148.095 69.630 148.445 ;
        RECT 69.825 147.915 70.155 148.275 ;
        RECT 70.325 148.140 70.555 148.445 ;
        RECT 70.745 148.595 70.945 148.765 ;
        RECT 71.700 148.635 71.930 149.625 ;
        RECT 70.745 148.220 70.915 148.595 ;
        RECT 71.265 148.465 71.930 148.635 ;
        RECT 71.265 148.175 71.435 148.465 ;
        RECT 71.605 147.915 71.935 148.295 ;
        RECT 72.105 148.175 72.290 150.295 ;
        RECT 72.530 150.005 72.795 150.465 ;
        RECT 72.965 149.870 73.215 150.295 ;
        RECT 73.425 150.020 74.530 150.190 ;
        RECT 72.910 149.740 73.215 149.870 ;
        RECT 72.460 148.545 72.740 149.495 ;
        RECT 72.910 148.635 73.080 149.740 ;
        RECT 73.250 148.955 73.490 149.550 ;
        RECT 73.660 149.485 74.190 149.850 ;
        RECT 73.660 148.785 73.830 149.485 ;
        RECT 74.360 149.405 74.530 150.020 ;
        RECT 74.700 149.665 74.870 150.465 ;
        RECT 75.040 149.965 75.290 150.295 ;
        RECT 75.515 149.995 76.400 150.165 ;
        RECT 74.360 149.315 74.870 149.405 ;
        RECT 72.910 148.505 73.135 148.635 ;
        RECT 73.305 148.565 73.830 148.785 ;
        RECT 74.000 149.145 74.870 149.315 ;
        RECT 72.545 147.915 72.795 148.375 ;
        RECT 72.965 148.365 73.135 148.505 ;
        RECT 74.000 148.365 74.170 149.145 ;
        RECT 74.700 149.075 74.870 149.145 ;
        RECT 74.380 148.895 74.580 148.925 ;
        RECT 75.040 148.895 75.210 149.965 ;
        RECT 75.380 149.075 75.570 149.795 ;
        RECT 74.380 148.595 75.210 148.895 ;
        RECT 75.740 148.865 76.060 149.825 ;
        RECT 72.965 148.195 73.300 148.365 ;
        RECT 73.495 148.195 74.170 148.365 ;
        RECT 74.490 147.915 74.860 148.415 ;
        RECT 75.040 148.365 75.210 148.595 ;
        RECT 75.595 148.535 76.060 148.865 ;
        RECT 76.230 149.155 76.400 149.995 ;
        RECT 76.580 149.965 76.895 150.465 ;
        RECT 77.125 149.735 77.465 150.295 ;
        RECT 76.570 149.360 77.465 149.735 ;
        RECT 77.635 149.455 77.805 150.465 ;
        RECT 77.275 149.155 77.465 149.360 ;
        RECT 77.975 149.405 78.305 150.250 ;
        RECT 78.540 150.085 78.875 150.465 ;
        RECT 77.975 149.325 78.365 149.405 ;
        RECT 78.150 149.275 78.365 149.325 ;
        RECT 76.230 148.825 77.105 149.155 ;
        RECT 77.275 148.825 78.025 149.155 ;
        RECT 76.230 148.365 76.400 148.825 ;
        RECT 77.275 148.655 77.475 148.825 ;
        RECT 78.195 148.695 78.365 149.275 ;
        RECT 78.140 148.655 78.365 148.695 ;
        RECT 75.040 148.195 75.445 148.365 ;
        RECT 75.615 148.195 76.400 148.365 ;
        RECT 76.675 147.915 76.885 148.445 ;
        RECT 77.145 148.130 77.475 148.655 ;
        RECT 77.985 148.570 78.365 148.655 ;
        RECT 78.535 148.595 78.775 149.905 ;
        RECT 79.045 149.495 79.295 150.295 ;
        RECT 79.515 149.745 79.845 150.465 ;
        RECT 80.030 149.495 80.280 150.295 ;
        RECT 80.745 149.665 81.075 150.465 ;
        RECT 81.245 150.035 81.585 150.295 ;
        RECT 78.945 149.325 81.135 149.495 ;
        RECT 77.645 147.915 77.815 148.525 ;
        RECT 77.985 148.135 78.315 148.570 ;
        RECT 78.945 148.415 79.115 149.325 ;
        RECT 80.820 149.155 81.135 149.325 ;
        RECT 78.620 148.085 79.115 148.415 ;
        RECT 79.335 148.190 79.685 149.155 ;
        RECT 79.865 148.185 80.165 149.155 ;
        RECT 80.345 148.185 80.625 149.155 ;
        RECT 80.820 148.905 81.150 149.155 ;
        RECT 80.805 147.915 81.075 148.715 ;
        RECT 81.325 148.635 81.585 150.035 ;
        RECT 81.755 149.300 82.045 150.465 ;
        RECT 82.215 149.705 82.730 150.115 ;
        RECT 82.965 149.705 83.135 150.465 ;
        RECT 83.305 150.125 85.335 150.295 ;
        RECT 82.215 148.895 82.555 149.705 ;
        RECT 83.305 149.460 83.475 150.125 ;
        RECT 83.870 149.785 84.995 149.955 ;
        RECT 82.725 149.270 83.475 149.460 ;
        RECT 83.645 149.445 84.655 149.615 ;
        RECT 82.215 148.725 83.445 148.895 ;
        RECT 81.245 148.125 81.585 148.635 ;
        RECT 81.755 147.915 82.045 148.640 ;
        RECT 82.490 148.120 82.735 148.725 ;
        RECT 82.955 147.915 83.465 148.450 ;
        RECT 83.645 148.085 83.835 149.445 ;
        RECT 84.005 148.765 84.280 149.245 ;
        RECT 84.005 148.595 84.285 148.765 ;
        RECT 84.485 148.645 84.655 149.445 ;
        RECT 84.825 148.655 84.995 149.785 ;
        RECT 85.165 149.155 85.335 150.125 ;
        RECT 85.505 149.325 85.675 150.465 ;
        RECT 85.845 149.325 86.180 150.295 ;
        RECT 86.375 149.575 86.635 150.285 ;
        RECT 86.805 149.755 87.135 150.465 ;
        RECT 87.305 149.575 87.535 150.285 ;
        RECT 86.375 149.335 87.535 149.575 ;
        RECT 87.715 149.555 87.985 150.285 ;
        RECT 88.165 149.735 88.505 150.465 ;
        RECT 87.715 149.335 88.485 149.555 ;
        RECT 85.165 148.825 85.360 149.155 ;
        RECT 85.585 148.825 85.840 149.155 ;
        RECT 85.585 148.655 85.755 148.825 ;
        RECT 86.010 148.655 86.180 149.325 ;
        RECT 86.365 148.825 86.665 149.155 ;
        RECT 86.845 148.845 87.370 149.155 ;
        RECT 87.550 148.845 88.015 149.155 ;
        RECT 84.005 148.085 84.280 148.595 ;
        RECT 84.825 148.485 85.755 148.655 ;
        RECT 84.825 148.450 85.000 148.485 ;
        RECT 84.470 148.085 85.000 148.450 ;
        RECT 85.425 147.915 85.755 148.315 ;
        RECT 85.925 148.085 86.180 148.655 ;
        RECT 86.375 147.915 86.665 148.645 ;
        RECT 86.845 148.205 87.075 148.845 ;
        RECT 88.195 148.665 88.485 149.335 ;
        RECT 87.255 148.465 88.485 148.665 ;
        RECT 87.255 148.095 87.565 148.465 ;
        RECT 87.745 147.915 88.415 148.285 ;
        RECT 88.675 148.095 88.935 150.285 ;
        RECT 89.115 149.375 90.325 150.465 ;
        RECT 90.585 149.795 90.755 150.295 ;
        RECT 90.925 149.965 91.255 150.465 ;
        RECT 90.585 149.625 91.250 149.795 ;
        RECT 89.115 148.665 89.635 149.205 ;
        RECT 89.805 148.835 90.325 149.375 ;
        RECT 90.500 148.805 90.850 149.455 ;
        RECT 89.115 147.915 90.325 148.665 ;
        RECT 91.020 148.635 91.250 149.625 ;
        RECT 90.585 148.465 91.250 148.635 ;
        RECT 90.585 148.175 90.755 148.465 ;
        RECT 90.925 147.915 91.255 148.295 ;
        RECT 91.425 148.175 91.610 150.295 ;
        RECT 91.850 150.005 92.115 150.465 ;
        RECT 92.285 149.870 92.535 150.295 ;
        RECT 92.745 150.020 93.850 150.190 ;
        RECT 92.230 149.740 92.535 149.870 ;
        RECT 91.780 148.545 92.060 149.495 ;
        RECT 92.230 148.635 92.400 149.740 ;
        RECT 92.570 148.955 92.810 149.550 ;
        RECT 92.980 149.485 93.510 149.850 ;
        RECT 92.980 148.785 93.150 149.485 ;
        RECT 93.680 149.405 93.850 150.020 ;
        RECT 94.020 149.665 94.190 150.465 ;
        RECT 94.360 149.965 94.610 150.295 ;
        RECT 94.835 149.995 95.720 150.165 ;
        RECT 93.680 149.315 94.190 149.405 ;
        RECT 92.230 148.505 92.455 148.635 ;
        RECT 92.625 148.565 93.150 148.785 ;
        RECT 93.320 149.145 94.190 149.315 ;
        RECT 91.865 147.915 92.115 148.375 ;
        RECT 92.285 148.365 92.455 148.505 ;
        RECT 93.320 148.365 93.490 149.145 ;
        RECT 94.020 149.075 94.190 149.145 ;
        RECT 93.700 148.895 93.900 148.925 ;
        RECT 94.360 148.895 94.530 149.965 ;
        RECT 94.700 149.075 94.890 149.795 ;
        RECT 93.700 148.595 94.530 148.895 ;
        RECT 95.060 148.865 95.380 149.825 ;
        RECT 92.285 148.195 92.620 148.365 ;
        RECT 92.815 148.195 93.490 148.365 ;
        RECT 93.810 147.915 94.180 148.415 ;
        RECT 94.360 148.365 94.530 148.595 ;
        RECT 94.915 148.535 95.380 148.865 ;
        RECT 95.550 149.155 95.720 149.995 ;
        RECT 95.900 149.965 96.215 150.465 ;
        RECT 96.445 149.735 96.785 150.295 ;
        RECT 95.890 149.360 96.785 149.735 ;
        RECT 96.955 149.455 97.125 150.465 ;
        RECT 96.595 149.155 96.785 149.360 ;
        RECT 97.295 149.405 97.625 150.250 ;
        RECT 97.855 149.495 98.165 150.295 ;
        RECT 98.335 149.665 98.645 150.465 ;
        RECT 98.815 149.835 99.075 150.295 ;
        RECT 99.245 150.005 99.500 150.465 ;
        RECT 99.675 149.835 99.935 150.295 ;
        RECT 98.815 149.665 99.935 149.835 ;
        RECT 97.295 149.325 97.685 149.405 ;
        RECT 97.470 149.275 97.685 149.325 ;
        RECT 95.550 148.825 96.425 149.155 ;
        RECT 96.595 148.825 97.345 149.155 ;
        RECT 95.550 148.365 95.720 148.825 ;
        RECT 96.595 148.655 96.795 148.825 ;
        RECT 97.515 148.695 97.685 149.275 ;
        RECT 97.460 148.655 97.685 148.695 ;
        RECT 94.360 148.195 94.765 148.365 ;
        RECT 94.935 148.195 95.720 148.365 ;
        RECT 95.995 147.915 96.205 148.445 ;
        RECT 96.465 148.130 96.795 148.655 ;
        RECT 97.305 148.570 97.685 148.655 ;
        RECT 97.855 149.325 98.885 149.495 ;
        RECT 96.965 147.915 97.135 148.525 ;
        RECT 97.305 148.135 97.635 148.570 ;
        RECT 97.855 148.415 98.025 149.325 ;
        RECT 98.195 148.585 98.545 149.155 ;
        RECT 98.715 149.075 98.885 149.325 ;
        RECT 99.675 149.415 99.935 149.665 ;
        RECT 100.105 149.595 100.390 150.465 ;
        RECT 99.675 149.245 100.430 149.415 ;
        RECT 98.715 148.905 99.855 149.075 ;
        RECT 100.025 148.735 100.430 149.245 ;
        RECT 98.780 148.565 100.430 148.735 ;
        RECT 101.555 149.410 101.860 150.195 ;
        RECT 102.040 149.995 102.725 150.465 ;
        RECT 102.035 149.475 102.730 149.785 ;
        RECT 101.555 148.605 101.730 149.410 ;
        RECT 102.905 149.305 103.190 150.250 ;
        RECT 103.365 150.015 103.695 150.465 ;
        RECT 103.865 149.845 104.035 150.275 ;
        RECT 102.330 149.155 103.190 149.305 ;
        RECT 101.905 149.135 103.190 149.155 ;
        RECT 103.360 149.615 104.035 149.845 ;
        RECT 104.385 149.845 104.555 150.275 ;
        RECT 104.725 150.015 105.055 150.465 ;
        RECT 104.385 149.615 105.060 149.845 ;
        RECT 101.905 148.775 102.890 149.135 ;
        RECT 103.360 148.965 103.595 149.615 ;
        RECT 97.855 148.085 98.155 148.415 ;
        RECT 98.325 147.915 98.600 148.395 ;
        RECT 98.780 148.175 99.075 148.565 ;
        RECT 99.245 147.915 99.500 148.395 ;
        RECT 99.675 148.175 99.935 148.565 ;
        RECT 100.105 147.915 100.385 148.395 ;
        RECT 101.555 148.085 101.795 148.605 ;
        RECT 102.720 148.440 102.890 148.775 ;
        RECT 103.060 148.635 103.595 148.965 ;
        RECT 103.375 148.485 103.595 148.635 ;
        RECT 103.765 148.595 104.065 149.445 ;
        RECT 104.355 148.595 104.655 149.445 ;
        RECT 104.825 148.965 105.060 149.615 ;
        RECT 105.230 149.305 105.515 150.250 ;
        RECT 105.695 149.995 106.380 150.465 ;
        RECT 105.690 149.475 106.385 149.785 ;
        RECT 106.560 149.410 106.865 150.195 ;
        RECT 105.230 149.155 106.090 149.305 ;
        RECT 105.230 149.135 106.515 149.155 ;
        RECT 104.825 148.635 105.360 148.965 ;
        RECT 105.530 148.775 106.515 149.135 ;
        RECT 104.825 148.485 105.045 148.635 ;
        RECT 101.965 147.915 102.360 148.410 ;
        RECT 102.720 148.245 103.095 148.440 ;
        RECT 102.925 148.100 103.095 148.245 ;
        RECT 103.375 148.110 103.615 148.485 ;
        RECT 103.785 147.915 104.120 148.420 ;
        RECT 104.300 147.915 104.635 148.420 ;
        RECT 104.805 148.110 105.045 148.485 ;
        RECT 105.530 148.440 105.700 148.775 ;
        RECT 106.690 148.605 106.865 149.410 ;
        RECT 107.515 149.300 107.805 150.465 ;
        RECT 107.975 150.030 113.320 150.465 ;
        RECT 113.495 150.030 118.840 150.465 ;
        RECT 105.325 148.245 105.700 148.440 ;
        RECT 105.325 148.100 105.495 148.245 ;
        RECT 106.060 147.915 106.455 148.410 ;
        RECT 106.625 148.085 106.865 148.605 ;
        RECT 107.515 147.915 107.805 148.640 ;
        RECT 109.560 148.460 109.900 149.290 ;
        RECT 111.380 148.780 111.730 150.030 ;
        RECT 115.080 148.460 115.420 149.290 ;
        RECT 116.900 148.780 117.250 150.030 ;
        RECT 119.015 149.375 120.225 150.465 ;
        RECT 119.015 148.665 119.535 149.205 ;
        RECT 119.705 148.835 120.225 149.375 ;
        RECT 120.400 150.075 120.735 150.295 ;
        RECT 121.740 150.085 122.095 150.465 ;
        RECT 120.400 149.455 120.655 150.075 ;
        RECT 120.905 149.915 121.135 149.955 ;
        RECT 122.265 149.915 122.515 150.295 ;
        RECT 120.905 149.715 122.515 149.915 ;
        RECT 120.905 149.625 121.090 149.715 ;
        RECT 121.680 149.705 122.515 149.715 ;
        RECT 122.765 149.685 123.015 150.465 ;
        RECT 123.185 149.615 123.445 150.295 ;
        RECT 121.245 149.515 121.575 149.545 ;
        RECT 121.245 149.455 123.045 149.515 ;
        RECT 120.400 149.345 123.105 149.455 ;
        RECT 120.400 149.285 121.575 149.345 ;
        RECT 122.905 149.310 123.105 149.345 ;
        RECT 120.395 148.905 120.885 149.105 ;
        RECT 121.075 148.905 121.550 149.115 ;
        RECT 107.975 147.915 113.320 148.460 ;
        RECT 113.495 147.915 118.840 148.460 ;
        RECT 119.015 147.915 120.225 148.665 ;
        RECT 120.400 147.915 120.855 148.680 ;
        RECT 121.330 148.505 121.550 148.905 ;
        RECT 121.795 148.905 122.125 149.115 ;
        RECT 121.795 148.505 122.005 148.905 ;
        RECT 122.295 148.870 122.705 149.175 ;
        RECT 122.935 148.735 123.105 149.310 ;
        RECT 122.835 148.615 123.105 148.735 ;
        RECT 122.260 148.570 123.105 148.615 ;
        RECT 122.260 148.445 123.015 148.570 ;
        RECT 122.260 148.295 122.430 148.445 ;
        RECT 123.275 148.415 123.445 149.615 ;
        RECT 123.615 149.325 123.895 150.465 ;
        RECT 124.065 149.315 124.395 150.295 ;
        RECT 124.565 149.325 124.825 150.465 ;
        RECT 124.995 149.375 128.505 150.465 ;
        RECT 128.675 149.375 129.885 150.465 ;
        RECT 123.625 148.885 123.960 149.155 ;
        RECT 124.130 148.715 124.300 149.315 ;
        RECT 124.470 148.905 124.805 149.155 ;
        RECT 121.130 148.085 122.430 148.295 ;
        RECT 122.685 147.915 123.015 148.275 ;
        RECT 123.185 148.085 123.445 148.415 ;
        RECT 123.615 147.915 123.925 148.715 ;
        RECT 124.130 148.085 124.825 148.715 ;
        RECT 124.995 148.685 126.645 149.205 ;
        RECT 126.815 148.855 128.505 149.375 ;
        RECT 124.995 147.915 128.505 148.685 ;
        RECT 128.675 148.665 129.195 149.205 ;
        RECT 129.365 148.835 129.885 149.375 ;
        RECT 130.060 150.075 130.395 150.295 ;
        RECT 131.400 150.085 131.755 150.465 ;
        RECT 130.060 149.455 130.315 150.075 ;
        RECT 130.565 149.915 130.795 149.955 ;
        RECT 131.925 149.915 132.175 150.295 ;
        RECT 130.565 149.715 132.175 149.915 ;
        RECT 130.565 149.625 130.750 149.715 ;
        RECT 131.340 149.705 132.175 149.715 ;
        RECT 132.425 149.685 132.675 150.465 ;
        RECT 132.845 149.615 133.105 150.295 ;
        RECT 130.905 149.515 131.235 149.545 ;
        RECT 130.905 149.455 132.705 149.515 ;
        RECT 130.060 149.345 132.765 149.455 ;
        RECT 130.060 149.285 131.235 149.345 ;
        RECT 132.565 149.310 132.765 149.345 ;
        RECT 130.055 148.905 130.545 149.105 ;
        RECT 130.735 148.905 131.210 149.115 ;
        RECT 128.675 147.915 129.885 148.665 ;
        RECT 130.060 147.915 130.515 148.680 ;
        RECT 130.990 148.505 131.210 148.905 ;
        RECT 131.455 148.905 131.785 149.115 ;
        RECT 131.455 148.505 131.665 148.905 ;
        RECT 131.955 148.870 132.365 149.175 ;
        RECT 132.595 148.735 132.765 149.310 ;
        RECT 132.495 148.615 132.765 148.735 ;
        RECT 131.920 148.570 132.765 148.615 ;
        RECT 131.920 148.445 132.675 148.570 ;
        RECT 131.920 148.295 132.090 148.445 ;
        RECT 132.935 148.425 133.105 149.615 ;
        RECT 133.275 149.300 133.565 150.465 ;
        RECT 134.660 149.325 134.995 150.295 ;
        RECT 135.165 149.325 135.335 150.465 ;
        RECT 135.505 150.125 137.535 150.295 ;
        RECT 134.660 148.655 134.830 149.325 ;
        RECT 135.505 149.155 135.675 150.125 ;
        RECT 135.000 148.825 135.255 149.155 ;
        RECT 135.480 148.825 135.675 149.155 ;
        RECT 135.845 149.785 136.970 149.955 ;
        RECT 135.085 148.655 135.255 148.825 ;
        RECT 135.845 148.655 136.015 149.785 ;
        RECT 132.875 148.415 133.105 148.425 ;
        RECT 130.790 148.085 132.090 148.295 ;
        RECT 132.345 147.915 132.675 148.275 ;
        RECT 132.845 148.085 133.105 148.415 ;
        RECT 133.275 147.915 133.565 148.640 ;
        RECT 134.660 148.085 134.915 148.655 ;
        RECT 135.085 148.485 136.015 148.655 ;
        RECT 136.185 149.445 137.195 149.615 ;
        RECT 136.185 148.645 136.355 149.445 ;
        RECT 136.560 148.765 136.835 149.245 ;
        RECT 136.555 148.595 136.835 148.765 ;
        RECT 135.840 148.450 136.015 148.485 ;
        RECT 135.085 147.915 135.415 148.315 ;
        RECT 135.840 148.085 136.370 148.450 ;
        RECT 136.560 148.085 136.835 148.595 ;
        RECT 137.005 148.085 137.195 149.445 ;
        RECT 137.365 149.460 137.535 150.125 ;
        RECT 137.705 149.705 137.875 150.465 ;
        RECT 138.110 149.705 138.625 150.115 ;
        RECT 137.365 149.270 138.115 149.460 ;
        RECT 138.285 148.895 138.625 149.705 ;
        RECT 137.395 148.725 138.625 148.895 ;
        RECT 138.795 149.325 139.180 150.295 ;
        RECT 139.350 150.005 139.675 150.465 ;
        RECT 140.195 149.835 140.475 150.295 ;
        RECT 139.350 149.615 140.475 149.835 ;
        RECT 137.375 147.915 137.885 148.450 ;
        RECT 138.105 148.120 138.350 148.725 ;
        RECT 138.795 148.655 139.075 149.325 ;
        RECT 139.350 149.155 139.800 149.615 ;
        RECT 140.665 149.445 141.065 150.295 ;
        RECT 141.465 150.005 141.735 150.465 ;
        RECT 141.905 149.835 142.190 150.295 ;
        RECT 139.245 148.825 139.800 149.155 ;
        RECT 139.970 148.885 141.065 149.445 ;
        RECT 139.350 148.715 139.800 148.825 ;
        RECT 138.795 148.085 139.180 148.655 ;
        RECT 139.350 148.545 140.475 148.715 ;
        RECT 139.350 147.915 139.675 148.375 ;
        RECT 140.195 148.085 140.475 148.545 ;
        RECT 140.665 148.085 141.065 148.885 ;
        RECT 141.235 149.615 142.190 149.835 ;
        RECT 141.235 148.715 141.445 149.615 ;
        RECT 141.615 148.885 142.305 149.445 ;
        RECT 142.475 149.390 142.745 150.295 ;
        RECT 142.915 149.705 143.245 150.465 ;
        RECT 143.425 149.535 143.595 150.295 ;
        RECT 141.235 148.545 142.190 148.715 ;
        RECT 141.465 147.915 141.735 148.375 ;
        RECT 141.905 148.085 142.190 148.545 ;
        RECT 142.475 148.590 142.645 149.390 ;
        RECT 142.930 149.365 143.595 149.535 ;
        RECT 143.945 149.535 144.115 150.295 ;
        RECT 144.330 149.705 144.660 150.465 ;
        RECT 143.945 149.365 144.660 149.535 ;
        RECT 144.830 149.390 145.085 150.295 ;
        RECT 142.930 149.220 143.100 149.365 ;
        RECT 142.815 148.890 143.100 149.220 ;
        RECT 142.930 148.635 143.100 148.890 ;
        RECT 143.335 148.815 143.665 149.185 ;
        RECT 143.855 148.815 144.210 149.185 ;
        RECT 144.490 149.155 144.660 149.365 ;
        RECT 144.490 148.825 144.745 149.155 ;
        RECT 144.490 148.635 144.660 148.825 ;
        RECT 144.915 148.660 145.085 149.390 ;
        RECT 145.260 149.315 145.520 150.465 ;
        RECT 145.695 149.375 146.905 150.465 ;
        RECT 145.695 148.835 146.215 149.375 ;
        RECT 142.475 148.085 142.735 148.590 ;
        RECT 142.930 148.465 143.595 148.635 ;
        RECT 142.915 147.915 143.245 148.295 ;
        RECT 143.425 148.085 143.595 148.465 ;
        RECT 143.945 148.465 144.660 148.635 ;
        RECT 143.945 148.085 144.115 148.465 ;
        RECT 144.330 147.915 144.660 148.295 ;
        RECT 144.830 148.085 145.085 148.660 ;
        RECT 145.260 147.915 145.520 148.755 ;
        RECT 146.385 148.665 146.905 149.205 ;
        RECT 145.695 147.915 146.905 148.665 ;
        RECT 17.270 147.745 146.990 147.915 ;
        RECT 17.355 146.995 18.565 147.745 ;
        RECT 17.355 146.455 17.875 146.995 ;
        RECT 18.740 146.905 19.000 147.745 ;
        RECT 19.175 147.000 19.430 147.575 ;
        RECT 19.600 147.365 19.930 147.745 ;
        RECT 20.145 147.195 20.315 147.575 ;
        RECT 20.575 147.200 25.920 147.745 ;
        RECT 19.600 147.025 20.315 147.195 ;
        RECT 18.045 146.285 18.565 146.825 ;
        RECT 17.355 145.195 18.565 146.285 ;
        RECT 18.740 145.195 19.000 146.345 ;
        RECT 19.175 146.270 19.345 147.000 ;
        RECT 19.600 146.835 19.770 147.025 ;
        RECT 19.515 146.505 19.770 146.835 ;
        RECT 19.600 146.295 19.770 146.505 ;
        RECT 20.050 146.475 20.405 146.845 ;
        RECT 22.160 146.370 22.500 147.200 ;
        RECT 26.095 146.975 28.685 147.745 ;
        RECT 29.365 147.090 29.695 147.525 ;
        RECT 29.865 147.135 30.035 147.745 ;
        RECT 29.315 147.005 29.695 147.090 ;
        RECT 30.205 147.005 30.535 147.530 ;
        RECT 30.795 147.215 31.005 147.745 ;
        RECT 31.280 147.295 32.065 147.465 ;
        RECT 32.235 147.295 32.640 147.465 ;
        RECT 19.175 145.365 19.430 146.270 ;
        RECT 19.600 146.125 20.315 146.295 ;
        RECT 19.600 145.195 19.930 145.955 ;
        RECT 20.145 145.365 20.315 146.125 ;
        RECT 23.980 145.630 24.330 146.880 ;
        RECT 26.095 146.455 27.305 146.975 ;
        RECT 29.315 146.965 29.540 147.005 ;
        RECT 27.475 146.285 28.685 146.805 ;
        RECT 20.575 145.195 25.920 145.630 ;
        RECT 26.095 145.195 28.685 146.285 ;
        RECT 29.315 146.385 29.485 146.965 ;
        RECT 30.205 146.835 30.405 147.005 ;
        RECT 31.280 146.835 31.450 147.295 ;
        RECT 29.655 146.505 30.405 146.835 ;
        RECT 30.575 146.505 31.450 146.835 ;
        RECT 29.315 146.335 29.530 146.385 ;
        RECT 29.315 146.255 29.705 146.335 ;
        RECT 29.375 145.410 29.705 146.255 ;
        RECT 30.215 146.300 30.405 146.505 ;
        RECT 29.875 145.195 30.045 146.205 ;
        RECT 30.215 145.925 31.110 146.300 ;
        RECT 30.215 145.365 30.555 145.925 ;
        RECT 30.785 145.195 31.100 145.695 ;
        RECT 31.280 145.665 31.450 146.505 ;
        RECT 31.620 146.795 32.085 147.125 ;
        RECT 32.470 147.065 32.640 147.295 ;
        RECT 32.820 147.245 33.190 147.745 ;
        RECT 33.510 147.295 34.185 147.465 ;
        RECT 34.380 147.295 34.715 147.465 ;
        RECT 31.620 145.835 31.940 146.795 ;
        RECT 32.470 146.765 33.300 147.065 ;
        RECT 32.110 145.865 32.300 146.585 ;
        RECT 32.470 145.695 32.640 146.765 ;
        RECT 33.100 146.735 33.300 146.765 ;
        RECT 32.810 146.515 32.980 146.585 ;
        RECT 33.510 146.515 33.680 147.295 ;
        RECT 34.545 147.155 34.715 147.295 ;
        RECT 34.885 147.285 35.135 147.745 ;
        RECT 32.810 146.345 33.680 146.515 ;
        RECT 33.850 146.875 34.375 147.095 ;
        RECT 34.545 147.025 34.770 147.155 ;
        RECT 32.810 146.255 33.320 146.345 ;
        RECT 31.280 145.495 32.165 145.665 ;
        RECT 32.390 145.365 32.640 145.695 ;
        RECT 32.810 145.195 32.980 145.995 ;
        RECT 33.150 145.640 33.320 146.255 ;
        RECT 33.850 146.175 34.020 146.875 ;
        RECT 33.490 145.810 34.020 146.175 ;
        RECT 34.190 146.110 34.430 146.705 ;
        RECT 34.600 145.920 34.770 147.025 ;
        RECT 34.940 146.165 35.220 147.115 ;
        RECT 34.465 145.790 34.770 145.920 ;
        RECT 33.150 145.470 34.255 145.640 ;
        RECT 34.465 145.365 34.715 145.790 ;
        RECT 34.885 145.195 35.150 145.655 ;
        RECT 35.390 145.365 35.575 147.485 ;
        RECT 35.745 147.365 36.075 147.745 ;
        RECT 36.245 147.195 36.415 147.485 ;
        RECT 35.750 147.025 36.415 147.195 ;
        RECT 35.750 146.035 35.980 147.025 ;
        RECT 36.675 146.995 37.885 147.745 ;
        RECT 38.090 147.005 38.705 147.575 ;
        RECT 38.875 147.235 39.090 147.745 ;
        RECT 39.320 147.235 39.600 147.565 ;
        RECT 39.780 147.235 40.020 147.745 ;
        RECT 36.150 146.205 36.500 146.855 ;
        RECT 36.675 146.455 37.195 146.995 ;
        RECT 37.365 146.285 37.885 146.825 ;
        RECT 35.750 145.865 36.415 146.035 ;
        RECT 35.745 145.195 36.075 145.695 ;
        RECT 36.245 145.365 36.415 145.865 ;
        RECT 36.675 145.195 37.885 146.285 ;
        RECT 38.090 145.985 38.405 147.005 ;
        RECT 38.575 146.335 38.745 146.835 ;
        RECT 38.995 146.505 39.260 147.065 ;
        RECT 39.430 146.335 39.600 147.235 ;
        RECT 39.770 146.505 40.125 147.065 ;
        RECT 38.575 146.165 40.000 146.335 ;
        RECT 38.090 145.365 38.625 145.985 ;
        RECT 38.795 145.195 39.125 145.995 ;
        RECT 39.610 145.990 40.000 146.165 ;
        RECT 40.365 145.375 40.625 147.565 ;
        RECT 40.885 147.375 41.555 147.745 ;
        RECT 41.735 147.195 42.045 147.565 ;
        RECT 40.815 146.995 42.045 147.195 ;
        RECT 40.815 146.325 41.105 146.995 ;
        RECT 42.225 146.815 42.455 147.455 ;
        RECT 42.635 147.015 42.925 147.745 ;
        RECT 43.115 147.020 43.405 147.745 ;
        RECT 44.665 147.285 44.920 147.745 ;
        RECT 45.090 147.115 45.420 147.575 ;
        RECT 45.590 147.285 45.760 147.745 ;
        RECT 45.930 147.115 46.260 147.575 ;
        RECT 46.430 147.285 46.600 147.745 ;
        RECT 46.770 147.115 47.100 147.575 ;
        RECT 47.270 147.285 47.440 147.745 ;
        RECT 47.610 147.115 47.940 147.575 ;
        RECT 48.110 147.285 48.415 147.745 ;
        RECT 49.295 147.115 49.625 147.475 ;
        RECT 50.245 147.285 50.495 147.745 ;
        RECT 50.665 147.285 51.225 147.575 ;
        RECT 44.495 146.925 48.465 147.115 ;
        RECT 49.295 146.925 50.685 147.115 ;
        RECT 41.285 146.505 41.750 146.815 ;
        RECT 41.930 146.505 42.455 146.815 ;
        RECT 42.635 146.505 42.935 146.835 ;
        RECT 40.815 146.105 41.585 146.325 ;
        RECT 40.795 145.195 41.135 145.925 ;
        RECT 41.315 145.375 41.585 146.105 ;
        RECT 41.765 146.085 42.925 146.325 ;
        RECT 41.765 145.375 41.995 146.085 ;
        RECT 42.165 145.195 42.495 145.905 ;
        RECT 42.665 145.375 42.925 146.085 ;
        RECT 43.115 145.195 43.405 146.360 ;
        RECT 44.495 146.335 44.840 146.925 ;
        RECT 45.090 146.505 47.945 146.755 ;
        RECT 48.145 146.335 48.465 146.925 ;
        RECT 50.515 146.835 50.685 146.925 ;
        RECT 44.495 146.165 48.465 146.335 ;
        RECT 49.110 146.505 49.785 146.755 ;
        RECT 50.005 146.505 50.345 146.755 ;
        RECT 50.515 146.505 50.805 146.835 ;
        RECT 44.665 145.195 44.920 145.995 ;
        RECT 45.090 145.365 45.420 146.165 ;
        RECT 45.590 145.195 45.760 145.995 ;
        RECT 45.930 145.365 46.260 146.165 ;
        RECT 46.430 145.195 46.600 145.995 ;
        RECT 46.770 145.365 47.100 146.165 ;
        RECT 47.270 145.195 47.440 145.995 ;
        RECT 47.610 145.365 47.940 146.165 ;
        RECT 49.110 146.145 49.375 146.505 ;
        RECT 50.515 146.255 50.685 146.505 ;
        RECT 49.745 146.085 50.685 146.255 ;
        RECT 48.110 145.195 48.410 145.995 ;
        RECT 49.295 145.195 49.575 145.865 ;
        RECT 49.745 145.535 50.045 146.085 ;
        RECT 50.975 145.915 51.225 147.285 ;
        RECT 51.395 146.925 51.655 147.745 ;
        RECT 51.825 146.925 52.155 147.345 ;
        RECT 52.335 147.260 53.125 147.525 ;
        RECT 51.905 146.835 52.155 146.925 ;
        RECT 50.245 145.195 50.575 145.915 ;
        RECT 50.765 145.365 51.225 145.915 ;
        RECT 51.395 145.875 51.735 146.755 ;
        RECT 51.905 146.585 52.700 146.835 ;
        RECT 51.395 145.195 51.655 145.705 ;
        RECT 51.905 145.365 52.075 146.585 ;
        RECT 52.870 146.405 53.125 147.260 ;
        RECT 53.295 147.105 53.495 147.525 ;
        RECT 53.685 147.285 54.015 147.745 ;
        RECT 53.295 146.585 53.705 147.105 ;
        RECT 54.185 147.095 54.445 147.575 ;
        RECT 53.875 146.405 54.105 146.835 ;
        RECT 52.315 146.235 54.105 146.405 ;
        RECT 52.315 145.870 52.565 146.235 ;
        RECT 52.735 145.875 53.065 146.065 ;
        RECT 53.285 145.940 54.000 146.235 ;
        RECT 54.275 146.065 54.445 147.095 ;
        RECT 55.585 147.090 55.915 147.525 ;
        RECT 56.085 147.135 56.255 147.745 ;
        RECT 55.535 147.005 55.915 147.090 ;
        RECT 56.425 147.005 56.755 147.530 ;
        RECT 57.015 147.215 57.225 147.745 ;
        RECT 57.500 147.295 58.285 147.465 ;
        RECT 58.455 147.295 58.860 147.465 ;
        RECT 55.535 146.965 55.760 147.005 ;
        RECT 55.535 146.385 55.705 146.965 ;
        RECT 56.425 146.835 56.625 147.005 ;
        RECT 57.500 146.835 57.670 147.295 ;
        RECT 55.875 146.505 56.625 146.835 ;
        RECT 56.795 146.505 57.670 146.835 ;
        RECT 55.535 146.335 55.750 146.385 ;
        RECT 55.535 146.255 55.925 146.335 ;
        RECT 52.735 145.700 52.930 145.875 ;
        RECT 52.315 145.195 52.930 145.700 ;
        RECT 53.100 145.365 53.575 145.705 ;
        RECT 53.745 145.195 53.960 145.740 ;
        RECT 54.170 145.365 54.445 146.065 ;
        RECT 55.595 145.410 55.925 146.255 ;
        RECT 56.435 146.300 56.625 146.505 ;
        RECT 56.095 145.195 56.265 146.205 ;
        RECT 56.435 145.925 57.330 146.300 ;
        RECT 56.435 145.365 56.775 145.925 ;
        RECT 57.005 145.195 57.320 145.695 ;
        RECT 57.500 145.665 57.670 146.505 ;
        RECT 57.840 146.795 58.305 147.125 ;
        RECT 58.690 147.065 58.860 147.295 ;
        RECT 59.040 147.245 59.410 147.745 ;
        RECT 59.730 147.295 60.405 147.465 ;
        RECT 60.600 147.295 60.935 147.465 ;
        RECT 57.840 145.835 58.160 146.795 ;
        RECT 58.690 146.765 59.520 147.065 ;
        RECT 58.330 145.865 58.520 146.585 ;
        RECT 58.690 145.695 58.860 146.765 ;
        RECT 59.320 146.735 59.520 146.765 ;
        RECT 59.030 146.515 59.200 146.585 ;
        RECT 59.730 146.515 59.900 147.295 ;
        RECT 60.765 147.155 60.935 147.295 ;
        RECT 61.105 147.285 61.355 147.745 ;
        RECT 59.030 146.345 59.900 146.515 ;
        RECT 60.070 146.875 60.595 147.095 ;
        RECT 60.765 147.025 60.990 147.155 ;
        RECT 59.030 146.255 59.540 146.345 ;
        RECT 57.500 145.495 58.385 145.665 ;
        RECT 58.610 145.365 58.860 145.695 ;
        RECT 59.030 145.195 59.200 145.995 ;
        RECT 59.370 145.640 59.540 146.255 ;
        RECT 60.070 146.175 60.240 146.875 ;
        RECT 59.710 145.810 60.240 146.175 ;
        RECT 60.410 146.110 60.650 146.705 ;
        RECT 60.820 145.920 60.990 147.025 ;
        RECT 61.160 146.165 61.440 147.115 ;
        RECT 60.685 145.790 60.990 145.920 ;
        RECT 59.370 145.470 60.475 145.640 ;
        RECT 60.685 145.365 60.935 145.790 ;
        RECT 61.105 145.195 61.370 145.655 ;
        RECT 61.610 145.365 61.795 147.485 ;
        RECT 61.965 147.365 62.295 147.745 ;
        RECT 62.465 147.195 62.635 147.485 ;
        RECT 61.970 147.025 62.635 147.195 ;
        RECT 61.970 146.035 62.200 147.025 ;
        RECT 62.930 147.005 63.545 147.575 ;
        RECT 63.715 147.235 63.930 147.745 ;
        RECT 64.160 147.235 64.440 147.565 ;
        RECT 64.620 147.235 64.860 147.745 ;
        RECT 62.370 146.205 62.720 146.855 ;
        RECT 61.970 145.865 62.635 146.035 ;
        RECT 61.965 145.195 62.295 145.695 ;
        RECT 62.465 145.365 62.635 145.865 ;
        RECT 62.930 145.985 63.245 147.005 ;
        RECT 63.415 146.335 63.585 146.835 ;
        RECT 63.835 146.505 64.100 147.065 ;
        RECT 64.270 146.335 64.440 147.235 ;
        RECT 64.610 146.505 64.965 147.065 ;
        RECT 65.195 146.975 68.705 147.745 ;
        RECT 68.875 147.020 69.165 147.745 ;
        RECT 70.345 147.195 70.515 147.485 ;
        RECT 70.685 147.365 71.015 147.745 ;
        RECT 70.345 147.025 71.010 147.195 ;
        RECT 65.195 146.455 66.845 146.975 ;
        RECT 63.415 146.165 64.840 146.335 ;
        RECT 67.015 146.285 68.705 146.805 ;
        RECT 62.930 145.365 63.465 145.985 ;
        RECT 63.635 145.195 63.965 145.995 ;
        RECT 64.450 145.990 64.840 146.165 ;
        RECT 65.195 145.195 68.705 146.285 ;
        RECT 68.875 145.195 69.165 146.360 ;
        RECT 70.260 146.205 70.610 146.855 ;
        RECT 70.780 146.035 71.010 147.025 ;
        RECT 70.345 145.865 71.010 146.035 ;
        RECT 70.345 145.365 70.515 145.865 ;
        RECT 70.685 145.195 71.015 145.695 ;
        RECT 71.185 145.365 71.370 147.485 ;
        RECT 71.625 147.285 71.875 147.745 ;
        RECT 72.045 147.295 72.380 147.465 ;
        RECT 72.575 147.295 73.250 147.465 ;
        RECT 72.045 147.155 72.215 147.295 ;
        RECT 71.540 146.165 71.820 147.115 ;
        RECT 71.990 147.025 72.215 147.155 ;
        RECT 71.990 145.920 72.160 147.025 ;
        RECT 72.385 146.875 72.910 147.095 ;
        RECT 72.330 146.110 72.570 146.705 ;
        RECT 72.740 146.175 72.910 146.875 ;
        RECT 73.080 146.515 73.250 147.295 ;
        RECT 73.570 147.245 73.940 147.745 ;
        RECT 74.120 147.295 74.525 147.465 ;
        RECT 74.695 147.295 75.480 147.465 ;
        RECT 74.120 147.065 74.290 147.295 ;
        RECT 73.460 146.765 74.290 147.065 ;
        RECT 74.675 146.795 75.140 147.125 ;
        RECT 73.460 146.735 73.660 146.765 ;
        RECT 73.780 146.515 73.950 146.585 ;
        RECT 73.080 146.345 73.950 146.515 ;
        RECT 73.440 146.255 73.950 146.345 ;
        RECT 71.990 145.790 72.295 145.920 ;
        RECT 72.740 145.810 73.270 146.175 ;
        RECT 71.610 145.195 71.875 145.655 ;
        RECT 72.045 145.365 72.295 145.790 ;
        RECT 73.440 145.640 73.610 146.255 ;
        RECT 72.505 145.470 73.610 145.640 ;
        RECT 73.780 145.195 73.950 145.995 ;
        RECT 74.120 145.695 74.290 146.765 ;
        RECT 74.460 145.865 74.650 146.585 ;
        RECT 74.820 145.835 75.140 146.795 ;
        RECT 75.310 146.835 75.480 147.295 ;
        RECT 75.755 147.215 75.965 147.745 ;
        RECT 76.225 147.005 76.555 147.530 ;
        RECT 76.725 147.135 76.895 147.745 ;
        RECT 77.065 147.090 77.395 147.525 ;
        RECT 78.650 147.115 78.935 147.575 ;
        RECT 79.105 147.285 79.375 147.745 ;
        RECT 77.065 147.005 77.445 147.090 ;
        RECT 76.355 146.835 76.555 147.005 ;
        RECT 77.220 146.965 77.445 147.005 ;
        RECT 75.310 146.505 76.185 146.835 ;
        RECT 76.355 146.505 77.105 146.835 ;
        RECT 74.120 145.365 74.370 145.695 ;
        RECT 75.310 145.665 75.480 146.505 ;
        RECT 76.355 146.300 76.545 146.505 ;
        RECT 77.275 146.385 77.445 146.965 ;
        RECT 78.650 146.945 79.605 147.115 ;
        RECT 77.230 146.335 77.445 146.385 ;
        RECT 75.650 145.925 76.545 146.300 ;
        RECT 77.055 146.255 77.445 146.335 ;
        RECT 74.595 145.495 75.480 145.665 ;
        RECT 75.660 145.195 75.975 145.695 ;
        RECT 76.205 145.365 76.545 145.925 ;
        RECT 76.715 145.195 76.885 146.205 ;
        RECT 77.055 145.410 77.385 146.255 ;
        RECT 78.535 146.215 79.225 146.775 ;
        RECT 79.395 146.045 79.605 146.945 ;
        RECT 78.650 145.825 79.605 146.045 ;
        RECT 79.775 146.775 80.175 147.575 ;
        RECT 80.365 147.115 80.645 147.575 ;
        RECT 81.165 147.285 81.490 147.745 ;
        RECT 80.365 146.945 81.490 147.115 ;
        RECT 81.660 147.005 82.045 147.575 ;
        RECT 81.040 146.835 81.490 146.945 ;
        RECT 79.775 146.215 80.870 146.775 ;
        RECT 81.040 146.505 81.595 146.835 ;
        RECT 78.650 145.365 78.935 145.825 ;
        RECT 79.105 145.195 79.375 145.655 ;
        RECT 79.775 145.365 80.175 146.215 ;
        RECT 81.040 146.045 81.490 146.505 ;
        RECT 81.765 146.335 82.045 147.005 ;
        RECT 82.330 147.115 82.615 147.575 ;
        RECT 82.785 147.285 83.055 147.745 ;
        RECT 82.330 146.945 83.285 147.115 ;
        RECT 80.365 145.825 81.490 146.045 ;
        RECT 80.365 145.365 80.645 145.825 ;
        RECT 81.165 145.195 81.490 145.655 ;
        RECT 81.660 145.365 82.045 146.335 ;
        RECT 82.215 146.215 82.905 146.775 ;
        RECT 83.075 146.045 83.285 146.945 ;
        RECT 82.330 145.825 83.285 146.045 ;
        RECT 83.455 146.775 83.855 147.575 ;
        RECT 84.045 147.115 84.325 147.575 ;
        RECT 84.845 147.285 85.170 147.745 ;
        RECT 84.045 146.945 85.170 147.115 ;
        RECT 85.340 147.005 85.725 147.575 ;
        RECT 85.915 147.175 86.170 147.525 ;
        RECT 86.340 147.345 86.670 147.745 ;
        RECT 86.840 147.175 87.010 147.525 ;
        RECT 87.180 147.345 87.560 147.745 ;
        RECT 85.915 147.005 87.580 147.175 ;
        RECT 87.750 147.070 88.025 147.415 ;
        RECT 84.720 146.835 85.170 146.945 ;
        RECT 83.455 146.215 84.550 146.775 ;
        RECT 84.720 146.505 85.275 146.835 ;
        RECT 82.330 145.365 82.615 145.825 ;
        RECT 82.785 145.195 83.055 145.655 ;
        RECT 83.455 145.365 83.855 146.215 ;
        RECT 84.720 146.045 85.170 146.505 ;
        RECT 85.445 146.335 85.725 147.005 ;
        RECT 87.410 146.835 87.580 147.005 ;
        RECT 85.895 146.505 86.245 146.835 ;
        RECT 86.415 146.505 87.240 146.835 ;
        RECT 87.410 146.505 87.685 146.835 ;
        RECT 84.045 145.825 85.170 146.045 ;
        RECT 84.045 145.365 84.325 145.825 ;
        RECT 84.845 145.195 85.170 145.655 ;
        RECT 85.340 145.365 85.725 146.335 ;
        RECT 85.915 146.045 86.245 146.335 ;
        RECT 86.415 146.215 86.640 146.505 ;
        RECT 87.410 146.335 87.580 146.505 ;
        RECT 87.855 146.335 88.025 147.070 ;
        RECT 88.195 146.915 88.485 147.745 ;
        RECT 88.655 147.200 94.000 147.745 ;
        RECT 86.910 146.165 87.580 146.335 ;
        RECT 86.910 146.045 87.080 146.165 ;
        RECT 85.915 145.875 87.080 146.045 ;
        RECT 85.895 145.415 87.090 145.705 ;
        RECT 87.260 145.195 87.540 145.995 ;
        RECT 87.750 145.365 88.025 146.335 ;
        RECT 88.195 145.195 88.485 146.400 ;
        RECT 90.240 146.370 90.580 147.200 ;
        RECT 94.635 147.020 94.925 147.745 ;
        RECT 95.095 146.975 97.685 147.745 ;
        RECT 97.905 147.205 98.130 147.565 ;
        RECT 98.310 147.375 98.640 147.745 ;
        RECT 98.820 147.205 99.075 147.565 ;
        RECT 99.640 147.375 100.385 147.745 ;
        RECT 97.905 147.015 100.390 147.205 ;
        RECT 92.060 145.630 92.410 146.880 ;
        RECT 95.095 146.455 96.305 146.975 ;
        RECT 88.655 145.195 94.000 145.630 ;
        RECT 94.635 145.195 94.925 146.360 ;
        RECT 96.475 146.285 97.685 146.805 ;
        RECT 97.865 146.505 98.135 146.835 ;
        RECT 98.315 146.505 98.750 146.835 ;
        RECT 98.930 146.505 99.505 146.835 ;
        RECT 99.685 146.505 99.965 146.835 ;
        RECT 100.165 146.325 100.390 147.015 ;
        RECT 95.095 145.195 97.685 146.285 ;
        RECT 97.895 146.145 100.390 146.325 ;
        RECT 100.565 146.145 100.900 147.565 ;
        RECT 102.085 147.195 102.255 147.485 ;
        RECT 102.425 147.365 102.755 147.745 ;
        RECT 102.085 147.025 102.750 147.195 ;
        RECT 102.000 146.205 102.350 146.855 ;
        RECT 97.895 145.375 98.185 146.145 ;
        RECT 98.755 145.735 99.945 145.965 ;
        RECT 98.755 145.375 99.015 145.735 ;
        RECT 99.185 145.195 99.515 145.565 ;
        RECT 99.685 145.375 99.945 145.735 ;
        RECT 100.135 145.195 100.465 145.915 ;
        RECT 100.635 145.375 100.900 146.145 ;
        RECT 102.520 146.035 102.750 147.025 ;
        RECT 102.085 145.865 102.750 146.035 ;
        RECT 102.085 145.365 102.255 145.865 ;
        RECT 102.425 145.195 102.755 145.695 ;
        RECT 102.925 145.365 103.110 147.485 ;
        RECT 103.365 147.285 103.615 147.745 ;
        RECT 103.785 147.295 104.120 147.465 ;
        RECT 104.315 147.295 104.990 147.465 ;
        RECT 103.785 147.155 103.955 147.295 ;
        RECT 103.280 146.165 103.560 147.115 ;
        RECT 103.730 147.025 103.955 147.155 ;
        RECT 103.730 145.920 103.900 147.025 ;
        RECT 104.125 146.875 104.650 147.095 ;
        RECT 104.070 146.110 104.310 146.705 ;
        RECT 104.480 146.175 104.650 146.875 ;
        RECT 104.820 146.515 104.990 147.295 ;
        RECT 105.310 147.245 105.680 147.745 ;
        RECT 105.860 147.295 106.265 147.465 ;
        RECT 106.435 147.295 107.220 147.465 ;
        RECT 105.860 147.065 106.030 147.295 ;
        RECT 105.200 146.765 106.030 147.065 ;
        RECT 106.415 146.795 106.880 147.125 ;
        RECT 105.200 146.735 105.400 146.765 ;
        RECT 105.520 146.515 105.690 146.585 ;
        RECT 104.820 146.345 105.690 146.515 ;
        RECT 105.180 146.255 105.690 146.345 ;
        RECT 103.730 145.790 104.035 145.920 ;
        RECT 104.480 145.810 105.010 146.175 ;
        RECT 103.350 145.195 103.615 145.655 ;
        RECT 103.785 145.365 104.035 145.790 ;
        RECT 105.180 145.640 105.350 146.255 ;
        RECT 104.245 145.470 105.350 145.640 ;
        RECT 105.520 145.195 105.690 145.995 ;
        RECT 105.860 145.695 106.030 146.765 ;
        RECT 106.200 145.865 106.390 146.585 ;
        RECT 106.560 145.835 106.880 146.795 ;
        RECT 107.050 146.835 107.220 147.295 ;
        RECT 107.495 147.215 107.705 147.745 ;
        RECT 107.965 147.005 108.295 147.530 ;
        RECT 108.465 147.135 108.635 147.745 ;
        RECT 108.805 147.090 109.135 147.525 ;
        RECT 109.445 147.195 109.615 147.485 ;
        RECT 109.785 147.365 110.115 147.745 ;
        RECT 108.805 147.005 109.185 147.090 ;
        RECT 109.445 147.025 110.110 147.195 ;
        RECT 108.095 146.835 108.295 147.005 ;
        RECT 108.960 146.965 109.185 147.005 ;
        RECT 107.050 146.505 107.925 146.835 ;
        RECT 108.095 146.505 108.845 146.835 ;
        RECT 105.860 145.365 106.110 145.695 ;
        RECT 107.050 145.665 107.220 146.505 ;
        RECT 108.095 146.300 108.285 146.505 ;
        RECT 109.015 146.385 109.185 146.965 ;
        RECT 108.970 146.335 109.185 146.385 ;
        RECT 107.390 145.925 108.285 146.300 ;
        RECT 108.795 146.255 109.185 146.335 ;
        RECT 106.335 145.495 107.220 145.665 ;
        RECT 107.400 145.195 107.715 145.695 ;
        RECT 107.945 145.365 108.285 145.925 ;
        RECT 108.455 145.195 108.625 146.205 ;
        RECT 108.795 145.410 109.125 146.255 ;
        RECT 109.360 146.205 109.710 146.855 ;
        RECT 109.880 146.035 110.110 147.025 ;
        RECT 109.445 145.865 110.110 146.035 ;
        RECT 109.445 145.365 109.615 145.865 ;
        RECT 109.785 145.195 110.115 145.695 ;
        RECT 110.285 145.365 110.470 147.485 ;
        RECT 110.725 147.285 110.975 147.745 ;
        RECT 111.145 147.295 111.480 147.465 ;
        RECT 111.675 147.295 112.350 147.465 ;
        RECT 111.145 147.155 111.315 147.295 ;
        RECT 110.640 146.165 110.920 147.115 ;
        RECT 111.090 147.025 111.315 147.155 ;
        RECT 111.090 145.920 111.260 147.025 ;
        RECT 111.485 146.875 112.010 147.095 ;
        RECT 111.430 146.110 111.670 146.705 ;
        RECT 111.840 146.175 112.010 146.875 ;
        RECT 112.180 146.515 112.350 147.295 ;
        RECT 112.670 147.245 113.040 147.745 ;
        RECT 113.220 147.295 113.625 147.465 ;
        RECT 113.795 147.295 114.580 147.465 ;
        RECT 113.220 147.065 113.390 147.295 ;
        RECT 112.560 146.765 113.390 147.065 ;
        RECT 113.775 146.795 114.240 147.125 ;
        RECT 112.560 146.735 112.760 146.765 ;
        RECT 112.880 146.515 113.050 146.585 ;
        RECT 112.180 146.345 113.050 146.515 ;
        RECT 112.540 146.255 113.050 146.345 ;
        RECT 111.090 145.790 111.395 145.920 ;
        RECT 111.840 145.810 112.370 146.175 ;
        RECT 110.710 145.195 110.975 145.655 ;
        RECT 111.145 145.365 111.395 145.790 ;
        RECT 112.540 145.640 112.710 146.255 ;
        RECT 111.605 145.470 112.710 145.640 ;
        RECT 112.880 145.195 113.050 145.995 ;
        RECT 113.220 145.695 113.390 146.765 ;
        RECT 113.560 145.865 113.750 146.585 ;
        RECT 113.920 145.835 114.240 146.795 ;
        RECT 114.410 146.835 114.580 147.295 ;
        RECT 114.855 147.215 115.065 147.745 ;
        RECT 115.325 147.005 115.655 147.530 ;
        RECT 115.825 147.135 115.995 147.745 ;
        RECT 116.165 147.090 116.495 147.525 ;
        RECT 116.165 147.005 116.545 147.090 ;
        RECT 115.455 146.835 115.655 147.005 ;
        RECT 116.320 146.965 116.545 147.005 ;
        RECT 114.410 146.505 115.285 146.835 ;
        RECT 115.455 146.505 116.205 146.835 ;
        RECT 113.220 145.365 113.470 145.695 ;
        RECT 114.410 145.665 114.580 146.505 ;
        RECT 115.455 146.300 115.645 146.505 ;
        RECT 116.375 146.385 116.545 146.965 ;
        RECT 116.715 146.975 120.225 147.745 ;
        RECT 120.395 147.020 120.685 147.745 ;
        RECT 120.855 147.005 121.240 147.575 ;
        RECT 121.410 147.285 121.735 147.745 ;
        RECT 122.255 147.115 122.535 147.575 ;
        RECT 116.715 146.455 118.365 146.975 ;
        RECT 116.330 146.335 116.545 146.385 ;
        RECT 114.750 145.925 115.645 146.300 ;
        RECT 116.155 146.255 116.545 146.335 ;
        RECT 118.535 146.285 120.225 146.805 ;
        RECT 113.695 145.495 114.580 145.665 ;
        RECT 114.760 145.195 115.075 145.695 ;
        RECT 115.305 145.365 115.645 145.925 ;
        RECT 115.815 145.195 115.985 146.205 ;
        RECT 116.155 145.410 116.485 146.255 ;
        RECT 116.715 145.195 120.225 146.285 ;
        RECT 120.395 145.195 120.685 146.360 ;
        RECT 120.855 146.335 121.135 147.005 ;
        RECT 121.410 146.945 122.535 147.115 ;
        RECT 121.410 146.835 121.860 146.945 ;
        RECT 121.305 146.505 121.860 146.835 ;
        RECT 122.725 146.775 123.125 147.575 ;
        RECT 123.525 147.285 123.795 147.745 ;
        RECT 123.965 147.115 124.250 147.575 ;
        RECT 120.855 145.365 121.240 146.335 ;
        RECT 121.410 146.045 121.860 146.505 ;
        RECT 122.030 146.215 123.125 146.775 ;
        RECT 121.410 145.825 122.535 146.045 ;
        RECT 121.410 145.195 121.735 145.655 ;
        RECT 122.255 145.365 122.535 145.825 ;
        RECT 122.725 145.365 123.125 146.215 ;
        RECT 123.295 146.945 124.250 147.115 ;
        RECT 124.535 146.975 128.045 147.745 ;
        RECT 128.215 146.995 129.425 147.745 ;
        RECT 123.295 146.045 123.505 146.945 ;
        RECT 123.675 146.215 124.365 146.775 ;
        RECT 124.535 146.455 126.185 146.975 ;
        RECT 126.355 146.285 128.045 146.805 ;
        RECT 128.215 146.455 128.735 146.995 ;
        RECT 129.600 146.980 130.055 147.745 ;
        RECT 130.330 147.365 131.630 147.575 ;
        RECT 131.885 147.385 132.215 147.745 ;
        RECT 131.460 147.215 131.630 147.365 ;
        RECT 132.385 147.245 132.645 147.575 ;
        RECT 128.905 146.285 129.425 146.825 ;
        RECT 130.530 146.755 130.750 147.155 ;
        RECT 129.595 146.555 130.085 146.755 ;
        RECT 130.275 146.545 130.750 146.755 ;
        RECT 130.995 146.755 131.205 147.155 ;
        RECT 131.460 147.090 132.215 147.215 ;
        RECT 131.460 147.045 132.305 147.090 ;
        RECT 132.035 146.925 132.305 147.045 ;
        RECT 130.995 146.545 131.325 146.755 ;
        RECT 131.495 146.485 131.905 146.790 ;
        RECT 123.295 145.825 124.250 146.045 ;
        RECT 123.525 145.195 123.795 145.655 ;
        RECT 123.965 145.365 124.250 145.825 ;
        RECT 124.535 145.195 128.045 146.285 ;
        RECT 128.215 145.195 129.425 146.285 ;
        RECT 129.600 146.315 130.775 146.375 ;
        RECT 132.135 146.350 132.305 146.925 ;
        RECT 132.105 146.315 132.305 146.350 ;
        RECT 129.600 146.205 132.305 146.315 ;
        RECT 129.600 145.585 129.855 146.205 ;
        RECT 130.445 146.145 132.245 146.205 ;
        RECT 130.445 146.115 130.775 146.145 ;
        RECT 132.475 146.045 132.645 147.245 ;
        RECT 133.365 147.195 133.535 147.485 ;
        RECT 133.705 147.365 134.035 147.745 ;
        RECT 133.365 147.025 134.030 147.195 ;
        RECT 133.280 146.205 133.630 146.855 ;
        RECT 130.105 145.945 130.290 146.035 ;
        RECT 130.880 145.945 131.715 145.955 ;
        RECT 130.105 145.745 131.715 145.945 ;
        RECT 130.105 145.705 130.335 145.745 ;
        RECT 129.600 145.365 129.935 145.585 ;
        RECT 130.940 145.195 131.295 145.575 ;
        RECT 131.465 145.365 131.715 145.745 ;
        RECT 131.965 145.195 132.215 145.975 ;
        RECT 132.385 145.365 132.645 146.045 ;
        RECT 133.800 146.035 134.030 147.025 ;
        RECT 133.365 145.865 134.030 146.035 ;
        RECT 133.365 145.365 133.535 145.865 ;
        RECT 133.705 145.195 134.035 145.695 ;
        RECT 134.205 145.365 134.390 147.485 ;
        RECT 134.645 147.285 134.895 147.745 ;
        RECT 135.065 147.295 135.400 147.465 ;
        RECT 135.595 147.295 136.270 147.465 ;
        RECT 135.065 147.155 135.235 147.295 ;
        RECT 134.560 146.165 134.840 147.115 ;
        RECT 135.010 147.025 135.235 147.155 ;
        RECT 135.010 145.920 135.180 147.025 ;
        RECT 135.405 146.875 135.930 147.095 ;
        RECT 135.350 146.110 135.590 146.705 ;
        RECT 135.760 146.175 135.930 146.875 ;
        RECT 136.100 146.515 136.270 147.295 ;
        RECT 136.590 147.245 136.960 147.745 ;
        RECT 137.140 147.295 137.545 147.465 ;
        RECT 137.715 147.295 138.500 147.465 ;
        RECT 137.140 147.065 137.310 147.295 ;
        RECT 136.480 146.765 137.310 147.065 ;
        RECT 137.695 146.795 138.160 147.125 ;
        RECT 136.480 146.735 136.680 146.765 ;
        RECT 136.800 146.515 136.970 146.585 ;
        RECT 136.100 146.345 136.970 146.515 ;
        RECT 136.460 146.255 136.970 146.345 ;
        RECT 135.010 145.790 135.315 145.920 ;
        RECT 135.760 145.810 136.290 146.175 ;
        RECT 134.630 145.195 134.895 145.655 ;
        RECT 135.065 145.365 135.315 145.790 ;
        RECT 136.460 145.640 136.630 146.255 ;
        RECT 135.525 145.470 136.630 145.640 ;
        RECT 136.800 145.195 136.970 145.995 ;
        RECT 137.140 145.695 137.310 146.765 ;
        RECT 137.480 145.865 137.670 146.585 ;
        RECT 137.840 145.835 138.160 146.795 ;
        RECT 138.330 146.835 138.500 147.295 ;
        RECT 138.775 147.215 138.985 147.745 ;
        RECT 139.245 147.005 139.575 147.530 ;
        RECT 139.745 147.135 139.915 147.745 ;
        RECT 140.085 147.090 140.415 147.525 ;
        RECT 140.725 147.195 140.895 147.575 ;
        RECT 141.075 147.365 141.405 147.745 ;
        RECT 140.085 147.005 140.465 147.090 ;
        RECT 140.725 147.025 141.390 147.195 ;
        RECT 141.585 147.070 141.845 147.575 ;
        RECT 139.375 146.835 139.575 147.005 ;
        RECT 140.240 146.965 140.465 147.005 ;
        RECT 138.330 146.505 139.205 146.835 ;
        RECT 139.375 146.505 140.125 146.835 ;
        RECT 137.140 145.365 137.390 145.695 ;
        RECT 138.330 145.665 138.500 146.505 ;
        RECT 139.375 146.300 139.565 146.505 ;
        RECT 140.295 146.385 140.465 146.965 ;
        RECT 140.655 146.475 140.985 146.845 ;
        RECT 141.220 146.770 141.390 147.025 ;
        RECT 140.250 146.335 140.465 146.385 ;
        RECT 138.670 145.925 139.565 146.300 ;
        RECT 140.075 146.255 140.465 146.335 ;
        RECT 141.220 146.440 141.505 146.770 ;
        RECT 141.220 146.295 141.390 146.440 ;
        RECT 137.615 145.495 138.500 145.665 ;
        RECT 138.680 145.195 138.995 145.695 ;
        RECT 139.225 145.365 139.565 145.925 ;
        RECT 139.735 145.195 139.905 146.205 ;
        RECT 140.075 145.410 140.405 146.255 ;
        RECT 140.725 146.125 141.390 146.295 ;
        RECT 141.675 146.270 141.845 147.070 ;
        RECT 142.105 147.195 142.275 147.575 ;
        RECT 142.490 147.365 142.820 147.745 ;
        RECT 142.105 147.025 142.820 147.195 ;
        RECT 142.015 146.475 142.370 146.845 ;
        RECT 142.650 146.835 142.820 147.025 ;
        RECT 142.990 147.000 143.245 147.575 ;
        RECT 142.650 146.505 142.905 146.835 ;
        RECT 142.650 146.295 142.820 146.505 ;
        RECT 140.725 145.365 140.895 146.125 ;
        RECT 141.075 145.195 141.405 145.955 ;
        RECT 141.575 145.365 141.845 146.270 ;
        RECT 142.105 146.125 142.820 146.295 ;
        RECT 143.075 146.270 143.245 147.000 ;
        RECT 143.420 146.905 143.680 147.745 ;
        RECT 143.945 147.195 144.115 147.575 ;
        RECT 144.330 147.365 144.660 147.745 ;
        RECT 143.945 147.025 144.660 147.195 ;
        RECT 143.855 146.475 144.210 146.845 ;
        RECT 144.490 146.835 144.660 147.025 ;
        RECT 144.830 147.000 145.085 147.575 ;
        RECT 144.490 146.505 144.745 146.835 ;
        RECT 142.105 145.365 142.275 146.125 ;
        RECT 142.490 145.195 142.820 145.955 ;
        RECT 142.990 145.365 143.245 146.270 ;
        RECT 143.420 145.195 143.680 146.345 ;
        RECT 144.490 146.295 144.660 146.505 ;
        RECT 143.945 146.125 144.660 146.295 ;
        RECT 144.915 146.270 145.085 147.000 ;
        RECT 145.260 146.905 145.520 147.745 ;
        RECT 145.695 146.995 146.905 147.745 ;
        RECT 143.945 145.365 144.115 146.125 ;
        RECT 144.330 145.195 144.660 145.955 ;
        RECT 144.830 145.365 145.085 146.270 ;
        RECT 145.260 145.195 145.520 146.345 ;
        RECT 145.695 146.285 146.215 146.825 ;
        RECT 146.385 146.455 146.905 146.995 ;
        RECT 145.695 145.195 146.905 146.285 ;
        RECT 17.270 145.025 146.990 145.195 ;
        RECT 17.355 143.935 18.565 145.025 ;
        RECT 17.355 143.225 17.875 143.765 ;
        RECT 18.045 143.395 18.565 143.935 ;
        RECT 18.740 143.875 19.000 145.025 ;
        RECT 19.175 143.950 19.430 144.855 ;
        RECT 19.600 144.265 19.930 145.025 ;
        RECT 20.145 144.095 20.315 144.855 ;
        RECT 20.575 144.590 25.920 145.025 ;
        RECT 17.355 142.475 18.565 143.225 ;
        RECT 18.740 142.475 19.000 143.315 ;
        RECT 19.175 143.220 19.345 143.950 ;
        RECT 19.600 143.925 20.315 144.095 ;
        RECT 19.600 143.715 19.770 143.925 ;
        RECT 19.515 143.385 19.770 143.715 ;
        RECT 19.175 142.645 19.430 143.220 ;
        RECT 19.600 143.195 19.770 143.385 ;
        RECT 20.050 143.375 20.405 143.745 ;
        RECT 19.600 143.025 20.315 143.195 ;
        RECT 19.600 142.475 19.930 142.855 ;
        RECT 20.145 142.645 20.315 143.025 ;
        RECT 22.160 143.020 22.500 143.850 ;
        RECT 23.980 143.340 24.330 144.590 ;
        RECT 26.095 143.935 29.605 145.025 ;
        RECT 26.095 143.245 27.745 143.765 ;
        RECT 27.915 143.415 29.605 143.935 ;
        RECT 30.235 143.860 30.525 145.025 ;
        RECT 30.695 143.935 34.205 145.025 ;
        RECT 35.295 144.470 35.900 145.025 ;
        RECT 36.075 144.515 36.555 144.855 ;
        RECT 36.725 144.480 36.980 145.025 ;
        RECT 35.295 144.370 35.910 144.470 ;
        RECT 35.725 144.345 35.910 144.370 ;
        RECT 30.695 143.245 32.345 143.765 ;
        RECT 32.515 143.415 34.205 143.935 ;
        RECT 35.295 143.750 35.555 144.200 ;
        RECT 35.725 144.100 36.055 144.345 ;
        RECT 36.225 144.025 36.980 144.275 ;
        RECT 37.150 144.155 37.425 144.855 ;
        RECT 37.595 144.515 37.855 145.025 ;
        RECT 36.210 143.990 36.980 144.025 ;
        RECT 36.195 143.980 36.980 143.990 ;
        RECT 36.190 143.965 37.085 143.980 ;
        RECT 36.170 143.950 37.085 143.965 ;
        RECT 36.150 143.940 37.085 143.950 ;
        RECT 36.125 143.930 37.085 143.940 ;
        RECT 36.055 143.900 37.085 143.930 ;
        RECT 36.035 143.870 37.085 143.900 ;
        RECT 36.015 143.840 37.085 143.870 ;
        RECT 35.985 143.815 37.085 143.840 ;
        RECT 35.950 143.780 37.085 143.815 ;
        RECT 35.920 143.775 37.085 143.780 ;
        RECT 35.920 143.770 36.310 143.775 ;
        RECT 35.920 143.760 36.285 143.770 ;
        RECT 35.920 143.755 36.270 143.760 ;
        RECT 35.920 143.750 36.255 143.755 ;
        RECT 35.295 143.745 36.255 143.750 ;
        RECT 35.295 143.735 36.245 143.745 ;
        RECT 35.295 143.730 36.235 143.735 ;
        RECT 35.295 143.720 36.225 143.730 ;
        RECT 35.295 143.710 36.220 143.720 ;
        RECT 35.295 143.705 36.215 143.710 ;
        RECT 35.295 143.690 36.205 143.705 ;
        RECT 35.295 143.675 36.200 143.690 ;
        RECT 35.295 143.650 36.190 143.675 ;
        RECT 35.295 143.580 36.185 143.650 ;
        RECT 20.575 142.475 25.920 143.020 ;
        RECT 26.095 142.475 29.605 143.245 ;
        RECT 30.235 142.475 30.525 143.200 ;
        RECT 30.695 142.475 34.205 143.245 ;
        RECT 35.295 143.025 35.845 143.410 ;
        RECT 36.015 142.855 36.185 143.580 ;
        RECT 35.295 142.685 36.185 142.855 ;
        RECT 36.355 143.180 36.685 143.605 ;
        RECT 36.855 143.380 37.085 143.775 ;
        RECT 36.355 142.695 36.575 143.180 ;
        RECT 37.255 143.125 37.425 144.155 ;
        RECT 37.595 143.465 37.935 144.345 ;
        RECT 38.105 143.635 38.275 144.855 ;
        RECT 38.515 144.520 39.130 145.025 ;
        RECT 38.515 143.985 38.765 144.350 ;
        RECT 38.935 144.345 39.130 144.520 ;
        RECT 39.300 144.515 39.775 144.855 ;
        RECT 39.945 144.480 40.160 145.025 ;
        RECT 38.935 144.155 39.265 144.345 ;
        RECT 39.485 143.985 40.200 144.280 ;
        RECT 40.370 144.155 40.645 144.855 ;
        RECT 40.905 144.355 41.075 144.855 ;
        RECT 41.245 144.525 41.575 145.025 ;
        RECT 40.905 144.185 41.570 144.355 ;
        RECT 38.515 143.815 40.305 143.985 ;
        RECT 38.105 143.385 38.900 143.635 ;
        RECT 38.105 143.295 38.355 143.385 ;
        RECT 36.745 142.475 36.995 143.015 ;
        RECT 37.165 142.645 37.425 143.125 ;
        RECT 37.595 142.475 37.855 143.295 ;
        RECT 38.025 142.875 38.355 143.295 ;
        RECT 39.070 142.960 39.325 143.815 ;
        RECT 38.535 142.695 39.325 142.960 ;
        RECT 39.495 143.115 39.905 143.635 ;
        RECT 40.075 143.385 40.305 143.815 ;
        RECT 40.475 143.125 40.645 144.155 ;
        RECT 40.820 143.365 41.170 144.015 ;
        RECT 41.340 143.195 41.570 144.185 ;
        RECT 39.495 142.695 39.695 143.115 ;
        RECT 39.885 142.475 40.215 142.935 ;
        RECT 40.385 142.645 40.645 143.125 ;
        RECT 40.905 143.025 41.570 143.195 ;
        RECT 40.905 142.735 41.075 143.025 ;
        RECT 41.245 142.475 41.575 142.855 ;
        RECT 41.745 142.735 41.930 144.855 ;
        RECT 42.170 144.565 42.435 145.025 ;
        RECT 42.605 144.430 42.855 144.855 ;
        RECT 43.065 144.580 44.170 144.750 ;
        RECT 42.550 144.300 42.855 144.430 ;
        RECT 42.100 143.105 42.380 144.055 ;
        RECT 42.550 143.195 42.720 144.300 ;
        RECT 42.890 143.515 43.130 144.110 ;
        RECT 43.300 144.045 43.830 144.410 ;
        RECT 43.300 143.345 43.470 144.045 ;
        RECT 44.000 143.965 44.170 144.580 ;
        RECT 44.340 144.225 44.510 145.025 ;
        RECT 44.680 144.525 44.930 144.855 ;
        RECT 45.155 144.555 46.040 144.725 ;
        RECT 44.000 143.875 44.510 143.965 ;
        RECT 42.550 143.065 42.775 143.195 ;
        RECT 42.945 143.125 43.470 143.345 ;
        RECT 43.640 143.705 44.510 143.875 ;
        RECT 42.185 142.475 42.435 142.935 ;
        RECT 42.605 142.925 42.775 143.065 ;
        RECT 43.640 142.925 43.810 143.705 ;
        RECT 44.340 143.635 44.510 143.705 ;
        RECT 44.020 143.455 44.220 143.485 ;
        RECT 44.680 143.455 44.850 144.525 ;
        RECT 45.020 143.635 45.210 144.355 ;
        RECT 44.020 143.155 44.850 143.455 ;
        RECT 45.380 143.425 45.700 144.385 ;
        RECT 42.605 142.755 42.940 142.925 ;
        RECT 43.135 142.755 43.810 142.925 ;
        RECT 44.130 142.475 44.500 142.975 ;
        RECT 44.680 142.925 44.850 143.155 ;
        RECT 45.235 143.095 45.700 143.425 ;
        RECT 45.870 143.715 46.040 144.555 ;
        RECT 46.220 144.525 46.535 145.025 ;
        RECT 46.765 144.295 47.105 144.855 ;
        RECT 46.210 143.920 47.105 144.295 ;
        RECT 47.275 144.015 47.445 145.025 ;
        RECT 46.915 143.715 47.105 143.920 ;
        RECT 47.615 143.965 47.945 144.810 ;
        RECT 48.175 144.470 48.780 145.025 ;
        RECT 48.955 144.515 49.435 144.855 ;
        RECT 49.605 144.480 49.860 145.025 ;
        RECT 48.175 144.370 48.790 144.470 ;
        RECT 48.605 144.345 48.790 144.370 ;
        RECT 47.615 143.885 48.005 143.965 ;
        RECT 47.790 143.835 48.005 143.885 ;
        RECT 45.870 143.385 46.745 143.715 ;
        RECT 46.915 143.385 47.665 143.715 ;
        RECT 45.870 142.925 46.040 143.385 ;
        RECT 46.915 143.215 47.115 143.385 ;
        RECT 47.835 143.255 48.005 143.835 ;
        RECT 48.175 143.750 48.435 144.200 ;
        RECT 48.605 144.100 48.935 144.345 ;
        RECT 49.105 144.025 49.860 144.275 ;
        RECT 50.030 144.155 50.305 144.855 ;
        RECT 49.090 143.990 49.860 144.025 ;
        RECT 49.075 143.980 49.860 143.990 ;
        RECT 49.070 143.965 49.965 143.980 ;
        RECT 49.050 143.950 49.965 143.965 ;
        RECT 49.030 143.940 49.965 143.950 ;
        RECT 49.005 143.930 49.965 143.940 ;
        RECT 48.935 143.900 49.965 143.930 ;
        RECT 48.915 143.870 49.965 143.900 ;
        RECT 48.895 143.840 49.965 143.870 ;
        RECT 48.865 143.815 49.965 143.840 ;
        RECT 48.830 143.780 49.965 143.815 ;
        RECT 48.800 143.775 49.965 143.780 ;
        RECT 48.800 143.770 49.190 143.775 ;
        RECT 48.800 143.760 49.165 143.770 ;
        RECT 48.800 143.755 49.150 143.760 ;
        RECT 48.800 143.750 49.135 143.755 ;
        RECT 48.175 143.745 49.135 143.750 ;
        RECT 48.175 143.735 49.125 143.745 ;
        RECT 48.175 143.730 49.115 143.735 ;
        RECT 48.175 143.720 49.105 143.730 ;
        RECT 48.175 143.710 49.100 143.720 ;
        RECT 48.175 143.705 49.095 143.710 ;
        RECT 48.175 143.690 49.085 143.705 ;
        RECT 48.175 143.675 49.080 143.690 ;
        RECT 48.175 143.650 49.070 143.675 ;
        RECT 48.175 143.580 49.065 143.650 ;
        RECT 47.780 143.215 48.005 143.255 ;
        RECT 44.680 142.755 45.085 142.925 ;
        RECT 45.255 142.755 46.040 142.925 ;
        RECT 46.315 142.475 46.525 143.005 ;
        RECT 46.785 142.690 47.115 143.215 ;
        RECT 47.625 143.130 48.005 143.215 ;
        RECT 47.285 142.475 47.455 143.085 ;
        RECT 47.625 142.695 47.955 143.130 ;
        RECT 48.175 143.025 48.725 143.410 ;
        RECT 48.895 142.855 49.065 143.580 ;
        RECT 48.175 142.685 49.065 142.855 ;
        RECT 49.235 143.180 49.565 143.605 ;
        RECT 49.735 143.380 49.965 143.775 ;
        RECT 49.235 142.695 49.455 143.180 ;
        RECT 50.135 143.125 50.305 144.155 ;
        RECT 51.580 144.055 51.970 144.230 ;
        RECT 52.455 144.225 52.785 145.025 ;
        RECT 52.955 144.235 53.490 144.855 ;
        RECT 53.695 144.470 54.300 145.025 ;
        RECT 54.475 144.515 54.955 144.855 ;
        RECT 55.125 144.480 55.380 145.025 ;
        RECT 53.695 144.370 54.310 144.470 ;
        RECT 51.580 143.885 53.005 144.055 ;
        RECT 51.455 143.155 51.810 143.715 ;
        RECT 49.625 142.475 49.875 143.015 ;
        RECT 50.045 142.645 50.305 143.125 ;
        RECT 51.980 142.985 52.150 143.885 ;
        RECT 52.320 143.155 52.585 143.715 ;
        RECT 52.835 143.385 53.005 143.885 ;
        RECT 53.175 143.215 53.490 144.235 ;
        RECT 54.125 144.345 54.310 144.370 ;
        RECT 53.695 143.750 53.955 144.200 ;
        RECT 54.125 144.100 54.455 144.345 ;
        RECT 54.625 144.025 55.380 144.275 ;
        RECT 55.550 144.155 55.825 144.855 ;
        RECT 54.610 143.990 55.380 144.025 ;
        RECT 54.595 143.980 55.380 143.990 ;
        RECT 54.590 143.965 55.485 143.980 ;
        RECT 54.570 143.950 55.485 143.965 ;
        RECT 54.550 143.940 55.485 143.950 ;
        RECT 54.525 143.930 55.485 143.940 ;
        RECT 54.455 143.900 55.485 143.930 ;
        RECT 54.435 143.870 55.485 143.900 ;
        RECT 54.415 143.840 55.485 143.870 ;
        RECT 54.385 143.815 55.485 143.840 ;
        RECT 54.350 143.780 55.485 143.815 ;
        RECT 54.320 143.775 55.485 143.780 ;
        RECT 54.320 143.770 54.710 143.775 ;
        RECT 54.320 143.760 54.685 143.770 ;
        RECT 54.320 143.755 54.670 143.760 ;
        RECT 54.320 143.750 54.655 143.755 ;
        RECT 53.695 143.745 54.655 143.750 ;
        RECT 53.695 143.735 54.645 143.745 ;
        RECT 53.695 143.730 54.635 143.735 ;
        RECT 53.695 143.720 54.625 143.730 ;
        RECT 53.695 143.710 54.620 143.720 ;
        RECT 53.695 143.705 54.615 143.710 ;
        RECT 53.695 143.690 54.605 143.705 ;
        RECT 53.695 143.675 54.600 143.690 ;
        RECT 53.695 143.650 54.590 143.675 ;
        RECT 53.695 143.580 54.585 143.650 ;
        RECT 51.560 142.475 51.800 142.985 ;
        RECT 51.980 142.655 52.260 142.985 ;
        RECT 52.490 142.475 52.705 142.985 ;
        RECT 52.875 142.645 53.490 143.215 ;
        RECT 53.695 143.025 54.245 143.410 ;
        RECT 54.415 142.855 54.585 143.580 ;
        RECT 53.695 142.685 54.585 142.855 ;
        RECT 54.755 143.180 55.085 143.605 ;
        RECT 55.255 143.380 55.485 143.775 ;
        RECT 54.755 142.695 54.975 143.180 ;
        RECT 55.655 143.125 55.825 144.155 ;
        RECT 55.995 143.860 56.285 145.025 ;
        RECT 56.545 144.355 56.715 144.855 ;
        RECT 56.885 144.525 57.215 145.025 ;
        RECT 56.545 144.185 57.210 144.355 ;
        RECT 56.460 143.365 56.810 144.015 ;
        RECT 55.145 142.475 55.395 143.015 ;
        RECT 55.565 142.645 55.825 143.125 ;
        RECT 55.995 142.475 56.285 143.200 ;
        RECT 56.980 143.195 57.210 144.185 ;
        RECT 56.545 143.025 57.210 143.195 ;
        RECT 56.545 142.735 56.715 143.025 ;
        RECT 56.885 142.475 57.215 142.855 ;
        RECT 57.385 142.735 57.570 144.855 ;
        RECT 57.810 144.565 58.075 145.025 ;
        RECT 58.245 144.430 58.495 144.855 ;
        RECT 58.705 144.580 59.810 144.750 ;
        RECT 58.190 144.300 58.495 144.430 ;
        RECT 57.740 143.105 58.020 144.055 ;
        RECT 58.190 143.195 58.360 144.300 ;
        RECT 58.530 143.515 58.770 144.110 ;
        RECT 58.940 144.045 59.470 144.410 ;
        RECT 58.940 143.345 59.110 144.045 ;
        RECT 59.640 143.965 59.810 144.580 ;
        RECT 59.980 144.225 60.150 145.025 ;
        RECT 60.320 144.525 60.570 144.855 ;
        RECT 60.795 144.555 61.680 144.725 ;
        RECT 59.640 143.875 60.150 143.965 ;
        RECT 58.190 143.065 58.415 143.195 ;
        RECT 58.585 143.125 59.110 143.345 ;
        RECT 59.280 143.705 60.150 143.875 ;
        RECT 57.825 142.475 58.075 142.935 ;
        RECT 58.245 142.925 58.415 143.065 ;
        RECT 59.280 142.925 59.450 143.705 ;
        RECT 59.980 143.635 60.150 143.705 ;
        RECT 59.660 143.455 59.860 143.485 ;
        RECT 60.320 143.455 60.490 144.525 ;
        RECT 60.660 143.635 60.850 144.355 ;
        RECT 59.660 143.155 60.490 143.455 ;
        RECT 61.020 143.425 61.340 144.385 ;
        RECT 58.245 142.755 58.580 142.925 ;
        RECT 58.775 142.755 59.450 142.925 ;
        RECT 59.770 142.475 60.140 142.975 ;
        RECT 60.320 142.925 60.490 143.155 ;
        RECT 60.875 143.095 61.340 143.425 ;
        RECT 61.510 143.715 61.680 144.555 ;
        RECT 61.860 144.525 62.175 145.025 ;
        RECT 62.405 144.295 62.745 144.855 ;
        RECT 61.850 143.920 62.745 144.295 ;
        RECT 62.915 144.015 63.085 145.025 ;
        RECT 62.555 143.715 62.745 143.920 ;
        RECT 63.255 143.965 63.585 144.810 ;
        RECT 63.815 144.590 69.160 145.025 ;
        RECT 63.255 143.885 63.645 143.965 ;
        RECT 63.430 143.835 63.645 143.885 ;
        RECT 61.510 143.385 62.385 143.715 ;
        RECT 62.555 143.385 63.305 143.715 ;
        RECT 61.510 142.925 61.680 143.385 ;
        RECT 62.555 143.215 62.755 143.385 ;
        RECT 63.475 143.255 63.645 143.835 ;
        RECT 63.420 143.215 63.645 143.255 ;
        RECT 60.320 142.755 60.725 142.925 ;
        RECT 60.895 142.755 61.680 142.925 ;
        RECT 61.955 142.475 62.165 143.005 ;
        RECT 62.425 142.690 62.755 143.215 ;
        RECT 63.265 143.130 63.645 143.215 ;
        RECT 62.925 142.475 63.095 143.085 ;
        RECT 63.265 142.695 63.595 143.130 ;
        RECT 65.400 143.020 65.740 143.850 ;
        RECT 67.220 143.340 67.570 144.590 ;
        RECT 69.335 143.935 71.925 145.025 ;
        RECT 72.185 144.355 72.355 144.855 ;
        RECT 72.525 144.525 72.855 145.025 ;
        RECT 72.185 144.185 72.850 144.355 ;
        RECT 69.335 143.245 70.545 143.765 ;
        RECT 70.715 143.415 71.925 143.935 ;
        RECT 72.100 143.365 72.450 144.015 ;
        RECT 63.815 142.475 69.160 143.020 ;
        RECT 69.335 142.475 71.925 143.245 ;
        RECT 72.620 143.195 72.850 144.185 ;
        RECT 72.185 143.025 72.850 143.195 ;
        RECT 72.185 142.735 72.355 143.025 ;
        RECT 72.525 142.475 72.855 142.855 ;
        RECT 73.025 142.735 73.210 144.855 ;
        RECT 73.450 144.565 73.715 145.025 ;
        RECT 73.885 144.430 74.135 144.855 ;
        RECT 74.345 144.580 75.450 144.750 ;
        RECT 73.830 144.300 74.135 144.430 ;
        RECT 73.380 143.105 73.660 144.055 ;
        RECT 73.830 143.195 74.000 144.300 ;
        RECT 74.170 143.515 74.410 144.110 ;
        RECT 74.580 144.045 75.110 144.410 ;
        RECT 74.580 143.345 74.750 144.045 ;
        RECT 75.280 143.965 75.450 144.580 ;
        RECT 75.620 144.225 75.790 145.025 ;
        RECT 75.960 144.525 76.210 144.855 ;
        RECT 76.435 144.555 77.320 144.725 ;
        RECT 75.280 143.875 75.790 143.965 ;
        RECT 73.830 143.065 74.055 143.195 ;
        RECT 74.225 143.125 74.750 143.345 ;
        RECT 74.920 143.705 75.790 143.875 ;
        RECT 73.465 142.475 73.715 142.935 ;
        RECT 73.885 142.925 74.055 143.065 ;
        RECT 74.920 142.925 75.090 143.705 ;
        RECT 75.620 143.635 75.790 143.705 ;
        RECT 75.300 143.455 75.500 143.485 ;
        RECT 75.960 143.455 76.130 144.525 ;
        RECT 76.300 143.635 76.490 144.355 ;
        RECT 75.300 143.155 76.130 143.455 ;
        RECT 76.660 143.425 76.980 144.385 ;
        RECT 73.885 142.755 74.220 142.925 ;
        RECT 74.415 142.755 75.090 142.925 ;
        RECT 75.410 142.475 75.780 142.975 ;
        RECT 75.960 142.925 76.130 143.155 ;
        RECT 76.515 143.095 76.980 143.425 ;
        RECT 77.150 143.715 77.320 144.555 ;
        RECT 77.500 144.525 77.815 145.025 ;
        RECT 78.045 144.295 78.385 144.855 ;
        RECT 77.490 143.920 78.385 144.295 ;
        RECT 78.555 144.015 78.725 145.025 ;
        RECT 78.195 143.715 78.385 143.920 ;
        RECT 78.895 143.965 79.225 144.810 ;
        RECT 78.895 143.885 79.285 143.965 ;
        RECT 79.460 143.885 79.780 145.025 ;
        RECT 79.070 143.835 79.285 143.885 ;
        RECT 77.150 143.385 78.025 143.715 ;
        RECT 78.195 143.385 78.945 143.715 ;
        RECT 77.150 142.925 77.320 143.385 ;
        RECT 78.195 143.215 78.395 143.385 ;
        RECT 79.115 143.255 79.285 143.835 ;
        RECT 79.960 143.715 80.155 144.765 ;
        RECT 80.335 144.175 80.665 144.855 ;
        RECT 80.865 144.225 81.120 145.025 ;
        RECT 80.335 143.895 80.685 144.175 ;
        RECT 79.520 143.665 79.780 143.715 ;
        RECT 79.515 143.495 79.780 143.665 ;
        RECT 79.520 143.385 79.780 143.495 ;
        RECT 79.960 143.385 80.345 143.715 ;
        RECT 80.515 143.515 80.685 143.895 ;
        RECT 80.875 143.685 81.120 144.045 ;
        RECT 81.755 143.860 82.045 145.025 ;
        RECT 82.215 143.885 82.600 144.855 ;
        RECT 82.770 144.565 83.095 145.025 ;
        RECT 83.615 144.395 83.895 144.855 ;
        RECT 82.770 144.175 83.895 144.395 ;
        RECT 80.515 143.345 81.035 143.515 ;
        RECT 79.060 143.215 79.285 143.255 ;
        RECT 75.960 142.755 76.365 142.925 ;
        RECT 76.535 142.755 77.320 142.925 ;
        RECT 77.595 142.475 77.805 143.005 ;
        RECT 78.065 142.690 78.395 143.215 ;
        RECT 78.905 143.130 79.285 143.215 ;
        RECT 78.565 142.475 78.735 143.085 ;
        RECT 78.905 142.695 79.235 143.130 ;
        RECT 79.460 143.005 80.675 143.175 ;
        RECT 79.460 142.655 79.750 143.005 ;
        RECT 79.945 142.475 80.275 142.835 ;
        RECT 80.445 142.700 80.675 143.005 ;
        RECT 80.865 142.780 81.035 143.345 ;
        RECT 82.215 143.215 82.495 143.885 ;
        RECT 82.770 143.715 83.220 144.175 ;
        RECT 84.085 144.005 84.485 144.855 ;
        RECT 84.885 144.565 85.155 145.025 ;
        RECT 85.325 144.395 85.610 144.855 ;
        RECT 82.665 143.385 83.220 143.715 ;
        RECT 83.390 143.445 84.485 144.005 ;
        RECT 82.770 143.275 83.220 143.385 ;
        RECT 81.755 142.475 82.045 143.200 ;
        RECT 82.215 142.645 82.600 143.215 ;
        RECT 82.770 143.105 83.895 143.275 ;
        RECT 82.770 142.475 83.095 142.935 ;
        RECT 83.615 142.645 83.895 143.105 ;
        RECT 84.085 142.645 84.485 143.445 ;
        RECT 84.655 144.175 85.610 144.395 ;
        RECT 84.655 143.275 84.865 144.175 ;
        RECT 85.035 143.445 85.725 144.005 ;
        RECT 85.895 143.885 86.175 145.025 ;
        RECT 86.345 143.875 86.675 144.855 ;
        RECT 86.845 143.885 87.105 145.025 ;
        RECT 88.285 144.355 88.455 144.855 ;
        RECT 88.625 144.525 88.955 145.025 ;
        RECT 88.285 144.185 88.950 144.355 ;
        RECT 85.905 143.445 86.240 143.715 ;
        RECT 86.410 143.325 86.580 143.875 ;
        RECT 86.750 143.465 87.085 143.715 ;
        RECT 88.200 143.365 88.550 144.015 ;
        RECT 86.410 143.275 86.585 143.325 ;
        RECT 84.655 143.105 85.610 143.275 ;
        RECT 84.885 142.475 85.155 142.935 ;
        RECT 85.325 142.645 85.610 143.105 ;
        RECT 85.895 142.475 86.205 143.275 ;
        RECT 86.410 142.645 87.105 143.275 ;
        RECT 88.720 143.195 88.950 144.185 ;
        RECT 88.285 143.025 88.950 143.195 ;
        RECT 88.285 142.735 88.455 143.025 ;
        RECT 88.625 142.475 88.955 142.855 ;
        RECT 89.125 142.735 89.310 144.855 ;
        RECT 89.550 144.565 89.815 145.025 ;
        RECT 89.985 144.430 90.235 144.855 ;
        RECT 90.445 144.580 91.550 144.750 ;
        RECT 89.930 144.300 90.235 144.430 ;
        RECT 89.480 143.105 89.760 144.055 ;
        RECT 89.930 143.195 90.100 144.300 ;
        RECT 90.270 143.515 90.510 144.110 ;
        RECT 90.680 144.045 91.210 144.410 ;
        RECT 90.680 143.345 90.850 144.045 ;
        RECT 91.380 143.965 91.550 144.580 ;
        RECT 91.720 144.225 91.890 145.025 ;
        RECT 92.060 144.525 92.310 144.855 ;
        RECT 92.535 144.555 93.420 144.725 ;
        RECT 91.380 143.875 91.890 143.965 ;
        RECT 89.930 143.065 90.155 143.195 ;
        RECT 90.325 143.125 90.850 143.345 ;
        RECT 91.020 143.705 91.890 143.875 ;
        RECT 89.565 142.475 89.815 142.935 ;
        RECT 89.985 142.925 90.155 143.065 ;
        RECT 91.020 142.925 91.190 143.705 ;
        RECT 91.720 143.635 91.890 143.705 ;
        RECT 91.400 143.455 91.600 143.485 ;
        RECT 92.060 143.455 92.230 144.525 ;
        RECT 92.400 143.635 92.590 144.355 ;
        RECT 91.400 143.155 92.230 143.455 ;
        RECT 92.760 143.425 93.080 144.385 ;
        RECT 89.985 142.755 90.320 142.925 ;
        RECT 90.515 142.755 91.190 142.925 ;
        RECT 91.510 142.475 91.880 142.975 ;
        RECT 92.060 142.925 92.230 143.155 ;
        RECT 92.615 143.095 93.080 143.425 ;
        RECT 93.250 143.715 93.420 144.555 ;
        RECT 93.600 144.525 93.915 145.025 ;
        RECT 94.145 144.295 94.485 144.855 ;
        RECT 93.590 143.920 94.485 144.295 ;
        RECT 94.655 144.015 94.825 145.025 ;
        RECT 94.295 143.715 94.485 143.920 ;
        RECT 94.995 143.965 95.325 144.810 ;
        RECT 94.995 143.885 95.385 143.965 ;
        RECT 95.555 143.935 96.765 145.025 ;
        RECT 95.170 143.835 95.385 143.885 ;
        RECT 93.250 143.385 94.125 143.715 ;
        RECT 94.295 143.385 95.045 143.715 ;
        RECT 93.250 142.925 93.420 143.385 ;
        RECT 94.295 143.215 94.495 143.385 ;
        RECT 95.215 143.255 95.385 143.835 ;
        RECT 95.160 143.215 95.385 143.255 ;
        RECT 92.060 142.755 92.465 142.925 ;
        RECT 92.635 142.755 93.420 142.925 ;
        RECT 93.695 142.475 93.905 143.005 ;
        RECT 94.165 142.690 94.495 143.215 ;
        RECT 95.005 143.130 95.385 143.215 ;
        RECT 95.555 143.225 96.075 143.765 ;
        RECT 96.245 143.395 96.765 143.935 ;
        RECT 96.940 144.075 97.205 144.845 ;
        RECT 97.375 144.305 97.705 145.025 ;
        RECT 97.895 144.485 98.155 144.845 ;
        RECT 98.325 144.655 98.655 145.025 ;
        RECT 98.825 144.485 99.085 144.845 ;
        RECT 97.895 144.255 99.085 144.485 ;
        RECT 99.655 144.075 99.945 144.845 ;
        RECT 94.665 142.475 94.835 143.085 ;
        RECT 95.005 142.695 95.335 143.130 ;
        RECT 95.555 142.475 96.765 143.225 ;
        RECT 96.940 142.655 97.275 144.075 ;
        RECT 97.450 143.895 99.945 144.075 ;
        RECT 100.155 143.935 102.745 145.025 ;
        RECT 97.450 143.205 97.675 143.895 ;
        RECT 97.875 143.385 98.155 143.715 ;
        RECT 98.335 143.385 98.910 143.715 ;
        RECT 99.090 143.385 99.525 143.715 ;
        RECT 99.705 143.385 99.975 143.715 ;
        RECT 100.155 143.245 101.365 143.765 ;
        RECT 101.535 143.415 102.745 143.935 ;
        RECT 103.380 143.885 103.715 144.855 ;
        RECT 103.885 143.885 104.055 145.025 ;
        RECT 104.225 144.685 106.255 144.855 ;
        RECT 97.450 143.015 99.935 143.205 ;
        RECT 97.455 142.475 98.200 142.845 ;
        RECT 98.765 142.655 99.020 143.015 ;
        RECT 99.200 142.475 99.530 142.845 ;
        RECT 99.710 142.655 99.935 143.015 ;
        RECT 100.155 142.475 102.745 143.245 ;
        RECT 103.380 143.215 103.550 143.885 ;
        RECT 104.225 143.715 104.395 144.685 ;
        RECT 103.720 143.385 103.975 143.715 ;
        RECT 104.200 143.385 104.395 143.715 ;
        RECT 104.565 144.345 105.690 144.515 ;
        RECT 103.805 143.215 103.975 143.385 ;
        RECT 104.565 143.215 104.735 144.345 ;
        RECT 103.380 142.645 103.635 143.215 ;
        RECT 103.805 143.045 104.735 143.215 ;
        RECT 104.905 144.005 105.915 144.175 ;
        RECT 104.905 143.205 105.075 144.005 ;
        RECT 105.280 143.665 105.555 143.805 ;
        RECT 105.275 143.495 105.555 143.665 ;
        RECT 104.560 143.010 104.735 143.045 ;
        RECT 103.805 142.475 104.135 142.875 ;
        RECT 104.560 142.645 105.090 143.010 ;
        RECT 105.280 142.645 105.555 143.495 ;
        RECT 105.725 142.645 105.915 144.005 ;
        RECT 106.085 144.020 106.255 144.685 ;
        RECT 106.425 144.265 106.595 145.025 ;
        RECT 106.830 144.265 107.345 144.675 ;
        RECT 106.085 143.830 106.835 144.020 ;
        RECT 107.005 143.455 107.345 144.265 ;
        RECT 107.515 143.860 107.805 145.025 ;
        RECT 107.980 143.885 108.315 144.855 ;
        RECT 108.485 143.885 108.655 145.025 ;
        RECT 108.825 144.685 110.855 144.855 ;
        RECT 106.115 143.285 107.345 143.455 ;
        RECT 106.095 142.475 106.605 143.010 ;
        RECT 106.825 142.680 107.070 143.285 ;
        RECT 107.980 143.215 108.150 143.885 ;
        RECT 108.825 143.715 108.995 144.685 ;
        RECT 108.320 143.385 108.575 143.715 ;
        RECT 108.800 143.385 108.995 143.715 ;
        RECT 109.165 144.345 110.290 144.515 ;
        RECT 108.405 143.215 108.575 143.385 ;
        RECT 109.165 143.215 109.335 144.345 ;
        RECT 107.515 142.475 107.805 143.200 ;
        RECT 107.980 142.645 108.235 143.215 ;
        RECT 108.405 143.045 109.335 143.215 ;
        RECT 109.505 144.005 110.515 144.175 ;
        RECT 109.505 143.205 109.675 144.005 ;
        RECT 109.160 143.010 109.335 143.045 ;
        RECT 108.405 142.475 108.735 142.875 ;
        RECT 109.160 142.645 109.690 143.010 ;
        RECT 109.880 142.985 110.155 143.805 ;
        RECT 109.875 142.815 110.155 142.985 ;
        RECT 109.880 142.645 110.155 142.815 ;
        RECT 110.325 142.645 110.515 144.005 ;
        RECT 110.685 144.020 110.855 144.685 ;
        RECT 111.025 144.265 111.195 145.025 ;
        RECT 111.430 144.265 111.945 144.675 ;
        RECT 112.115 144.590 117.460 145.025 ;
        RECT 110.685 143.830 111.435 144.020 ;
        RECT 111.605 143.455 111.945 144.265 ;
        RECT 110.715 143.285 111.945 143.455 ;
        RECT 110.695 142.475 111.205 143.010 ;
        RECT 111.425 142.680 111.670 143.285 ;
        RECT 113.700 143.020 114.040 143.850 ;
        RECT 115.520 143.340 115.870 144.590 ;
        RECT 118.615 143.965 118.945 144.810 ;
        RECT 119.115 144.015 119.285 145.025 ;
        RECT 119.455 144.295 119.795 144.855 ;
        RECT 120.025 144.525 120.340 145.025 ;
        RECT 120.520 144.555 121.405 144.725 ;
        RECT 118.555 143.885 118.945 143.965 ;
        RECT 119.455 143.920 120.350 144.295 ;
        RECT 118.555 143.835 118.770 143.885 ;
        RECT 118.555 143.255 118.725 143.835 ;
        RECT 119.455 143.715 119.645 143.920 ;
        RECT 120.520 143.715 120.690 144.555 ;
        RECT 121.630 144.525 121.880 144.855 ;
        RECT 118.895 143.385 119.645 143.715 ;
        RECT 119.815 143.385 120.690 143.715 ;
        RECT 118.555 143.215 118.780 143.255 ;
        RECT 119.445 143.215 119.645 143.385 ;
        RECT 118.555 143.130 118.935 143.215 ;
        RECT 112.115 142.475 117.460 143.020 ;
        RECT 118.605 142.695 118.935 143.130 ;
        RECT 119.105 142.475 119.275 143.085 ;
        RECT 119.445 142.690 119.775 143.215 ;
        RECT 120.035 142.475 120.245 143.005 ;
        RECT 120.520 142.925 120.690 143.385 ;
        RECT 120.860 143.425 121.180 144.385 ;
        RECT 121.350 143.635 121.540 144.355 ;
        RECT 121.710 143.455 121.880 144.525 ;
        RECT 122.050 144.225 122.220 145.025 ;
        RECT 122.390 144.580 123.495 144.750 ;
        RECT 122.390 143.965 122.560 144.580 ;
        RECT 123.705 144.430 123.955 144.855 ;
        RECT 124.125 144.565 124.390 145.025 ;
        RECT 122.730 144.045 123.260 144.410 ;
        RECT 123.705 144.300 124.010 144.430 ;
        RECT 122.050 143.875 122.560 143.965 ;
        RECT 122.050 143.705 122.920 143.875 ;
        RECT 122.050 143.635 122.220 143.705 ;
        RECT 122.340 143.455 122.540 143.485 ;
        RECT 120.860 143.095 121.325 143.425 ;
        RECT 121.710 143.155 122.540 143.455 ;
        RECT 121.710 142.925 121.880 143.155 ;
        RECT 120.520 142.755 121.305 142.925 ;
        RECT 121.475 142.755 121.880 142.925 ;
        RECT 122.060 142.475 122.430 142.975 ;
        RECT 122.750 142.925 122.920 143.705 ;
        RECT 123.090 143.345 123.260 144.045 ;
        RECT 123.430 143.515 123.670 144.110 ;
        RECT 123.090 143.125 123.615 143.345 ;
        RECT 123.840 143.195 124.010 144.300 ;
        RECT 123.785 143.065 124.010 143.195 ;
        RECT 124.180 143.105 124.460 144.055 ;
        RECT 123.785 142.925 123.955 143.065 ;
        RECT 122.750 142.755 123.425 142.925 ;
        RECT 123.620 142.755 123.955 142.925 ;
        RECT 124.125 142.475 124.375 142.935 ;
        RECT 124.630 142.735 124.815 144.855 ;
        RECT 124.985 144.525 125.315 145.025 ;
        RECT 125.485 144.355 125.655 144.855 ;
        RECT 124.990 144.185 125.655 144.355 ;
        RECT 126.030 144.395 126.315 144.855 ;
        RECT 126.485 144.565 126.755 145.025 ;
        RECT 124.990 143.195 125.220 144.185 ;
        RECT 126.030 144.175 126.985 144.395 ;
        RECT 125.390 143.365 125.740 144.015 ;
        RECT 125.915 143.445 126.605 144.005 ;
        RECT 126.775 143.275 126.985 144.175 ;
        RECT 124.990 143.025 125.655 143.195 ;
        RECT 124.985 142.475 125.315 142.855 ;
        RECT 125.485 142.735 125.655 143.025 ;
        RECT 126.030 143.105 126.985 143.275 ;
        RECT 127.155 144.005 127.555 144.855 ;
        RECT 127.745 144.395 128.025 144.855 ;
        RECT 128.545 144.565 128.870 145.025 ;
        RECT 127.745 144.175 128.870 144.395 ;
        RECT 127.155 143.445 128.250 144.005 ;
        RECT 128.420 143.715 128.870 144.175 ;
        RECT 129.040 143.885 129.425 144.855 ;
        RECT 129.595 143.935 133.105 145.025 ;
        RECT 126.030 142.645 126.315 143.105 ;
        RECT 126.485 142.475 126.755 142.935 ;
        RECT 127.155 142.645 127.555 143.445 ;
        RECT 128.420 143.385 128.975 143.715 ;
        RECT 128.420 143.275 128.870 143.385 ;
        RECT 127.745 143.105 128.870 143.275 ;
        RECT 129.145 143.215 129.425 143.885 ;
        RECT 127.745 142.645 128.025 143.105 ;
        RECT 128.545 142.475 128.870 142.935 ;
        RECT 129.040 142.645 129.425 143.215 ;
        RECT 129.595 143.245 131.245 143.765 ;
        RECT 131.415 143.415 133.105 143.935 ;
        RECT 133.275 143.860 133.565 145.025 ;
        RECT 133.825 144.355 133.995 144.855 ;
        RECT 134.165 144.525 134.495 145.025 ;
        RECT 133.825 144.185 134.490 144.355 ;
        RECT 133.740 143.365 134.090 144.015 ;
        RECT 129.595 142.475 133.105 143.245 ;
        RECT 133.275 142.475 133.565 143.200 ;
        RECT 134.260 143.195 134.490 144.185 ;
        RECT 133.825 143.025 134.490 143.195 ;
        RECT 133.825 142.735 133.995 143.025 ;
        RECT 134.165 142.475 134.495 142.855 ;
        RECT 134.665 142.735 134.850 144.855 ;
        RECT 135.090 144.565 135.355 145.025 ;
        RECT 135.525 144.430 135.775 144.855 ;
        RECT 135.985 144.580 137.090 144.750 ;
        RECT 135.470 144.300 135.775 144.430 ;
        RECT 135.020 143.105 135.300 144.055 ;
        RECT 135.470 143.195 135.640 144.300 ;
        RECT 135.810 143.515 136.050 144.110 ;
        RECT 136.220 144.045 136.750 144.410 ;
        RECT 136.220 143.345 136.390 144.045 ;
        RECT 136.920 143.965 137.090 144.580 ;
        RECT 137.260 144.225 137.430 145.025 ;
        RECT 137.600 144.525 137.850 144.855 ;
        RECT 138.075 144.555 138.960 144.725 ;
        RECT 136.920 143.875 137.430 143.965 ;
        RECT 135.470 143.065 135.695 143.195 ;
        RECT 135.865 143.125 136.390 143.345 ;
        RECT 136.560 143.705 137.430 143.875 ;
        RECT 135.105 142.475 135.355 142.935 ;
        RECT 135.525 142.925 135.695 143.065 ;
        RECT 136.560 142.925 136.730 143.705 ;
        RECT 137.260 143.635 137.430 143.705 ;
        RECT 136.940 143.455 137.140 143.485 ;
        RECT 137.600 143.455 137.770 144.525 ;
        RECT 137.940 143.635 138.130 144.355 ;
        RECT 136.940 143.155 137.770 143.455 ;
        RECT 138.300 143.425 138.620 144.385 ;
        RECT 135.525 142.755 135.860 142.925 ;
        RECT 136.055 142.755 136.730 142.925 ;
        RECT 137.050 142.475 137.420 142.975 ;
        RECT 137.600 142.925 137.770 143.155 ;
        RECT 138.155 143.095 138.620 143.425 ;
        RECT 138.790 143.715 138.960 144.555 ;
        RECT 139.140 144.525 139.455 145.025 ;
        RECT 139.685 144.295 140.025 144.855 ;
        RECT 139.130 143.920 140.025 144.295 ;
        RECT 140.195 144.015 140.365 145.025 ;
        RECT 139.835 143.715 140.025 143.920 ;
        RECT 140.535 143.965 140.865 144.810 ;
        RECT 140.535 143.885 140.925 143.965 ;
        RECT 140.710 143.835 140.925 143.885 ;
        RECT 138.790 143.385 139.665 143.715 ;
        RECT 139.835 143.385 140.585 143.715 ;
        RECT 138.790 142.925 138.960 143.385 ;
        RECT 139.835 143.215 140.035 143.385 ;
        RECT 140.755 143.255 140.925 143.835 ;
        RECT 140.700 143.215 140.925 143.255 ;
        RECT 137.600 142.755 138.005 142.925 ;
        RECT 138.175 142.755 138.960 142.925 ;
        RECT 139.235 142.475 139.445 143.005 ;
        RECT 139.705 142.690 140.035 143.215 ;
        RECT 140.545 143.130 140.925 143.215 ;
        RECT 141.095 143.885 141.480 144.855 ;
        RECT 141.650 144.565 141.975 145.025 ;
        RECT 142.495 144.395 142.775 144.855 ;
        RECT 141.650 144.175 142.775 144.395 ;
        RECT 141.095 143.215 141.375 143.885 ;
        RECT 141.650 143.715 142.100 144.175 ;
        RECT 142.965 144.005 143.365 144.855 ;
        RECT 143.765 144.565 144.035 145.025 ;
        RECT 144.205 144.395 144.490 144.855 ;
        RECT 141.545 143.385 142.100 143.715 ;
        RECT 142.270 143.445 143.365 144.005 ;
        RECT 141.650 143.275 142.100 143.385 ;
        RECT 140.205 142.475 140.375 143.085 ;
        RECT 140.545 142.695 140.875 143.130 ;
        RECT 141.095 142.645 141.480 143.215 ;
        RECT 141.650 143.105 142.775 143.275 ;
        RECT 141.650 142.475 141.975 142.935 ;
        RECT 142.495 142.645 142.775 143.105 ;
        RECT 142.965 142.645 143.365 143.445 ;
        RECT 143.535 144.175 144.490 144.395 ;
        RECT 143.535 143.275 143.745 144.175 ;
        RECT 143.915 143.445 144.605 144.005 ;
        RECT 145.695 143.935 146.905 145.025 ;
        RECT 145.695 143.395 146.215 143.935 ;
        RECT 143.535 143.105 144.490 143.275 ;
        RECT 146.385 143.225 146.905 143.765 ;
        RECT 143.765 142.475 144.035 142.935 ;
        RECT 144.205 142.645 144.490 143.105 ;
        RECT 145.695 142.475 146.905 143.225 ;
        RECT 17.270 142.305 146.990 142.475 ;
        RECT 17.355 141.555 18.565 142.305 ;
        RECT 19.285 141.755 19.455 142.045 ;
        RECT 19.625 141.925 19.955 142.305 ;
        RECT 19.285 141.585 19.950 141.755 ;
        RECT 17.355 141.015 17.875 141.555 ;
        RECT 18.045 140.845 18.565 141.385 ;
        RECT 17.355 139.755 18.565 140.845 ;
        RECT 19.200 140.765 19.550 141.415 ;
        RECT 19.720 140.595 19.950 141.585 ;
        RECT 19.285 140.425 19.950 140.595 ;
        RECT 19.285 139.925 19.455 140.425 ;
        RECT 19.625 139.755 19.955 140.255 ;
        RECT 20.125 139.925 20.310 142.045 ;
        RECT 20.565 141.845 20.815 142.305 ;
        RECT 20.985 141.855 21.320 142.025 ;
        RECT 21.515 141.855 22.190 142.025 ;
        RECT 20.985 141.715 21.155 141.855 ;
        RECT 20.480 140.725 20.760 141.675 ;
        RECT 20.930 141.585 21.155 141.715 ;
        RECT 20.930 140.480 21.100 141.585 ;
        RECT 21.325 141.435 21.850 141.655 ;
        RECT 21.270 140.670 21.510 141.265 ;
        RECT 21.680 140.735 21.850 141.435 ;
        RECT 22.020 141.075 22.190 141.855 ;
        RECT 22.510 141.805 22.880 142.305 ;
        RECT 23.060 141.855 23.465 142.025 ;
        RECT 23.635 141.855 24.420 142.025 ;
        RECT 23.060 141.625 23.230 141.855 ;
        RECT 22.400 141.325 23.230 141.625 ;
        RECT 23.615 141.355 24.080 141.685 ;
        RECT 22.400 141.295 22.600 141.325 ;
        RECT 22.720 141.075 22.890 141.145 ;
        RECT 22.020 140.905 22.890 141.075 ;
        RECT 22.380 140.815 22.890 140.905 ;
        RECT 20.930 140.350 21.235 140.480 ;
        RECT 21.680 140.370 22.210 140.735 ;
        RECT 20.550 139.755 20.815 140.215 ;
        RECT 20.985 139.925 21.235 140.350 ;
        RECT 22.380 140.200 22.550 140.815 ;
        RECT 21.445 140.030 22.550 140.200 ;
        RECT 22.720 139.755 22.890 140.555 ;
        RECT 23.060 140.255 23.230 141.325 ;
        RECT 23.400 140.425 23.590 141.145 ;
        RECT 23.760 140.395 24.080 141.355 ;
        RECT 24.250 141.395 24.420 141.855 ;
        RECT 24.695 141.775 24.905 142.305 ;
        RECT 25.165 141.565 25.495 142.090 ;
        RECT 25.665 141.695 25.835 142.305 ;
        RECT 26.005 141.650 26.335 142.085 ;
        RECT 27.640 141.795 27.880 142.305 ;
        RECT 28.060 141.795 28.340 142.125 ;
        RECT 28.570 141.795 28.785 142.305 ;
        RECT 26.005 141.565 26.385 141.650 ;
        RECT 25.295 141.395 25.495 141.565 ;
        RECT 26.160 141.525 26.385 141.565 ;
        RECT 24.250 141.065 25.125 141.395 ;
        RECT 25.295 141.065 26.045 141.395 ;
        RECT 23.060 139.925 23.310 140.255 ;
        RECT 24.250 140.225 24.420 141.065 ;
        RECT 25.295 140.860 25.485 141.065 ;
        RECT 26.215 140.945 26.385 141.525 ;
        RECT 27.535 141.065 27.890 141.625 ;
        RECT 26.170 140.895 26.385 140.945 ;
        RECT 28.060 140.895 28.230 141.795 ;
        RECT 28.400 141.065 28.665 141.625 ;
        RECT 28.955 141.565 29.570 142.135 ;
        RECT 29.775 141.760 35.120 142.305 ;
        RECT 28.915 140.895 29.085 141.395 ;
        RECT 24.590 140.485 25.485 140.860 ;
        RECT 25.995 140.815 26.385 140.895 ;
        RECT 23.535 140.055 24.420 140.225 ;
        RECT 24.600 139.755 24.915 140.255 ;
        RECT 25.145 139.925 25.485 140.485 ;
        RECT 25.655 139.755 25.825 140.765 ;
        RECT 25.995 139.970 26.325 140.815 ;
        RECT 27.660 140.725 29.085 140.895 ;
        RECT 27.660 140.550 28.050 140.725 ;
        RECT 28.535 139.755 28.865 140.555 ;
        RECT 29.255 140.545 29.570 141.565 ;
        RECT 31.360 140.930 31.700 141.760 ;
        RECT 35.845 141.755 36.015 142.045 ;
        RECT 36.185 141.925 36.515 142.305 ;
        RECT 35.845 141.585 36.510 141.755 ;
        RECT 29.035 139.925 29.570 140.545 ;
        RECT 33.180 140.190 33.530 141.440 ;
        RECT 35.760 140.765 36.110 141.415 ;
        RECT 36.280 140.595 36.510 141.585 ;
        RECT 35.845 140.425 36.510 140.595 ;
        RECT 29.775 139.755 35.120 140.190 ;
        RECT 35.845 139.925 36.015 140.425 ;
        RECT 36.185 139.755 36.515 140.255 ;
        RECT 36.685 139.925 36.870 142.045 ;
        RECT 37.125 141.845 37.375 142.305 ;
        RECT 37.545 141.855 37.880 142.025 ;
        RECT 38.075 141.855 38.750 142.025 ;
        RECT 37.545 141.715 37.715 141.855 ;
        RECT 37.040 140.725 37.320 141.675 ;
        RECT 37.490 141.585 37.715 141.715 ;
        RECT 37.490 140.480 37.660 141.585 ;
        RECT 37.885 141.435 38.410 141.655 ;
        RECT 37.830 140.670 38.070 141.265 ;
        RECT 38.240 140.735 38.410 141.435 ;
        RECT 38.580 141.075 38.750 141.855 ;
        RECT 39.070 141.805 39.440 142.305 ;
        RECT 39.620 141.855 40.025 142.025 ;
        RECT 40.195 141.855 40.980 142.025 ;
        RECT 39.620 141.625 39.790 141.855 ;
        RECT 38.960 141.325 39.790 141.625 ;
        RECT 40.175 141.355 40.640 141.685 ;
        RECT 38.960 141.295 39.160 141.325 ;
        RECT 39.280 141.075 39.450 141.145 ;
        RECT 38.580 140.905 39.450 141.075 ;
        RECT 38.940 140.815 39.450 140.905 ;
        RECT 37.490 140.350 37.795 140.480 ;
        RECT 38.240 140.370 38.770 140.735 ;
        RECT 37.110 139.755 37.375 140.215 ;
        RECT 37.545 139.925 37.795 140.350 ;
        RECT 38.940 140.200 39.110 140.815 ;
        RECT 38.005 140.030 39.110 140.200 ;
        RECT 39.280 139.755 39.450 140.555 ;
        RECT 39.620 140.255 39.790 141.325 ;
        RECT 39.960 140.425 40.150 141.145 ;
        RECT 40.320 140.395 40.640 141.355 ;
        RECT 40.810 141.395 40.980 141.855 ;
        RECT 41.255 141.775 41.465 142.305 ;
        RECT 41.725 141.565 42.055 142.090 ;
        RECT 42.225 141.695 42.395 142.305 ;
        RECT 42.565 141.650 42.895 142.085 ;
        RECT 42.565 141.565 42.945 141.650 ;
        RECT 43.115 141.580 43.405 142.305 ;
        RECT 41.855 141.395 42.055 141.565 ;
        RECT 42.720 141.525 42.945 141.565 ;
        RECT 40.810 141.065 41.685 141.395 ;
        RECT 41.855 141.065 42.605 141.395 ;
        RECT 39.620 139.925 39.870 140.255 ;
        RECT 40.810 140.225 40.980 141.065 ;
        RECT 41.855 140.860 42.045 141.065 ;
        RECT 42.775 140.945 42.945 141.525 ;
        RECT 43.575 141.505 44.270 142.135 ;
        RECT 44.475 141.505 44.785 142.305 ;
        RECT 44.955 141.760 50.300 142.305 ;
        RECT 43.595 141.065 43.930 141.315 ;
        RECT 42.730 140.895 42.945 140.945 ;
        RECT 41.150 140.485 42.045 140.860 ;
        RECT 42.555 140.815 42.945 140.895 ;
        RECT 40.095 140.055 40.980 140.225 ;
        RECT 41.160 139.755 41.475 140.255 ;
        RECT 41.705 139.925 42.045 140.485 ;
        RECT 42.215 139.755 42.385 140.765 ;
        RECT 42.555 139.970 42.885 140.815 ;
        RECT 43.115 139.755 43.405 140.920 ;
        RECT 44.100 140.905 44.270 141.505 ;
        RECT 44.440 141.065 44.775 141.335 ;
        RECT 46.540 140.930 46.880 141.760 ;
        RECT 51.445 141.650 51.775 142.085 ;
        RECT 51.945 141.695 52.115 142.305 ;
        RECT 51.395 141.565 51.775 141.650 ;
        RECT 52.285 141.565 52.615 142.090 ;
        RECT 52.875 141.775 53.085 142.305 ;
        RECT 53.360 141.855 54.145 142.025 ;
        RECT 54.315 141.855 54.720 142.025 ;
        RECT 51.395 141.525 51.620 141.565 ;
        RECT 43.575 139.755 43.835 140.895 ;
        RECT 44.005 139.925 44.335 140.905 ;
        RECT 44.505 139.755 44.785 140.895 ;
        RECT 48.360 140.190 48.710 141.440 ;
        RECT 51.395 140.945 51.565 141.525 ;
        RECT 52.285 141.395 52.485 141.565 ;
        RECT 53.360 141.395 53.530 141.855 ;
        RECT 51.735 141.065 52.485 141.395 ;
        RECT 52.655 141.065 53.530 141.395 ;
        RECT 51.395 140.895 51.610 140.945 ;
        RECT 51.395 140.815 51.785 140.895 ;
        RECT 44.955 139.755 50.300 140.190 ;
        RECT 51.455 139.970 51.785 140.815 ;
        RECT 52.295 140.860 52.485 141.065 ;
        RECT 51.955 139.755 52.125 140.765 ;
        RECT 52.295 140.485 53.190 140.860 ;
        RECT 52.295 139.925 52.635 140.485 ;
        RECT 52.865 139.755 53.180 140.255 ;
        RECT 53.360 140.225 53.530 141.065 ;
        RECT 53.700 141.355 54.165 141.685 ;
        RECT 54.550 141.625 54.720 141.855 ;
        RECT 54.900 141.805 55.270 142.305 ;
        RECT 55.590 141.855 56.265 142.025 ;
        RECT 56.460 141.855 56.795 142.025 ;
        RECT 53.700 140.395 54.020 141.355 ;
        RECT 54.550 141.325 55.380 141.625 ;
        RECT 54.190 140.425 54.380 141.145 ;
        RECT 54.550 140.255 54.720 141.325 ;
        RECT 55.180 141.295 55.380 141.325 ;
        RECT 54.890 141.075 55.060 141.145 ;
        RECT 55.590 141.075 55.760 141.855 ;
        RECT 56.625 141.715 56.795 141.855 ;
        RECT 56.965 141.845 57.215 142.305 ;
        RECT 54.890 140.905 55.760 141.075 ;
        RECT 55.930 141.435 56.455 141.655 ;
        RECT 56.625 141.585 56.850 141.715 ;
        RECT 54.890 140.815 55.400 140.905 ;
        RECT 53.360 140.055 54.245 140.225 ;
        RECT 54.470 139.925 54.720 140.255 ;
        RECT 54.890 139.755 55.060 140.555 ;
        RECT 55.230 140.200 55.400 140.815 ;
        RECT 55.930 140.735 56.100 141.435 ;
        RECT 55.570 140.370 56.100 140.735 ;
        RECT 56.270 140.670 56.510 141.265 ;
        RECT 56.680 140.480 56.850 141.585 ;
        RECT 57.020 140.725 57.300 141.675 ;
        RECT 56.545 140.350 56.850 140.480 ;
        RECT 55.230 140.030 56.335 140.200 ;
        RECT 56.545 139.925 56.795 140.350 ;
        RECT 56.965 139.755 57.230 140.215 ;
        RECT 57.470 139.925 57.655 142.045 ;
        RECT 57.825 141.925 58.155 142.305 ;
        RECT 58.325 141.755 58.495 142.045 ;
        RECT 58.755 141.760 64.100 142.305 ;
        RECT 57.830 141.585 58.495 141.755 ;
        RECT 57.830 140.595 58.060 141.585 ;
        RECT 58.230 140.765 58.580 141.415 ;
        RECT 60.340 140.930 60.680 141.760 ;
        RECT 64.275 141.555 65.485 142.305 ;
        RECT 65.700 141.845 65.965 142.305 ;
        RECT 66.335 141.665 66.505 142.135 ;
        RECT 66.755 141.845 66.925 142.305 ;
        RECT 67.175 141.665 67.345 142.135 ;
        RECT 67.595 141.845 67.765 142.305 ;
        RECT 68.015 141.665 68.185 142.135 ;
        RECT 68.355 141.840 68.605 142.305 ;
        RECT 57.830 140.425 58.495 140.595 ;
        RECT 57.825 139.755 58.155 140.255 ;
        RECT 58.325 139.925 58.495 140.425 ;
        RECT 62.160 140.190 62.510 141.440 ;
        RECT 64.275 141.015 64.795 141.555 ;
        RECT 66.335 141.485 68.705 141.665 ;
        RECT 68.875 141.580 69.165 142.305 ;
        RECT 69.395 141.845 69.640 142.305 ;
        RECT 64.965 140.845 65.485 141.385 ;
        RECT 65.675 141.065 68.185 141.315 ;
        RECT 68.355 140.895 68.705 141.485 ;
        RECT 69.335 141.065 69.650 141.675 ;
        RECT 69.820 141.315 70.070 142.125 ;
        RECT 70.240 141.780 70.500 142.305 ;
        RECT 70.670 141.655 70.930 142.110 ;
        RECT 71.100 141.825 71.360 142.305 ;
        RECT 71.530 141.655 71.790 142.110 ;
        RECT 71.960 141.825 72.220 142.305 ;
        RECT 72.390 141.655 72.650 142.110 ;
        RECT 72.820 141.825 73.080 142.305 ;
        RECT 73.250 141.655 73.510 142.110 ;
        RECT 73.680 141.825 73.980 142.305 ;
        RECT 70.670 141.485 73.980 141.655 ;
        RECT 69.820 141.065 72.840 141.315 ;
        RECT 58.755 139.755 64.100 140.190 ;
        RECT 64.275 139.755 65.485 140.845 ;
        RECT 65.700 139.755 65.995 140.895 ;
        RECT 66.255 140.725 68.705 140.895 ;
        RECT 66.255 139.925 66.585 140.725 ;
        RECT 66.755 139.755 66.925 140.555 ;
        RECT 67.095 139.925 67.425 140.725 ;
        RECT 67.935 140.705 68.705 140.725 ;
        RECT 67.595 139.755 67.765 140.555 ;
        RECT 67.935 139.925 68.265 140.705 ;
        RECT 68.435 139.755 68.605 140.215 ;
        RECT 68.875 139.755 69.165 140.920 ;
        RECT 69.345 139.755 69.640 140.865 ;
        RECT 69.820 139.930 70.070 141.065 ;
        RECT 73.010 140.895 73.980 141.485 ;
        RECT 74.395 141.535 76.985 142.305 ;
        RECT 77.160 141.815 77.415 142.305 ;
        RECT 77.585 141.795 78.815 142.135 ;
        RECT 74.395 141.015 75.605 141.535 ;
        RECT 70.240 139.755 70.500 140.865 ;
        RECT 70.670 140.655 73.980 140.895 ;
        RECT 75.775 140.845 76.985 141.365 ;
        RECT 77.180 141.065 77.400 141.645 ;
        RECT 77.585 140.895 77.765 141.795 ;
        RECT 77.935 141.065 78.310 141.625 ;
        RECT 78.485 141.565 78.815 141.795 ;
        RECT 78.995 141.760 84.340 142.305 ;
        RECT 78.515 141.065 78.825 141.395 ;
        RECT 80.580 140.930 80.920 141.760 ;
        RECT 85.015 141.485 85.245 142.305 ;
        RECT 85.415 141.505 85.745 142.135 ;
        RECT 70.670 139.930 70.930 140.655 ;
        RECT 71.100 139.755 71.360 140.485 ;
        RECT 71.530 139.930 71.790 140.655 ;
        RECT 71.960 139.755 72.220 140.485 ;
        RECT 72.390 139.930 72.650 140.655 ;
        RECT 72.820 139.755 73.080 140.485 ;
        RECT 73.250 139.930 73.510 140.655 ;
        RECT 73.680 139.755 73.975 140.485 ;
        RECT 74.395 139.755 76.985 140.845 ;
        RECT 77.160 139.755 77.415 140.895 ;
        RECT 77.585 140.725 78.815 140.895 ;
        RECT 77.585 139.925 77.915 140.725 ;
        RECT 78.085 139.755 78.315 140.555 ;
        RECT 78.485 139.925 78.815 140.725 ;
        RECT 82.400 140.190 82.750 141.440 ;
        RECT 84.995 141.065 85.325 141.315 ;
        RECT 85.495 140.905 85.745 141.505 ;
        RECT 85.915 141.485 86.125 142.305 ;
        RECT 86.355 141.925 87.245 142.095 ;
        RECT 86.355 141.370 86.905 141.755 ;
        RECT 87.075 141.200 87.245 141.925 ;
        RECT 78.995 139.755 84.340 140.190 ;
        RECT 85.015 139.755 85.245 140.895 ;
        RECT 85.415 139.925 85.745 140.905 ;
        RECT 86.355 141.130 87.245 141.200 ;
        RECT 87.415 141.600 87.635 142.085 ;
        RECT 87.805 141.765 88.055 142.305 ;
        RECT 88.225 141.655 88.485 142.135 ;
        RECT 87.415 141.175 87.745 141.600 ;
        RECT 86.355 141.105 87.250 141.130 ;
        RECT 86.355 141.090 87.260 141.105 ;
        RECT 86.355 141.075 87.265 141.090 ;
        RECT 86.355 141.070 87.275 141.075 ;
        RECT 86.355 141.060 87.280 141.070 ;
        RECT 86.355 141.050 87.285 141.060 ;
        RECT 86.355 141.045 87.295 141.050 ;
        RECT 86.355 141.035 87.305 141.045 ;
        RECT 86.355 141.030 87.315 141.035 ;
        RECT 85.915 139.755 86.125 140.895 ;
        RECT 86.355 140.580 86.615 141.030 ;
        RECT 86.980 141.025 87.315 141.030 ;
        RECT 86.980 141.020 87.330 141.025 ;
        RECT 86.980 141.010 87.345 141.020 ;
        RECT 86.980 141.005 87.370 141.010 ;
        RECT 87.915 141.005 88.145 141.400 ;
        RECT 86.980 141.000 88.145 141.005 ;
        RECT 87.010 140.965 88.145 141.000 ;
        RECT 87.045 140.940 88.145 140.965 ;
        RECT 87.075 140.910 88.145 140.940 ;
        RECT 87.095 140.880 88.145 140.910 ;
        RECT 87.115 140.850 88.145 140.880 ;
        RECT 87.185 140.840 88.145 140.850 ;
        RECT 87.210 140.830 88.145 140.840 ;
        RECT 87.230 140.815 88.145 140.830 ;
        RECT 87.250 140.800 88.145 140.815 ;
        RECT 87.255 140.790 88.040 140.800 ;
        RECT 87.270 140.755 88.040 140.790 ;
        RECT 86.785 140.435 87.115 140.680 ;
        RECT 87.285 140.505 88.040 140.755 ;
        RECT 88.315 140.625 88.485 141.655 ;
        RECT 86.785 140.410 86.970 140.435 ;
        RECT 86.355 140.310 86.970 140.410 ;
        RECT 86.355 139.755 86.960 140.310 ;
        RECT 87.135 139.925 87.615 140.265 ;
        RECT 87.785 139.755 88.040 140.300 ;
        RECT 88.210 139.925 88.485 140.625 ;
        RECT 89.120 141.565 89.375 142.135 ;
        RECT 89.545 141.905 89.875 142.305 ;
        RECT 90.300 141.770 90.830 142.135 ;
        RECT 91.020 141.965 91.295 142.135 ;
        RECT 91.015 141.795 91.295 141.965 ;
        RECT 90.300 141.735 90.475 141.770 ;
        RECT 89.545 141.565 90.475 141.735 ;
        RECT 89.120 140.895 89.290 141.565 ;
        RECT 89.545 141.395 89.715 141.565 ;
        RECT 89.460 141.065 89.715 141.395 ;
        RECT 89.940 141.065 90.135 141.395 ;
        RECT 89.120 139.925 89.455 140.895 ;
        RECT 89.625 139.755 89.795 140.895 ;
        RECT 89.965 140.095 90.135 141.065 ;
        RECT 90.305 140.435 90.475 141.565 ;
        RECT 90.645 140.775 90.815 141.575 ;
        RECT 91.020 140.975 91.295 141.795 ;
        RECT 91.465 140.775 91.655 142.135 ;
        RECT 91.835 141.770 92.345 142.305 ;
        RECT 92.565 141.495 92.810 142.100 ;
        RECT 93.255 141.555 94.465 142.305 ;
        RECT 94.635 141.580 94.925 142.305 ;
        RECT 95.095 141.760 100.440 142.305 ;
        RECT 91.855 141.325 93.085 141.495 ;
        RECT 90.645 140.605 91.655 140.775 ;
        RECT 91.825 140.760 92.575 140.950 ;
        RECT 90.305 140.265 91.430 140.435 ;
        RECT 91.825 140.095 91.995 140.760 ;
        RECT 92.745 140.515 93.085 141.325 ;
        RECT 93.255 141.015 93.775 141.555 ;
        RECT 93.945 140.845 94.465 141.385 ;
        RECT 96.680 140.930 97.020 141.760 ;
        RECT 100.615 141.535 102.285 142.305 ;
        RECT 102.570 141.675 102.855 142.135 ;
        RECT 103.025 141.845 103.295 142.305 ;
        RECT 89.965 139.925 91.995 140.095 ;
        RECT 92.165 139.755 92.335 140.515 ;
        RECT 92.570 140.105 93.085 140.515 ;
        RECT 93.255 139.755 94.465 140.845 ;
        RECT 94.635 139.755 94.925 140.920 ;
        RECT 98.500 140.190 98.850 141.440 ;
        RECT 100.615 141.015 101.365 141.535 ;
        RECT 102.570 141.505 103.525 141.675 ;
        RECT 101.535 140.845 102.285 141.365 ;
        RECT 95.095 139.755 100.440 140.190 ;
        RECT 100.615 139.755 102.285 140.845 ;
        RECT 102.455 140.775 103.145 141.335 ;
        RECT 103.315 140.605 103.525 141.505 ;
        RECT 102.570 140.385 103.525 140.605 ;
        RECT 103.695 141.335 104.095 142.135 ;
        RECT 104.285 141.675 104.565 142.135 ;
        RECT 105.085 141.845 105.410 142.305 ;
        RECT 104.285 141.505 105.410 141.675 ;
        RECT 105.580 141.565 105.965 142.135 ;
        RECT 104.960 141.395 105.410 141.505 ;
        RECT 103.695 140.775 104.790 141.335 ;
        RECT 104.960 141.065 105.515 141.395 ;
        RECT 102.570 139.925 102.855 140.385 ;
        RECT 103.025 139.755 103.295 140.215 ;
        RECT 103.695 139.925 104.095 140.775 ;
        RECT 104.960 140.605 105.410 141.065 ;
        RECT 105.685 140.895 105.965 141.565 ;
        RECT 106.135 141.535 107.805 142.305 ;
        RECT 106.135 141.015 106.885 141.535 ;
        RECT 104.285 140.385 105.410 140.605 ;
        RECT 104.285 139.925 104.565 140.385 ;
        RECT 105.085 139.755 105.410 140.215 ;
        RECT 105.580 139.925 105.965 140.895 ;
        RECT 107.055 140.845 107.805 141.365 ;
        RECT 106.135 139.755 107.805 140.845 ;
        RECT 107.975 141.360 108.315 142.135 ;
        RECT 108.485 141.845 108.655 142.305 ;
        RECT 108.895 141.870 109.255 142.135 ;
        RECT 108.895 141.865 109.250 141.870 ;
        RECT 108.895 141.855 109.245 141.865 ;
        RECT 108.895 141.850 109.240 141.855 ;
        RECT 108.895 141.840 109.235 141.850 ;
        RECT 109.885 141.845 110.055 142.305 ;
        RECT 108.895 141.835 109.230 141.840 ;
        RECT 108.895 141.825 109.220 141.835 ;
        RECT 108.895 141.815 109.210 141.825 ;
        RECT 108.895 141.675 109.195 141.815 ;
        RECT 108.485 141.485 109.195 141.675 ;
        RECT 109.385 141.675 109.715 141.755 ;
        RECT 110.225 141.675 110.565 142.135 ;
        RECT 110.795 141.825 111.075 142.305 ;
        RECT 109.385 141.485 110.565 141.675 ;
        RECT 111.245 141.655 111.505 142.045 ;
        RECT 111.680 141.825 111.935 142.305 ;
        RECT 112.105 141.655 112.400 142.045 ;
        RECT 112.580 141.825 112.855 142.305 ;
        RECT 113.025 141.805 113.325 142.135 ;
        RECT 110.750 141.485 112.400 141.655 ;
        RECT 107.975 139.925 108.255 141.360 ;
        RECT 108.485 140.915 108.770 141.485 ;
        RECT 108.955 141.085 109.425 141.315 ;
        RECT 109.595 141.295 109.925 141.315 ;
        RECT 109.595 141.115 110.045 141.295 ;
        RECT 110.235 141.115 110.565 141.315 ;
        RECT 108.485 140.700 109.635 140.915 ;
        RECT 108.425 139.755 109.135 140.530 ;
        RECT 109.305 139.925 109.635 140.700 ;
        RECT 109.830 140.000 110.045 141.115 ;
        RECT 110.335 140.775 110.565 141.115 ;
        RECT 110.750 140.975 111.155 141.485 ;
        RECT 111.325 141.145 112.465 141.315 ;
        RECT 110.750 140.805 111.505 140.975 ;
        RECT 110.225 139.755 110.555 140.475 ;
        RECT 110.790 139.755 111.075 140.625 ;
        RECT 111.245 140.555 111.505 140.805 ;
        RECT 112.295 140.895 112.465 141.145 ;
        RECT 112.635 141.065 112.985 141.635 ;
        RECT 113.155 140.895 113.325 141.805 ;
        RECT 113.495 141.535 117.005 142.305 ;
        RECT 117.635 141.675 117.975 142.135 ;
        RECT 118.145 141.845 118.315 142.305 ;
        RECT 118.945 141.870 119.305 142.135 ;
        RECT 118.950 141.865 119.305 141.870 ;
        RECT 118.955 141.855 119.305 141.865 ;
        RECT 118.960 141.850 119.305 141.855 ;
        RECT 118.965 141.840 119.305 141.850 ;
        RECT 119.545 141.845 119.715 142.305 ;
        RECT 118.970 141.835 119.305 141.840 ;
        RECT 118.980 141.825 119.305 141.835 ;
        RECT 118.990 141.815 119.305 141.825 ;
        RECT 118.485 141.675 118.815 141.755 ;
        RECT 113.495 141.015 115.145 141.535 ;
        RECT 117.635 141.485 118.815 141.675 ;
        RECT 119.005 141.675 119.305 141.815 ;
        RECT 119.005 141.485 119.715 141.675 ;
        RECT 112.295 140.725 113.325 140.895 ;
        RECT 115.315 140.845 117.005 141.365 ;
        RECT 111.245 140.385 112.365 140.555 ;
        RECT 111.245 139.925 111.505 140.385 ;
        RECT 111.680 139.755 111.935 140.215 ;
        RECT 112.105 139.925 112.365 140.385 ;
        RECT 112.535 139.755 112.845 140.555 ;
        RECT 113.015 139.925 113.325 140.725 ;
        RECT 113.495 139.755 117.005 140.845 ;
        RECT 117.635 141.115 117.965 141.315 ;
        RECT 118.275 141.295 118.605 141.315 ;
        RECT 118.155 141.115 118.605 141.295 ;
        RECT 117.635 140.775 117.865 141.115 ;
        RECT 117.645 139.755 117.975 140.475 ;
        RECT 118.155 140.000 118.370 141.115 ;
        RECT 118.775 141.085 119.245 141.315 ;
        RECT 119.430 140.915 119.715 141.485 ;
        RECT 119.885 141.360 120.225 142.135 ;
        RECT 120.395 141.580 120.685 142.305 ;
        RECT 120.905 141.650 121.235 142.085 ;
        RECT 121.405 141.695 121.575 142.305 ;
        RECT 118.565 140.700 119.715 140.915 ;
        RECT 118.565 139.925 118.895 140.700 ;
        RECT 119.065 139.755 119.775 140.530 ;
        RECT 119.945 139.925 120.225 141.360 ;
        RECT 120.855 141.565 121.235 141.650 ;
        RECT 121.745 141.565 122.075 142.090 ;
        RECT 122.335 141.775 122.545 142.305 ;
        RECT 122.820 141.855 123.605 142.025 ;
        RECT 123.775 141.855 124.180 142.025 ;
        RECT 120.855 141.525 121.080 141.565 ;
        RECT 120.855 140.945 121.025 141.525 ;
        RECT 121.745 141.395 121.945 141.565 ;
        RECT 122.820 141.395 122.990 141.855 ;
        RECT 121.195 141.065 121.945 141.395 ;
        RECT 122.115 141.065 122.990 141.395 ;
        RECT 120.395 139.755 120.685 140.920 ;
        RECT 120.855 140.895 121.070 140.945 ;
        RECT 120.855 140.815 121.245 140.895 ;
        RECT 120.915 139.970 121.245 140.815 ;
        RECT 121.755 140.860 121.945 141.065 ;
        RECT 121.415 139.755 121.585 140.765 ;
        RECT 121.755 140.485 122.650 140.860 ;
        RECT 121.755 139.925 122.095 140.485 ;
        RECT 122.325 139.755 122.640 140.255 ;
        RECT 122.820 140.225 122.990 141.065 ;
        RECT 123.160 141.355 123.625 141.685 ;
        RECT 124.010 141.625 124.180 141.855 ;
        RECT 124.360 141.805 124.730 142.305 ;
        RECT 125.050 141.855 125.725 142.025 ;
        RECT 125.920 141.855 126.255 142.025 ;
        RECT 123.160 140.395 123.480 141.355 ;
        RECT 124.010 141.325 124.840 141.625 ;
        RECT 123.650 140.425 123.840 141.145 ;
        RECT 124.010 140.255 124.180 141.325 ;
        RECT 124.640 141.295 124.840 141.325 ;
        RECT 124.350 141.075 124.520 141.145 ;
        RECT 125.050 141.075 125.220 141.855 ;
        RECT 126.085 141.715 126.255 141.855 ;
        RECT 126.425 141.845 126.675 142.305 ;
        RECT 124.350 140.905 125.220 141.075 ;
        RECT 125.390 141.435 125.915 141.655 ;
        RECT 126.085 141.585 126.310 141.715 ;
        RECT 124.350 140.815 124.860 140.905 ;
        RECT 122.820 140.055 123.705 140.225 ;
        RECT 123.930 139.925 124.180 140.255 ;
        RECT 124.350 139.755 124.520 140.555 ;
        RECT 124.690 140.200 124.860 140.815 ;
        RECT 125.390 140.735 125.560 141.435 ;
        RECT 125.030 140.370 125.560 140.735 ;
        RECT 125.730 140.670 125.970 141.265 ;
        RECT 126.140 140.480 126.310 141.585 ;
        RECT 126.480 140.725 126.760 141.675 ;
        RECT 126.005 140.350 126.310 140.480 ;
        RECT 124.690 140.030 125.795 140.200 ;
        RECT 126.005 139.925 126.255 140.350 ;
        RECT 126.425 139.755 126.690 140.215 ;
        RECT 126.930 139.925 127.115 142.045 ;
        RECT 127.285 141.925 127.615 142.305 ;
        RECT 127.785 141.755 127.955 142.045 ;
        RECT 127.290 141.585 127.955 141.755 ;
        RECT 127.290 140.595 127.520 141.585 ;
        RECT 127.690 140.765 128.040 141.415 ;
        RECT 128.215 141.360 128.555 142.135 ;
        RECT 128.725 141.845 128.895 142.305 ;
        RECT 129.135 141.870 129.495 142.135 ;
        RECT 129.135 141.865 129.490 141.870 ;
        RECT 129.135 141.855 129.485 141.865 ;
        RECT 129.135 141.850 129.480 141.855 ;
        RECT 129.135 141.840 129.475 141.850 ;
        RECT 130.125 141.845 130.295 142.305 ;
        RECT 129.135 141.835 129.470 141.840 ;
        RECT 129.135 141.825 129.460 141.835 ;
        RECT 129.135 141.815 129.450 141.825 ;
        RECT 129.135 141.675 129.435 141.815 ;
        RECT 128.725 141.485 129.435 141.675 ;
        RECT 129.625 141.675 129.955 141.755 ;
        RECT 130.465 141.675 130.805 142.135 ;
        RECT 129.625 141.485 130.805 141.675 ;
        RECT 130.975 141.535 133.565 142.305 ;
        RECT 133.740 141.565 133.995 142.135 ;
        RECT 134.165 141.905 134.495 142.305 ;
        RECT 134.920 141.770 135.450 142.135 ;
        RECT 135.640 141.965 135.915 142.135 ;
        RECT 135.635 141.795 135.915 141.965 ;
        RECT 134.920 141.735 135.095 141.770 ;
        RECT 134.165 141.565 135.095 141.735 ;
        RECT 127.290 140.425 127.955 140.595 ;
        RECT 127.285 139.755 127.615 140.255 ;
        RECT 127.785 139.925 127.955 140.425 ;
        RECT 128.215 139.925 128.495 141.360 ;
        RECT 128.725 140.915 129.010 141.485 ;
        RECT 129.195 141.085 129.665 141.315 ;
        RECT 129.835 141.295 130.165 141.315 ;
        RECT 129.835 141.115 130.285 141.295 ;
        RECT 130.475 141.115 130.805 141.315 ;
        RECT 128.725 140.700 129.875 140.915 ;
        RECT 128.665 139.755 129.375 140.530 ;
        RECT 129.545 139.925 129.875 140.700 ;
        RECT 130.070 140.000 130.285 141.115 ;
        RECT 130.575 140.775 130.805 141.115 ;
        RECT 130.975 141.015 132.185 141.535 ;
        RECT 132.355 140.845 133.565 141.365 ;
        RECT 130.465 139.755 130.795 140.475 ;
        RECT 130.975 139.755 133.565 140.845 ;
        RECT 133.740 140.895 133.910 141.565 ;
        RECT 134.165 141.395 134.335 141.565 ;
        RECT 134.080 141.065 134.335 141.395 ;
        RECT 134.560 141.065 134.755 141.395 ;
        RECT 133.740 139.925 134.075 140.895 ;
        RECT 134.245 139.755 134.415 140.895 ;
        RECT 134.585 140.095 134.755 141.065 ;
        RECT 134.925 140.435 135.095 141.565 ;
        RECT 135.265 140.775 135.435 141.575 ;
        RECT 135.640 140.975 135.915 141.795 ;
        RECT 136.085 140.775 136.275 142.135 ;
        RECT 136.455 141.770 136.965 142.305 ;
        RECT 137.185 141.495 137.430 142.100 ;
        RECT 137.880 141.565 138.135 142.135 ;
        RECT 138.305 141.905 138.635 142.305 ;
        RECT 139.060 141.770 139.590 142.135 ;
        RECT 139.060 141.735 139.235 141.770 ;
        RECT 138.305 141.565 139.235 141.735 ;
        RECT 139.780 141.625 140.055 142.135 ;
        RECT 136.475 141.325 137.705 141.495 ;
        RECT 135.265 140.605 136.275 140.775 ;
        RECT 136.445 140.760 137.195 140.950 ;
        RECT 134.925 140.265 136.050 140.435 ;
        RECT 136.445 140.095 136.615 140.760 ;
        RECT 137.365 140.515 137.705 141.325 ;
        RECT 134.585 139.925 136.615 140.095 ;
        RECT 136.785 139.755 136.955 140.515 ;
        RECT 137.190 140.105 137.705 140.515 ;
        RECT 137.880 140.895 138.050 141.565 ;
        RECT 138.305 141.395 138.475 141.565 ;
        RECT 138.220 141.065 138.475 141.395 ;
        RECT 138.700 141.065 138.895 141.395 ;
        RECT 137.880 139.925 138.215 140.895 ;
        RECT 138.385 139.755 138.555 140.895 ;
        RECT 138.725 140.095 138.895 141.065 ;
        RECT 139.065 140.435 139.235 141.565 ;
        RECT 139.405 140.775 139.575 141.575 ;
        RECT 139.775 141.455 140.055 141.625 ;
        RECT 139.780 140.975 140.055 141.455 ;
        RECT 140.225 140.775 140.415 142.135 ;
        RECT 140.595 141.770 141.105 142.305 ;
        RECT 141.325 141.495 141.570 142.100 ;
        RECT 142.105 141.755 142.275 142.135 ;
        RECT 142.455 141.925 142.785 142.305 ;
        RECT 142.105 141.585 142.770 141.755 ;
        RECT 142.965 141.630 143.225 142.135 ;
        RECT 140.615 141.325 141.845 141.495 ;
        RECT 139.405 140.605 140.415 140.775 ;
        RECT 140.585 140.760 141.335 140.950 ;
        RECT 139.065 140.265 140.190 140.435 ;
        RECT 140.585 140.095 140.755 140.760 ;
        RECT 141.505 140.515 141.845 141.325 ;
        RECT 142.035 141.035 142.365 141.405 ;
        RECT 142.600 141.330 142.770 141.585 ;
        RECT 142.600 141.000 142.885 141.330 ;
        RECT 142.600 140.855 142.770 141.000 ;
        RECT 138.725 139.925 140.755 140.095 ;
        RECT 140.925 139.755 141.095 140.515 ;
        RECT 141.330 140.105 141.845 140.515 ;
        RECT 142.105 140.685 142.770 140.855 ;
        RECT 143.055 140.830 143.225 141.630 ;
        RECT 143.945 141.755 144.115 142.135 ;
        RECT 144.330 141.925 144.660 142.305 ;
        RECT 143.945 141.585 144.660 141.755 ;
        RECT 143.855 141.035 144.210 141.405 ;
        RECT 144.490 141.395 144.660 141.585 ;
        RECT 144.830 141.560 145.085 142.135 ;
        RECT 144.490 141.065 144.745 141.395 ;
        RECT 144.490 140.855 144.660 141.065 ;
        RECT 142.105 139.925 142.275 140.685 ;
        RECT 142.455 139.755 142.785 140.515 ;
        RECT 142.955 139.925 143.225 140.830 ;
        RECT 143.945 140.685 144.660 140.855 ;
        RECT 144.915 140.830 145.085 141.560 ;
        RECT 145.260 141.465 145.520 142.305 ;
        RECT 145.695 141.555 146.905 142.305 ;
        RECT 143.945 139.925 144.115 140.685 ;
        RECT 144.330 139.755 144.660 140.515 ;
        RECT 144.830 139.925 145.085 140.830 ;
        RECT 145.260 139.755 145.520 140.905 ;
        RECT 145.695 140.845 146.215 141.385 ;
        RECT 146.385 141.015 146.905 141.555 ;
        RECT 145.695 139.755 146.905 140.845 ;
        RECT 17.270 139.585 146.990 139.755 ;
        RECT 17.355 138.495 18.565 139.585 ;
        RECT 17.355 137.785 17.875 138.325 ;
        RECT 18.045 137.955 18.565 138.495 ;
        RECT 18.740 138.445 19.075 139.415 ;
        RECT 19.245 138.445 19.415 139.585 ;
        RECT 19.585 139.245 21.615 139.415 ;
        RECT 17.355 137.035 18.565 137.785 ;
        RECT 18.740 137.775 18.910 138.445 ;
        RECT 19.585 138.275 19.755 139.245 ;
        RECT 19.080 137.945 19.335 138.275 ;
        RECT 19.560 137.945 19.755 138.275 ;
        RECT 19.925 138.905 21.050 139.075 ;
        RECT 19.165 137.775 19.335 137.945 ;
        RECT 19.925 137.775 20.095 138.905 ;
        RECT 18.740 137.205 18.995 137.775 ;
        RECT 19.165 137.605 20.095 137.775 ;
        RECT 20.265 138.565 21.275 138.735 ;
        RECT 20.265 137.765 20.435 138.565 ;
        RECT 20.640 138.225 20.915 138.365 ;
        RECT 20.635 138.055 20.915 138.225 ;
        RECT 19.920 137.570 20.095 137.605 ;
        RECT 19.165 137.035 19.495 137.435 ;
        RECT 19.920 137.205 20.450 137.570 ;
        RECT 20.640 137.205 20.915 138.055 ;
        RECT 21.085 137.205 21.275 138.565 ;
        RECT 21.445 138.580 21.615 139.245 ;
        RECT 21.785 138.825 21.955 139.585 ;
        RECT 22.190 138.825 22.705 139.235 ;
        RECT 21.445 138.390 22.195 138.580 ;
        RECT 22.365 138.015 22.705 138.825 ;
        RECT 22.935 138.525 23.265 139.370 ;
        RECT 23.435 138.575 23.605 139.585 ;
        RECT 23.775 138.855 24.115 139.415 ;
        RECT 24.345 139.085 24.660 139.585 ;
        RECT 24.840 139.115 25.725 139.285 ;
        RECT 21.475 137.845 22.705 138.015 ;
        RECT 22.875 138.445 23.265 138.525 ;
        RECT 23.775 138.480 24.670 138.855 ;
        RECT 22.875 138.395 23.090 138.445 ;
        RECT 21.455 137.035 21.965 137.570 ;
        RECT 22.185 137.240 22.430 137.845 ;
        RECT 22.875 137.815 23.045 138.395 ;
        RECT 23.775 138.275 23.965 138.480 ;
        RECT 24.840 138.275 25.010 139.115 ;
        RECT 25.950 139.085 26.200 139.415 ;
        RECT 23.215 137.945 23.965 138.275 ;
        RECT 24.135 137.945 25.010 138.275 ;
        RECT 22.875 137.775 23.100 137.815 ;
        RECT 23.765 137.775 23.965 137.945 ;
        RECT 22.875 137.690 23.255 137.775 ;
        RECT 22.925 137.255 23.255 137.690 ;
        RECT 23.425 137.035 23.595 137.645 ;
        RECT 23.765 137.250 24.095 137.775 ;
        RECT 24.355 137.035 24.565 137.565 ;
        RECT 24.840 137.485 25.010 137.945 ;
        RECT 25.180 137.985 25.500 138.945 ;
        RECT 25.670 138.195 25.860 138.915 ;
        RECT 26.030 138.015 26.200 139.085 ;
        RECT 26.370 138.785 26.540 139.585 ;
        RECT 26.710 139.140 27.815 139.310 ;
        RECT 26.710 138.525 26.880 139.140 ;
        RECT 28.025 138.990 28.275 139.415 ;
        RECT 28.445 139.125 28.710 139.585 ;
        RECT 27.050 138.605 27.580 138.970 ;
        RECT 28.025 138.860 28.330 138.990 ;
        RECT 26.370 138.435 26.880 138.525 ;
        RECT 26.370 138.265 27.240 138.435 ;
        RECT 26.370 138.195 26.540 138.265 ;
        RECT 26.660 138.015 26.860 138.045 ;
        RECT 25.180 137.655 25.645 137.985 ;
        RECT 26.030 137.715 26.860 138.015 ;
        RECT 26.030 137.485 26.200 137.715 ;
        RECT 24.840 137.315 25.625 137.485 ;
        RECT 25.795 137.315 26.200 137.485 ;
        RECT 26.380 137.035 26.750 137.535 ;
        RECT 27.070 137.485 27.240 138.265 ;
        RECT 27.410 137.905 27.580 138.605 ;
        RECT 27.750 138.075 27.990 138.670 ;
        RECT 27.410 137.685 27.935 137.905 ;
        RECT 28.160 137.755 28.330 138.860 ;
        RECT 28.105 137.625 28.330 137.755 ;
        RECT 28.500 137.665 28.780 138.615 ;
        RECT 28.105 137.485 28.275 137.625 ;
        RECT 27.070 137.315 27.745 137.485 ;
        RECT 27.940 137.315 28.275 137.485 ;
        RECT 28.445 137.035 28.695 137.495 ;
        RECT 28.950 137.295 29.135 139.415 ;
        RECT 29.305 139.085 29.635 139.585 ;
        RECT 29.805 138.915 29.975 139.415 ;
        RECT 29.310 138.745 29.975 138.915 ;
        RECT 29.310 137.755 29.540 138.745 ;
        RECT 29.710 137.925 30.060 138.575 ;
        RECT 30.235 138.420 30.525 139.585 ;
        RECT 30.695 138.785 31.135 139.415 ;
        RECT 30.695 137.775 31.005 138.785 ;
        RECT 31.310 138.735 31.625 139.585 ;
        RECT 31.795 139.245 33.225 139.415 ;
        RECT 31.795 138.565 31.965 139.245 ;
        RECT 31.175 138.395 31.965 138.565 ;
        RECT 31.175 137.945 31.345 138.395 ;
        RECT 32.135 138.275 32.335 139.075 ;
        RECT 31.515 137.945 31.905 138.225 ;
        RECT 32.090 137.945 32.335 138.275 ;
        RECT 32.535 137.945 32.785 139.075 ;
        RECT 32.975 138.615 33.225 139.245 ;
        RECT 33.405 138.785 33.735 139.585 ;
        RECT 33.915 139.150 39.260 139.585 ;
        RECT 39.435 139.150 44.780 139.585 ;
        RECT 44.955 139.150 50.300 139.585 ;
        RECT 50.475 139.150 55.820 139.585 ;
        RECT 32.975 138.445 33.745 138.615 ;
        RECT 33.000 137.945 33.405 138.275 ;
        RECT 33.575 137.775 33.745 138.445 ;
        RECT 29.310 137.585 29.975 137.755 ;
        RECT 29.305 137.035 29.635 137.415 ;
        RECT 29.805 137.295 29.975 137.585 ;
        RECT 30.235 137.035 30.525 137.760 ;
        RECT 30.695 137.215 31.135 137.775 ;
        RECT 31.305 137.035 31.755 137.775 ;
        RECT 31.925 137.605 33.085 137.775 ;
        RECT 31.925 137.205 32.095 137.605 ;
        RECT 32.265 137.035 32.685 137.435 ;
        RECT 32.855 137.205 33.085 137.605 ;
        RECT 33.255 137.205 33.745 137.775 ;
        RECT 35.500 137.580 35.840 138.410 ;
        RECT 37.320 137.900 37.670 139.150 ;
        RECT 41.020 137.580 41.360 138.410 ;
        RECT 42.840 137.900 43.190 139.150 ;
        RECT 46.540 137.580 46.880 138.410 ;
        RECT 48.360 137.900 48.710 139.150 ;
        RECT 52.060 137.580 52.400 138.410 ;
        RECT 53.880 137.900 54.230 139.150 ;
        RECT 55.995 138.420 56.285 139.585 ;
        RECT 56.455 139.150 61.800 139.585 ;
        RECT 61.975 139.150 67.320 139.585 ;
        RECT 33.915 137.035 39.260 137.580 ;
        RECT 39.435 137.035 44.780 137.580 ;
        RECT 44.955 137.035 50.300 137.580 ;
        RECT 50.475 137.035 55.820 137.580 ;
        RECT 55.995 137.035 56.285 137.760 ;
        RECT 58.040 137.580 58.380 138.410 ;
        RECT 59.860 137.900 60.210 139.150 ;
        RECT 63.560 137.580 63.900 138.410 ;
        RECT 65.380 137.900 65.730 139.150 ;
        RECT 67.495 138.495 68.705 139.585 ;
        RECT 67.495 137.785 68.015 138.325 ;
        RECT 68.185 137.955 68.705 138.495 ;
        RECT 68.875 138.735 69.255 139.415 ;
        RECT 69.845 138.735 70.015 139.585 ;
        RECT 70.185 138.905 70.515 139.415 ;
        RECT 70.685 139.075 70.855 139.585 ;
        RECT 71.025 138.905 71.425 139.415 ;
        RECT 70.185 138.735 71.425 138.905 ;
        RECT 56.455 137.035 61.800 137.580 ;
        RECT 61.975 137.035 67.320 137.580 ;
        RECT 67.495 137.035 68.705 137.785 ;
        RECT 68.875 137.775 69.045 138.735 ;
        RECT 69.215 138.395 70.520 138.565 ;
        RECT 71.605 138.485 71.925 139.415 ;
        RECT 69.215 137.945 69.460 138.395 ;
        RECT 69.630 138.025 70.180 138.225 ;
        RECT 70.350 138.195 70.520 138.395 ;
        RECT 71.295 138.315 71.925 138.485 ;
        RECT 72.095 138.715 72.370 139.415 ;
        RECT 72.580 139.040 72.795 139.585 ;
        RECT 72.965 139.075 73.440 139.415 ;
        RECT 73.610 139.080 74.225 139.585 ;
        RECT 73.610 138.905 73.805 139.080 ;
        RECT 70.350 138.025 70.725 138.195 ;
        RECT 70.895 137.775 71.125 138.275 ;
        RECT 68.875 137.605 71.125 137.775 ;
        RECT 68.925 137.035 69.255 137.425 ;
        RECT 69.425 137.285 69.595 137.605 ;
        RECT 71.295 137.435 71.465 138.315 ;
        RECT 69.765 137.035 70.095 137.425 ;
        RECT 70.510 137.265 71.465 137.435 ;
        RECT 71.635 137.035 71.925 137.870 ;
        RECT 72.095 137.685 72.265 138.715 ;
        RECT 72.540 138.545 73.255 138.840 ;
        RECT 73.475 138.715 73.805 138.905 ;
        RECT 73.975 138.545 74.225 138.910 ;
        RECT 72.435 138.375 74.225 138.545 ;
        RECT 72.435 137.945 72.665 138.375 ;
        RECT 72.095 137.205 72.355 137.685 ;
        RECT 72.835 137.675 73.245 138.195 ;
        RECT 72.525 137.035 72.855 137.495 ;
        RECT 73.045 137.255 73.245 137.675 ;
        RECT 73.415 137.520 73.670 138.375 ;
        RECT 74.465 138.195 74.635 139.415 ;
        RECT 74.885 139.075 75.145 139.585 ;
        RECT 75.315 139.150 80.660 139.585 ;
        RECT 73.840 137.945 74.635 138.195 ;
        RECT 74.805 138.025 75.145 138.905 ;
        RECT 74.385 137.855 74.635 137.945 ;
        RECT 73.415 137.255 74.205 137.520 ;
        RECT 74.385 137.435 74.715 137.855 ;
        RECT 74.885 137.035 75.145 137.855 ;
        RECT 76.900 137.580 77.240 138.410 ;
        RECT 78.720 137.900 79.070 139.150 ;
        RECT 81.755 138.420 82.045 139.585 ;
        RECT 82.675 139.075 83.865 139.365 ;
        RECT 82.695 138.735 83.865 138.905 ;
        RECT 84.035 138.785 84.315 139.585 ;
        RECT 82.695 138.445 83.020 138.735 ;
        RECT 83.695 138.615 83.865 138.735 ;
        RECT 83.190 138.275 83.385 138.565 ;
        RECT 83.695 138.445 84.355 138.615 ;
        RECT 84.525 138.445 84.800 139.415 ;
        RECT 84.975 138.445 85.235 139.585 ;
        RECT 85.475 139.075 87.090 139.405 ;
        RECT 84.185 138.275 84.355 138.445 ;
        RECT 82.675 137.945 83.020 138.275 ;
        RECT 83.190 137.945 84.015 138.275 ;
        RECT 84.185 137.945 84.460 138.275 ;
        RECT 84.185 137.775 84.355 137.945 ;
        RECT 75.315 137.035 80.660 137.580 ;
        RECT 81.755 137.035 82.045 137.760 ;
        RECT 82.690 137.605 84.355 137.775 ;
        RECT 84.630 137.710 84.800 138.445 ;
        RECT 85.485 138.275 85.655 138.835 ;
        RECT 85.915 138.735 87.090 138.905 ;
        RECT 87.260 138.785 87.540 139.585 ;
        RECT 85.915 138.445 86.245 138.735 ;
        RECT 86.920 138.615 87.090 138.735 ;
        RECT 86.415 138.275 86.660 138.565 ;
        RECT 86.920 138.445 87.580 138.615 ;
        RECT 87.750 138.445 88.025 139.415 ;
        RECT 87.410 138.275 87.580 138.445 ;
        RECT 84.980 138.025 85.315 138.275 ;
        RECT 85.485 137.945 86.200 138.275 ;
        RECT 86.415 137.945 87.240 138.275 ;
        RECT 87.410 137.945 87.685 138.275 ;
        RECT 85.485 137.855 85.735 137.945 ;
        RECT 82.690 137.255 82.945 137.605 ;
        RECT 83.115 137.035 83.445 137.435 ;
        RECT 83.615 137.255 83.785 137.605 ;
        RECT 83.955 137.035 84.335 137.435 ;
        RECT 84.525 137.365 84.800 137.710 ;
        RECT 84.975 137.035 85.235 137.855 ;
        RECT 85.405 137.435 85.735 137.855 ;
        RECT 87.410 137.775 87.580 137.945 ;
        RECT 85.915 137.605 87.580 137.775 ;
        RECT 87.855 137.710 88.025 138.445 ;
        RECT 85.915 137.205 86.175 137.605 ;
        RECT 86.345 137.035 86.675 137.435 ;
        RECT 86.845 137.255 87.015 137.605 ;
        RECT 87.185 137.035 87.560 137.435 ;
        RECT 87.750 137.365 88.025 137.710 ;
        RECT 88.200 138.445 88.535 139.415 ;
        RECT 88.705 138.445 88.875 139.585 ;
        RECT 89.045 139.245 91.075 139.415 ;
        RECT 88.200 137.775 88.370 138.445 ;
        RECT 89.045 138.275 89.215 139.245 ;
        RECT 88.540 137.945 88.795 138.275 ;
        RECT 89.020 137.945 89.215 138.275 ;
        RECT 89.385 138.905 90.510 139.075 ;
        RECT 88.625 137.775 88.795 137.945 ;
        RECT 89.385 137.775 89.555 138.905 ;
        RECT 88.200 137.205 88.455 137.775 ;
        RECT 88.625 137.605 89.555 137.775 ;
        RECT 89.725 138.565 90.735 138.735 ;
        RECT 89.725 137.765 89.895 138.565 ;
        RECT 90.100 138.225 90.375 138.365 ;
        RECT 90.095 138.055 90.375 138.225 ;
        RECT 89.380 137.570 89.555 137.605 ;
        RECT 88.625 137.035 88.955 137.435 ;
        RECT 89.380 137.205 89.910 137.570 ;
        RECT 90.100 137.205 90.375 138.055 ;
        RECT 90.545 137.205 90.735 138.565 ;
        RECT 90.905 138.580 91.075 139.245 ;
        RECT 91.245 138.825 91.415 139.585 ;
        RECT 91.650 138.825 92.165 139.235 ;
        RECT 90.905 138.390 91.655 138.580 ;
        RECT 91.825 138.015 92.165 138.825 ;
        RECT 90.935 137.845 92.165 138.015 ;
        RECT 92.340 138.445 92.675 139.415 ;
        RECT 92.845 138.445 93.015 139.585 ;
        RECT 93.185 139.245 95.215 139.415 ;
        RECT 90.915 137.035 91.425 137.570 ;
        RECT 91.645 137.240 91.890 137.845 ;
        RECT 92.340 137.775 92.510 138.445 ;
        RECT 93.185 138.275 93.355 139.245 ;
        RECT 92.680 137.945 92.935 138.275 ;
        RECT 93.160 137.945 93.355 138.275 ;
        RECT 93.525 138.905 94.650 139.075 ;
        RECT 92.765 137.775 92.935 137.945 ;
        RECT 93.525 137.775 93.695 138.905 ;
        RECT 92.340 137.205 92.595 137.775 ;
        RECT 92.765 137.605 93.695 137.775 ;
        RECT 93.865 138.565 94.875 138.735 ;
        RECT 93.865 137.765 94.035 138.565 ;
        RECT 94.240 137.885 94.515 138.365 ;
        RECT 94.235 137.715 94.515 137.885 ;
        RECT 93.520 137.570 93.695 137.605 ;
        RECT 92.765 137.035 93.095 137.435 ;
        RECT 93.520 137.205 94.050 137.570 ;
        RECT 94.240 137.205 94.515 137.715 ;
        RECT 94.685 137.205 94.875 138.565 ;
        RECT 95.045 138.580 95.215 139.245 ;
        RECT 95.385 138.825 95.555 139.585 ;
        RECT 95.790 138.825 96.305 139.235 ;
        RECT 95.045 138.390 95.795 138.580 ;
        RECT 95.965 138.015 96.305 138.825 ;
        RECT 96.475 138.495 99.985 139.585 ;
        RECT 95.075 137.845 96.305 138.015 ;
        RECT 95.055 137.035 95.565 137.570 ;
        RECT 95.785 137.240 96.030 137.845 ;
        RECT 96.475 137.805 98.125 138.325 ;
        RECT 98.295 137.975 99.985 138.495 ;
        RECT 100.620 138.445 100.875 139.585 ;
        RECT 101.045 138.615 101.375 139.415 ;
        RECT 101.545 138.785 101.715 139.585 ;
        RECT 101.885 138.615 102.215 139.415 ;
        RECT 102.385 138.785 102.555 139.585 ;
        RECT 102.725 138.615 103.055 139.415 ;
        RECT 103.225 138.785 103.395 139.585 ;
        RECT 103.565 138.615 103.895 139.415 ;
        RECT 104.065 138.785 104.315 139.585 ;
        RECT 101.045 138.445 103.895 138.615 ;
        RECT 100.640 138.025 102.260 138.275 ;
        RECT 102.440 138.025 102.975 138.445 ;
        RECT 103.145 138.025 104.585 138.275 ;
        RECT 96.475 137.035 99.985 137.805 ;
        RECT 100.620 137.665 102.555 137.855 ;
        RECT 100.620 137.205 100.955 137.665 ;
        RECT 101.125 137.035 101.295 137.495 ;
        RECT 101.465 137.205 101.795 137.665 ;
        RECT 101.965 137.035 102.135 137.495 ;
        RECT 102.305 137.415 102.555 137.665 ;
        RECT 102.725 137.755 102.975 138.025 ;
        RECT 104.755 137.980 105.035 139.415 ;
        RECT 105.205 138.810 105.915 139.585 ;
        RECT 106.085 138.640 106.415 139.415 ;
        RECT 105.265 138.425 106.415 138.640 ;
        RECT 102.725 137.585 103.895 137.755 ;
        RECT 104.065 137.415 104.315 137.835 ;
        RECT 102.305 137.205 104.315 137.415 ;
        RECT 104.755 137.205 105.095 137.980 ;
        RECT 105.265 137.855 105.550 138.425 ;
        RECT 105.735 138.025 106.205 138.255 ;
        RECT 106.610 138.225 106.825 139.340 ;
        RECT 107.005 138.865 107.335 139.585 ;
        RECT 107.115 138.225 107.345 138.565 ;
        RECT 107.515 138.420 107.805 139.585 ;
        RECT 107.975 138.495 109.645 139.585 ;
        RECT 106.375 138.045 106.825 138.225 ;
        RECT 106.375 138.025 106.705 138.045 ;
        RECT 107.015 138.025 107.345 138.225 ;
        RECT 105.265 137.665 105.975 137.855 ;
        RECT 105.675 137.525 105.975 137.665 ;
        RECT 106.165 137.665 107.345 137.855 ;
        RECT 107.975 137.805 108.725 138.325 ;
        RECT 108.895 137.975 109.645 138.495 ;
        RECT 110.275 138.445 110.660 139.415 ;
        RECT 110.830 139.125 111.155 139.585 ;
        RECT 111.675 138.955 111.955 139.415 ;
        RECT 110.830 138.735 111.955 138.955 ;
        RECT 106.165 137.585 106.495 137.665 ;
        RECT 105.675 137.515 105.990 137.525 ;
        RECT 105.675 137.505 106.000 137.515 ;
        RECT 105.675 137.500 106.010 137.505 ;
        RECT 105.265 137.035 105.435 137.495 ;
        RECT 105.675 137.490 106.015 137.500 ;
        RECT 105.675 137.485 106.020 137.490 ;
        RECT 105.675 137.475 106.025 137.485 ;
        RECT 105.675 137.470 106.030 137.475 ;
        RECT 105.675 137.205 106.035 137.470 ;
        RECT 106.665 137.035 106.835 137.495 ;
        RECT 107.005 137.205 107.345 137.665 ;
        RECT 107.515 137.035 107.805 137.760 ;
        RECT 107.975 137.035 109.645 137.805 ;
        RECT 110.275 137.775 110.555 138.445 ;
        RECT 110.830 138.275 111.280 138.735 ;
        RECT 112.145 138.565 112.545 139.415 ;
        RECT 112.945 139.125 113.215 139.585 ;
        RECT 113.385 138.955 113.670 139.415 ;
        RECT 110.725 137.945 111.280 138.275 ;
        RECT 111.450 138.005 112.545 138.565 ;
        RECT 110.830 137.835 111.280 137.945 ;
        RECT 110.275 137.205 110.660 137.775 ;
        RECT 110.830 137.665 111.955 137.835 ;
        RECT 110.830 137.035 111.155 137.495 ;
        RECT 111.675 137.205 111.955 137.665 ;
        RECT 112.145 137.205 112.545 138.005 ;
        RECT 112.715 138.735 113.670 138.955 ;
        RECT 114.045 138.915 114.215 139.415 ;
        RECT 114.385 139.085 114.715 139.585 ;
        RECT 114.045 138.745 114.710 138.915 ;
        RECT 112.715 137.835 112.925 138.735 ;
        RECT 113.095 138.005 113.785 138.565 ;
        RECT 113.960 137.925 114.310 138.575 ;
        RECT 112.715 137.665 113.670 137.835 ;
        RECT 114.480 137.755 114.710 138.745 ;
        RECT 112.945 137.035 113.215 137.495 ;
        RECT 113.385 137.205 113.670 137.665 ;
        RECT 114.045 137.585 114.710 137.755 ;
        RECT 114.045 137.295 114.215 137.585 ;
        RECT 114.385 137.035 114.715 137.415 ;
        RECT 114.885 137.295 115.070 139.415 ;
        RECT 115.310 139.125 115.575 139.585 ;
        RECT 115.745 138.990 115.995 139.415 ;
        RECT 116.205 139.140 117.310 139.310 ;
        RECT 115.690 138.860 115.995 138.990 ;
        RECT 115.240 137.665 115.520 138.615 ;
        RECT 115.690 137.755 115.860 138.860 ;
        RECT 116.030 138.075 116.270 138.670 ;
        RECT 116.440 138.605 116.970 138.970 ;
        RECT 116.440 137.905 116.610 138.605 ;
        RECT 117.140 138.525 117.310 139.140 ;
        RECT 117.480 138.785 117.650 139.585 ;
        RECT 117.820 139.085 118.070 139.415 ;
        RECT 118.295 139.115 119.180 139.285 ;
        RECT 117.140 138.435 117.650 138.525 ;
        RECT 115.690 137.625 115.915 137.755 ;
        RECT 116.085 137.685 116.610 137.905 ;
        RECT 116.780 138.265 117.650 138.435 ;
        RECT 115.325 137.035 115.575 137.495 ;
        RECT 115.745 137.485 115.915 137.625 ;
        RECT 116.780 137.485 116.950 138.265 ;
        RECT 117.480 138.195 117.650 138.265 ;
        RECT 117.160 138.015 117.360 138.045 ;
        RECT 117.820 138.015 117.990 139.085 ;
        RECT 118.160 138.195 118.350 138.915 ;
        RECT 117.160 137.715 117.990 138.015 ;
        RECT 118.520 137.985 118.840 138.945 ;
        RECT 115.745 137.315 116.080 137.485 ;
        RECT 116.275 137.315 116.950 137.485 ;
        RECT 117.270 137.035 117.640 137.535 ;
        RECT 117.820 137.485 117.990 137.715 ;
        RECT 118.375 137.655 118.840 137.985 ;
        RECT 119.010 138.275 119.180 139.115 ;
        RECT 119.360 139.085 119.675 139.585 ;
        RECT 119.905 138.855 120.245 139.415 ;
        RECT 119.350 138.480 120.245 138.855 ;
        RECT 120.415 138.575 120.585 139.585 ;
        RECT 120.055 138.275 120.245 138.480 ;
        RECT 120.755 138.525 121.085 139.370 ;
        RECT 121.405 138.915 121.575 139.415 ;
        RECT 121.745 139.085 122.075 139.585 ;
        RECT 121.405 138.745 122.070 138.915 ;
        RECT 120.755 138.445 121.145 138.525 ;
        RECT 120.930 138.395 121.145 138.445 ;
        RECT 119.010 137.945 119.885 138.275 ;
        RECT 120.055 137.945 120.805 138.275 ;
        RECT 119.010 137.485 119.180 137.945 ;
        RECT 120.055 137.775 120.255 137.945 ;
        RECT 120.975 137.815 121.145 138.395 ;
        RECT 121.320 137.925 121.670 138.575 ;
        RECT 120.920 137.775 121.145 137.815 ;
        RECT 117.820 137.315 118.225 137.485 ;
        RECT 118.395 137.315 119.180 137.485 ;
        RECT 119.455 137.035 119.665 137.565 ;
        RECT 119.925 137.250 120.255 137.775 ;
        RECT 120.765 137.690 121.145 137.775 ;
        RECT 121.840 137.755 122.070 138.745 ;
        RECT 120.425 137.035 120.595 137.645 ;
        RECT 120.765 137.255 121.095 137.690 ;
        RECT 121.405 137.585 122.070 137.755 ;
        RECT 121.405 137.295 121.575 137.585 ;
        RECT 121.745 137.035 122.075 137.415 ;
        RECT 122.245 137.295 122.430 139.415 ;
        RECT 122.670 139.125 122.935 139.585 ;
        RECT 123.105 138.990 123.355 139.415 ;
        RECT 123.565 139.140 124.670 139.310 ;
        RECT 123.050 138.860 123.355 138.990 ;
        RECT 122.600 137.665 122.880 138.615 ;
        RECT 123.050 137.755 123.220 138.860 ;
        RECT 123.390 138.075 123.630 138.670 ;
        RECT 123.800 138.605 124.330 138.970 ;
        RECT 123.800 137.905 123.970 138.605 ;
        RECT 124.500 138.525 124.670 139.140 ;
        RECT 124.840 138.785 125.010 139.585 ;
        RECT 125.180 139.085 125.430 139.415 ;
        RECT 125.655 139.115 126.540 139.285 ;
        RECT 124.500 138.435 125.010 138.525 ;
        RECT 123.050 137.625 123.275 137.755 ;
        RECT 123.445 137.685 123.970 137.905 ;
        RECT 124.140 138.265 125.010 138.435 ;
        RECT 122.685 137.035 122.935 137.495 ;
        RECT 123.105 137.485 123.275 137.625 ;
        RECT 124.140 137.485 124.310 138.265 ;
        RECT 124.840 138.195 125.010 138.265 ;
        RECT 124.520 138.015 124.720 138.045 ;
        RECT 125.180 138.015 125.350 139.085 ;
        RECT 125.520 138.195 125.710 138.915 ;
        RECT 124.520 137.715 125.350 138.015 ;
        RECT 125.880 137.985 126.200 138.945 ;
        RECT 123.105 137.315 123.440 137.485 ;
        RECT 123.635 137.315 124.310 137.485 ;
        RECT 124.630 137.035 125.000 137.535 ;
        RECT 125.180 137.485 125.350 137.715 ;
        RECT 125.735 137.655 126.200 137.985 ;
        RECT 126.370 138.275 126.540 139.115 ;
        RECT 126.720 139.085 127.035 139.585 ;
        RECT 127.265 138.855 127.605 139.415 ;
        RECT 126.710 138.480 127.605 138.855 ;
        RECT 127.775 138.575 127.945 139.585 ;
        RECT 127.415 138.275 127.605 138.480 ;
        RECT 128.115 138.525 128.445 139.370 ;
        RECT 128.115 138.445 128.505 138.525 ;
        RECT 128.675 138.495 130.345 139.585 ;
        RECT 130.605 138.965 130.775 139.395 ;
        RECT 130.945 139.135 131.275 139.585 ;
        RECT 130.605 138.735 131.280 138.965 ;
        RECT 128.290 138.395 128.505 138.445 ;
        RECT 126.370 137.945 127.245 138.275 ;
        RECT 127.415 137.945 128.165 138.275 ;
        RECT 126.370 137.485 126.540 137.945 ;
        RECT 127.415 137.775 127.615 137.945 ;
        RECT 128.335 137.815 128.505 138.395 ;
        RECT 128.280 137.775 128.505 137.815 ;
        RECT 125.180 137.315 125.585 137.485 ;
        RECT 125.755 137.315 126.540 137.485 ;
        RECT 126.815 137.035 127.025 137.565 ;
        RECT 127.285 137.250 127.615 137.775 ;
        RECT 128.125 137.690 128.505 137.775 ;
        RECT 128.675 137.805 129.425 138.325 ;
        RECT 129.595 137.975 130.345 138.495 ;
        RECT 127.785 137.035 127.955 137.645 ;
        RECT 128.125 137.255 128.455 137.690 ;
        RECT 128.675 137.035 130.345 137.805 ;
        RECT 130.575 137.715 130.875 138.565 ;
        RECT 131.045 138.085 131.280 138.735 ;
        RECT 131.450 138.425 131.735 139.370 ;
        RECT 131.915 139.115 132.600 139.585 ;
        RECT 131.910 138.595 132.605 138.905 ;
        RECT 132.780 138.530 133.085 139.315 ;
        RECT 131.450 138.275 132.310 138.425 ;
        RECT 131.450 138.255 132.735 138.275 ;
        RECT 131.045 137.755 131.580 138.085 ;
        RECT 131.750 137.895 132.735 138.255 ;
        RECT 131.045 137.605 131.265 137.755 ;
        RECT 130.520 137.035 130.855 137.540 ;
        RECT 131.025 137.230 131.265 137.605 ;
        RECT 131.750 137.560 131.920 137.895 ;
        RECT 132.910 137.725 133.085 138.530 ;
        RECT 133.275 138.420 133.565 139.585 ;
        RECT 133.740 138.635 134.005 139.405 ;
        RECT 134.175 138.865 134.505 139.585 ;
        RECT 134.695 139.045 134.955 139.405 ;
        RECT 135.125 139.215 135.455 139.585 ;
        RECT 135.625 139.045 135.885 139.405 ;
        RECT 134.695 138.815 135.885 139.045 ;
        RECT 136.455 138.635 136.745 139.405 ;
        RECT 137.505 138.915 137.675 139.415 ;
        RECT 137.845 139.085 138.175 139.585 ;
        RECT 137.505 138.745 138.170 138.915 ;
        RECT 131.545 137.365 131.920 137.560 ;
        RECT 131.545 137.220 131.715 137.365 ;
        RECT 132.280 137.035 132.675 137.530 ;
        RECT 132.845 137.205 133.085 137.725 ;
        RECT 133.275 137.035 133.565 137.760 ;
        RECT 133.740 137.215 134.075 138.635 ;
        RECT 134.250 138.455 136.745 138.635 ;
        RECT 134.250 137.765 134.475 138.455 ;
        RECT 134.675 137.945 134.955 138.275 ;
        RECT 135.135 137.945 135.710 138.275 ;
        RECT 135.890 137.945 136.325 138.275 ;
        RECT 136.505 137.945 136.775 138.275 ;
        RECT 137.420 137.925 137.770 138.575 ;
        RECT 134.250 137.575 136.735 137.765 ;
        RECT 137.940 137.755 138.170 138.745 ;
        RECT 134.255 137.035 135.000 137.405 ;
        RECT 135.565 137.215 135.820 137.575 ;
        RECT 136.000 137.035 136.330 137.405 ;
        RECT 136.510 137.215 136.735 137.575 ;
        RECT 137.505 137.585 138.170 137.755 ;
        RECT 137.505 137.295 137.675 137.585 ;
        RECT 137.845 137.035 138.175 137.415 ;
        RECT 138.345 137.295 138.530 139.415 ;
        RECT 138.770 139.125 139.035 139.585 ;
        RECT 139.205 138.990 139.455 139.415 ;
        RECT 139.665 139.140 140.770 139.310 ;
        RECT 139.150 138.860 139.455 138.990 ;
        RECT 138.700 137.665 138.980 138.615 ;
        RECT 139.150 137.755 139.320 138.860 ;
        RECT 139.490 138.075 139.730 138.670 ;
        RECT 139.900 138.605 140.430 138.970 ;
        RECT 139.900 137.905 140.070 138.605 ;
        RECT 140.600 138.525 140.770 139.140 ;
        RECT 140.940 138.785 141.110 139.585 ;
        RECT 141.280 139.085 141.530 139.415 ;
        RECT 141.755 139.115 142.640 139.285 ;
        RECT 140.600 138.435 141.110 138.525 ;
        RECT 139.150 137.625 139.375 137.755 ;
        RECT 139.545 137.685 140.070 137.905 ;
        RECT 140.240 138.265 141.110 138.435 ;
        RECT 138.785 137.035 139.035 137.495 ;
        RECT 139.205 137.485 139.375 137.625 ;
        RECT 140.240 137.485 140.410 138.265 ;
        RECT 140.940 138.195 141.110 138.265 ;
        RECT 140.620 138.015 140.820 138.045 ;
        RECT 141.280 138.015 141.450 139.085 ;
        RECT 141.620 138.195 141.810 138.915 ;
        RECT 140.620 137.715 141.450 138.015 ;
        RECT 141.980 137.985 142.300 138.945 ;
        RECT 139.205 137.315 139.540 137.485 ;
        RECT 139.735 137.315 140.410 137.485 ;
        RECT 140.730 137.035 141.100 137.535 ;
        RECT 141.280 137.485 141.450 137.715 ;
        RECT 141.835 137.655 142.300 137.985 ;
        RECT 142.470 138.275 142.640 139.115 ;
        RECT 142.820 139.085 143.135 139.585 ;
        RECT 143.365 138.855 143.705 139.415 ;
        RECT 142.810 138.480 143.705 138.855 ;
        RECT 143.875 138.575 144.045 139.585 ;
        RECT 143.515 138.275 143.705 138.480 ;
        RECT 144.215 138.525 144.545 139.370 ;
        RECT 144.215 138.445 144.605 138.525 ;
        RECT 144.390 138.395 144.605 138.445 ;
        RECT 142.470 137.945 143.345 138.275 ;
        RECT 143.515 137.945 144.265 138.275 ;
        RECT 142.470 137.485 142.640 137.945 ;
        RECT 143.515 137.775 143.715 137.945 ;
        RECT 144.435 137.815 144.605 138.395 ;
        RECT 145.695 138.495 146.905 139.585 ;
        RECT 145.695 137.955 146.215 138.495 ;
        RECT 144.380 137.775 144.605 137.815 ;
        RECT 146.385 137.785 146.905 138.325 ;
        RECT 141.280 137.315 141.685 137.485 ;
        RECT 141.855 137.315 142.640 137.485 ;
        RECT 142.915 137.035 143.125 137.565 ;
        RECT 143.385 137.250 143.715 137.775 ;
        RECT 144.225 137.690 144.605 137.775 ;
        RECT 143.885 137.035 144.055 137.645 ;
        RECT 144.225 137.255 144.555 137.690 ;
        RECT 145.695 137.035 146.905 137.785 ;
        RECT 17.270 136.865 146.990 137.035 ;
        RECT 17.355 136.115 18.565 136.865 ;
        RECT 17.355 135.575 17.875 136.115 ;
        RECT 18.740 136.025 19.000 136.865 ;
        RECT 19.175 136.120 19.430 136.695 ;
        RECT 19.600 136.485 19.930 136.865 ;
        RECT 20.145 136.315 20.315 136.695 ;
        RECT 19.600 136.145 20.315 136.315 ;
        RECT 20.665 136.315 20.835 136.695 ;
        RECT 21.015 136.485 21.345 136.865 ;
        RECT 20.665 136.145 21.330 136.315 ;
        RECT 21.525 136.190 21.785 136.695 ;
        RECT 18.045 135.405 18.565 135.945 ;
        RECT 17.355 134.315 18.565 135.405 ;
        RECT 18.740 134.315 19.000 135.465 ;
        RECT 19.175 135.390 19.345 136.120 ;
        RECT 19.600 135.955 19.770 136.145 ;
        RECT 19.515 135.625 19.770 135.955 ;
        RECT 19.600 135.415 19.770 135.625 ;
        RECT 20.050 135.595 20.405 135.965 ;
        RECT 20.595 135.595 20.935 135.965 ;
        RECT 21.160 135.890 21.330 136.145 ;
        RECT 21.160 135.560 21.435 135.890 ;
        RECT 21.160 135.415 21.330 135.560 ;
        RECT 19.175 134.485 19.430 135.390 ;
        RECT 19.600 135.245 20.315 135.415 ;
        RECT 19.600 134.315 19.930 135.075 ;
        RECT 20.145 134.485 20.315 135.245 ;
        RECT 20.655 135.245 21.330 135.415 ;
        RECT 21.605 135.390 21.785 136.190 ;
        RECT 21.955 136.095 24.545 136.865 ;
        RECT 24.805 136.315 24.975 136.605 ;
        RECT 25.145 136.485 25.475 136.865 ;
        RECT 24.805 136.145 25.470 136.315 ;
        RECT 21.955 135.575 23.165 136.095 ;
        RECT 23.335 135.405 24.545 135.925 ;
        RECT 20.655 134.485 20.835 135.245 ;
        RECT 21.015 134.315 21.345 135.075 ;
        RECT 21.515 134.485 21.785 135.390 ;
        RECT 21.955 134.315 24.545 135.405 ;
        RECT 24.720 135.325 25.070 135.975 ;
        RECT 25.240 135.155 25.470 136.145 ;
        RECT 24.805 134.985 25.470 135.155 ;
        RECT 24.805 134.485 24.975 134.985 ;
        RECT 25.145 134.315 25.475 134.815 ;
        RECT 25.645 134.485 25.830 136.605 ;
        RECT 26.085 136.405 26.335 136.865 ;
        RECT 26.505 136.415 26.840 136.585 ;
        RECT 27.035 136.415 27.710 136.585 ;
        RECT 26.505 136.275 26.675 136.415 ;
        RECT 26.000 135.285 26.280 136.235 ;
        RECT 26.450 136.145 26.675 136.275 ;
        RECT 26.450 135.040 26.620 136.145 ;
        RECT 26.845 135.995 27.370 136.215 ;
        RECT 26.790 135.230 27.030 135.825 ;
        RECT 27.200 135.295 27.370 135.995 ;
        RECT 27.540 135.635 27.710 136.415 ;
        RECT 28.030 136.365 28.400 136.865 ;
        RECT 28.580 136.415 28.985 136.585 ;
        RECT 29.155 136.415 29.940 136.585 ;
        RECT 28.580 136.185 28.750 136.415 ;
        RECT 27.920 135.885 28.750 136.185 ;
        RECT 29.135 135.915 29.600 136.245 ;
        RECT 27.920 135.855 28.120 135.885 ;
        RECT 28.240 135.635 28.410 135.705 ;
        RECT 27.540 135.465 28.410 135.635 ;
        RECT 27.900 135.375 28.410 135.465 ;
        RECT 26.450 134.910 26.755 135.040 ;
        RECT 27.200 134.930 27.730 135.295 ;
        RECT 26.070 134.315 26.335 134.775 ;
        RECT 26.505 134.485 26.755 134.910 ;
        RECT 27.900 134.760 28.070 135.375 ;
        RECT 26.965 134.590 28.070 134.760 ;
        RECT 28.240 134.315 28.410 135.115 ;
        RECT 28.580 134.815 28.750 135.885 ;
        RECT 28.920 134.985 29.110 135.705 ;
        RECT 29.280 134.955 29.600 135.915 ;
        RECT 29.770 135.955 29.940 136.415 ;
        RECT 30.215 136.335 30.425 136.865 ;
        RECT 30.685 136.125 31.015 136.650 ;
        RECT 31.185 136.255 31.355 136.865 ;
        RECT 31.525 136.210 31.855 136.645 ;
        RECT 31.525 136.125 31.905 136.210 ;
        RECT 30.815 135.955 31.015 136.125 ;
        RECT 31.680 136.085 31.905 136.125 ;
        RECT 29.770 135.625 30.645 135.955 ;
        RECT 30.815 135.625 31.565 135.955 ;
        RECT 28.580 134.485 28.830 134.815 ;
        RECT 29.770 134.785 29.940 135.625 ;
        RECT 30.815 135.420 31.005 135.625 ;
        RECT 31.735 135.505 31.905 136.085 ;
        RECT 32.115 136.045 32.345 136.865 ;
        RECT 32.515 136.065 32.845 136.695 ;
        RECT 32.095 135.625 32.425 135.875 ;
        RECT 31.690 135.455 31.905 135.505 ;
        RECT 32.595 135.465 32.845 136.065 ;
        RECT 33.015 136.045 33.225 136.865 ;
        RECT 33.455 136.320 38.800 136.865 ;
        RECT 35.040 135.490 35.380 136.320 ;
        RECT 38.975 136.095 42.485 136.865 ;
        RECT 43.115 136.140 43.405 136.865 ;
        RECT 43.575 136.320 48.920 136.865 ;
        RECT 49.095 136.320 54.440 136.865 ;
        RECT 54.615 136.320 59.960 136.865 ;
        RECT 30.110 135.045 31.005 135.420 ;
        RECT 31.515 135.375 31.905 135.455 ;
        RECT 29.055 134.615 29.940 134.785 ;
        RECT 30.120 134.315 30.435 134.815 ;
        RECT 30.665 134.485 31.005 135.045 ;
        RECT 31.175 134.315 31.345 135.325 ;
        RECT 31.515 134.530 31.845 135.375 ;
        RECT 32.115 134.315 32.345 135.455 ;
        RECT 32.515 134.485 32.845 135.465 ;
        RECT 33.015 134.315 33.225 135.455 ;
        RECT 36.860 134.750 37.210 136.000 ;
        RECT 38.975 135.575 40.625 136.095 ;
        RECT 40.795 135.405 42.485 135.925 ;
        RECT 45.160 135.490 45.500 136.320 ;
        RECT 33.455 134.315 38.800 134.750 ;
        RECT 38.975 134.315 42.485 135.405 ;
        RECT 43.115 134.315 43.405 135.480 ;
        RECT 46.980 134.750 47.330 136.000 ;
        RECT 50.680 135.490 51.020 136.320 ;
        RECT 52.500 134.750 52.850 136.000 ;
        RECT 56.200 135.490 56.540 136.320 ;
        RECT 60.135 136.095 63.645 136.865 ;
        RECT 63.815 136.115 65.025 136.865 ;
        RECT 58.020 134.750 58.370 136.000 ;
        RECT 60.135 135.575 61.785 136.095 ;
        RECT 61.955 135.405 63.645 135.925 ;
        RECT 63.815 135.575 64.335 136.115 ;
        RECT 65.205 136.055 65.475 136.865 ;
        RECT 65.645 136.055 65.975 136.695 ;
        RECT 66.145 136.055 66.385 136.865 ;
        RECT 66.610 136.125 67.225 136.695 ;
        RECT 67.395 136.355 67.610 136.865 ;
        RECT 67.840 136.355 68.120 136.685 ;
        RECT 68.300 136.355 68.540 136.865 ;
        RECT 64.505 135.405 65.025 135.945 ;
        RECT 65.195 135.625 65.545 135.875 ;
        RECT 65.715 135.455 65.885 136.055 ;
        RECT 66.055 135.625 66.405 135.875 ;
        RECT 43.575 134.315 48.920 134.750 ;
        RECT 49.095 134.315 54.440 134.750 ;
        RECT 54.615 134.315 59.960 134.750 ;
        RECT 60.135 134.315 63.645 135.405 ;
        RECT 63.815 134.315 65.025 135.405 ;
        RECT 65.205 134.315 65.535 135.455 ;
        RECT 65.715 135.285 66.395 135.455 ;
        RECT 66.065 134.500 66.395 135.285 ;
        RECT 66.610 135.105 66.925 136.125 ;
        RECT 67.095 135.455 67.265 135.955 ;
        RECT 67.515 135.625 67.780 136.185 ;
        RECT 67.950 135.455 68.120 136.355 ;
        RECT 68.290 135.625 68.645 136.185 ;
        RECT 68.875 136.140 69.165 136.865 ;
        RECT 69.425 136.315 69.595 136.605 ;
        RECT 69.765 136.485 70.095 136.865 ;
        RECT 69.425 136.145 70.090 136.315 ;
        RECT 67.095 135.285 68.520 135.455 ;
        RECT 66.610 134.485 67.145 135.105 ;
        RECT 67.315 134.315 67.645 135.115 ;
        RECT 68.130 135.110 68.520 135.285 ;
        RECT 68.875 134.315 69.165 135.480 ;
        RECT 69.340 135.325 69.690 135.975 ;
        RECT 69.860 135.155 70.090 136.145 ;
        RECT 69.425 134.985 70.090 135.155 ;
        RECT 69.425 134.485 69.595 134.985 ;
        RECT 69.765 134.315 70.095 134.815 ;
        RECT 70.265 134.485 70.450 136.605 ;
        RECT 70.705 136.405 70.955 136.865 ;
        RECT 71.125 136.415 71.460 136.585 ;
        RECT 71.655 136.415 72.330 136.585 ;
        RECT 71.125 136.275 71.295 136.415 ;
        RECT 70.620 135.285 70.900 136.235 ;
        RECT 71.070 136.145 71.295 136.275 ;
        RECT 71.070 135.040 71.240 136.145 ;
        RECT 71.465 135.995 71.990 136.215 ;
        RECT 71.410 135.230 71.650 135.825 ;
        RECT 71.820 135.295 71.990 135.995 ;
        RECT 72.160 135.635 72.330 136.415 ;
        RECT 72.650 136.365 73.020 136.865 ;
        RECT 73.200 136.415 73.605 136.585 ;
        RECT 73.775 136.415 74.560 136.585 ;
        RECT 73.200 136.185 73.370 136.415 ;
        RECT 72.540 135.885 73.370 136.185 ;
        RECT 73.755 135.915 74.220 136.245 ;
        RECT 72.540 135.855 72.740 135.885 ;
        RECT 72.860 135.635 73.030 135.705 ;
        RECT 72.160 135.465 73.030 135.635 ;
        RECT 72.520 135.375 73.030 135.465 ;
        RECT 71.070 134.910 71.375 135.040 ;
        RECT 71.820 134.930 72.350 135.295 ;
        RECT 70.690 134.315 70.955 134.775 ;
        RECT 71.125 134.485 71.375 134.910 ;
        RECT 72.520 134.760 72.690 135.375 ;
        RECT 71.585 134.590 72.690 134.760 ;
        RECT 72.860 134.315 73.030 135.115 ;
        RECT 73.200 134.815 73.370 135.885 ;
        RECT 73.540 134.985 73.730 135.705 ;
        RECT 73.900 134.955 74.220 135.915 ;
        RECT 74.390 135.955 74.560 136.415 ;
        RECT 74.835 136.335 75.045 136.865 ;
        RECT 75.305 136.125 75.635 136.650 ;
        RECT 75.805 136.255 75.975 136.865 ;
        RECT 76.145 136.210 76.475 136.645 ;
        RECT 76.145 136.125 76.525 136.210 ;
        RECT 75.435 135.955 75.635 136.125 ;
        RECT 76.300 136.085 76.525 136.125 ;
        RECT 74.390 135.625 75.265 135.955 ;
        RECT 75.435 135.625 76.185 135.955 ;
        RECT 73.200 134.485 73.450 134.815 ;
        RECT 74.390 134.785 74.560 135.625 ;
        RECT 75.435 135.420 75.625 135.625 ;
        RECT 76.355 135.505 76.525 136.085 ;
        RECT 76.695 136.065 77.390 136.695 ;
        RECT 77.595 136.065 77.905 136.865 ;
        RECT 78.075 136.115 79.285 136.865 ;
        RECT 76.715 135.625 77.050 135.875 ;
        RECT 76.310 135.455 76.525 135.505 ;
        RECT 77.220 135.465 77.390 136.065 ;
        RECT 77.560 135.625 77.895 135.895 ;
        RECT 78.075 135.575 78.595 136.115 ;
        RECT 79.455 136.045 79.715 136.865 ;
        RECT 79.885 136.045 80.215 136.465 ;
        RECT 80.395 136.295 80.655 136.695 ;
        RECT 80.825 136.465 81.155 136.865 ;
        RECT 81.325 136.295 81.495 136.645 ;
        RECT 81.665 136.465 82.040 136.865 ;
        RECT 80.395 136.125 82.060 136.295 ;
        RECT 82.230 136.190 82.505 136.535 ;
        RECT 79.965 135.955 80.215 136.045 ;
        RECT 81.890 135.955 82.060 136.125 ;
        RECT 74.730 135.045 75.625 135.420 ;
        RECT 76.135 135.375 76.525 135.455 ;
        RECT 73.675 134.615 74.560 134.785 ;
        RECT 74.740 134.315 75.055 134.815 ;
        RECT 75.285 134.485 75.625 135.045 ;
        RECT 75.795 134.315 75.965 135.325 ;
        RECT 76.135 134.530 76.465 135.375 ;
        RECT 76.695 134.315 76.955 135.455 ;
        RECT 77.125 134.485 77.455 135.465 ;
        RECT 77.625 134.315 77.905 135.455 ;
        RECT 78.765 135.405 79.285 135.945 ;
        RECT 79.460 135.625 79.795 135.875 ;
        RECT 79.965 135.625 80.680 135.955 ;
        RECT 80.895 135.625 81.720 135.955 ;
        RECT 81.890 135.625 82.165 135.955 ;
        RECT 78.075 134.315 79.285 135.405 ;
        RECT 79.455 134.315 79.715 135.455 ;
        RECT 79.965 135.065 80.135 135.625 ;
        RECT 80.395 135.165 80.725 135.455 ;
        RECT 80.895 135.335 81.140 135.625 ;
        RECT 81.890 135.455 82.060 135.625 ;
        RECT 82.335 135.455 82.505 136.190 ;
        RECT 82.675 136.045 82.935 136.865 ;
        RECT 83.105 136.045 83.435 136.465 ;
        RECT 83.615 136.295 83.875 136.695 ;
        RECT 84.045 136.465 84.375 136.865 ;
        RECT 84.545 136.295 84.715 136.645 ;
        RECT 84.885 136.465 85.260 136.865 ;
        RECT 83.615 136.125 85.280 136.295 ;
        RECT 85.450 136.190 85.725 136.535 ;
        RECT 83.185 135.955 83.435 136.045 ;
        RECT 85.110 135.955 85.280 136.125 ;
        RECT 82.680 135.625 83.015 135.875 ;
        RECT 83.185 135.625 83.900 135.955 ;
        RECT 84.115 135.625 84.940 135.955 ;
        RECT 85.110 135.625 85.385 135.955 ;
        RECT 81.400 135.285 82.060 135.455 ;
        RECT 81.400 135.165 81.570 135.285 ;
        RECT 80.395 134.995 81.570 135.165 ;
        RECT 79.955 134.495 81.570 134.825 ;
        RECT 81.740 134.315 82.020 135.115 ;
        RECT 82.230 134.485 82.505 135.455 ;
        RECT 82.675 134.315 82.935 135.455 ;
        RECT 83.185 135.065 83.355 135.625 ;
        RECT 83.615 135.165 83.945 135.455 ;
        RECT 84.115 135.335 84.360 135.625 ;
        RECT 85.110 135.455 85.280 135.625 ;
        RECT 85.555 135.455 85.725 136.190 ;
        RECT 86.905 136.315 87.075 136.605 ;
        RECT 87.245 136.485 87.575 136.865 ;
        RECT 86.905 136.145 87.570 136.315 ;
        RECT 84.620 135.285 85.280 135.455 ;
        RECT 84.620 135.165 84.790 135.285 ;
        RECT 83.615 134.995 84.790 135.165 ;
        RECT 83.175 134.495 84.790 134.825 ;
        RECT 84.960 134.315 85.240 135.115 ;
        RECT 85.450 134.485 85.725 135.455 ;
        RECT 86.820 135.325 87.170 135.975 ;
        RECT 87.340 135.155 87.570 136.145 ;
        RECT 86.905 134.985 87.570 135.155 ;
        RECT 86.905 134.485 87.075 134.985 ;
        RECT 87.245 134.315 87.575 134.815 ;
        RECT 87.745 134.485 87.930 136.605 ;
        RECT 88.185 136.405 88.435 136.865 ;
        RECT 88.605 136.415 88.940 136.585 ;
        RECT 89.135 136.415 89.810 136.585 ;
        RECT 88.605 136.275 88.775 136.415 ;
        RECT 88.100 135.285 88.380 136.235 ;
        RECT 88.550 136.145 88.775 136.275 ;
        RECT 88.550 135.040 88.720 136.145 ;
        RECT 88.945 135.995 89.470 136.215 ;
        RECT 88.890 135.230 89.130 135.825 ;
        RECT 89.300 135.295 89.470 135.995 ;
        RECT 89.640 135.635 89.810 136.415 ;
        RECT 90.130 136.365 90.500 136.865 ;
        RECT 90.680 136.415 91.085 136.585 ;
        RECT 91.255 136.415 92.040 136.585 ;
        RECT 90.680 136.185 90.850 136.415 ;
        RECT 90.020 135.885 90.850 136.185 ;
        RECT 91.235 135.915 91.700 136.245 ;
        RECT 90.020 135.855 90.220 135.885 ;
        RECT 90.340 135.635 90.510 135.705 ;
        RECT 89.640 135.465 90.510 135.635 ;
        RECT 90.000 135.375 90.510 135.465 ;
        RECT 88.550 134.910 88.855 135.040 ;
        RECT 89.300 134.930 89.830 135.295 ;
        RECT 88.170 134.315 88.435 134.775 ;
        RECT 88.605 134.485 88.855 134.910 ;
        RECT 90.000 134.760 90.170 135.375 ;
        RECT 89.065 134.590 90.170 134.760 ;
        RECT 90.340 134.315 90.510 135.115 ;
        RECT 90.680 134.815 90.850 135.885 ;
        RECT 91.020 134.985 91.210 135.705 ;
        RECT 91.380 134.955 91.700 135.915 ;
        RECT 91.870 135.955 92.040 136.415 ;
        RECT 92.315 136.335 92.525 136.865 ;
        RECT 92.785 136.125 93.115 136.650 ;
        RECT 93.285 136.255 93.455 136.865 ;
        RECT 93.625 136.210 93.955 136.645 ;
        RECT 94.125 136.350 94.295 136.865 ;
        RECT 93.625 136.125 94.005 136.210 ;
        RECT 94.635 136.140 94.925 136.865 ;
        RECT 92.915 135.955 93.115 136.125 ;
        RECT 93.780 136.085 94.005 136.125 ;
        RECT 91.870 135.625 92.745 135.955 ;
        RECT 92.915 135.625 93.665 135.955 ;
        RECT 90.680 134.485 90.930 134.815 ;
        RECT 91.870 134.785 92.040 135.625 ;
        RECT 92.915 135.420 93.105 135.625 ;
        RECT 93.835 135.505 94.005 136.085 ;
        RECT 95.095 136.095 98.605 136.865 ;
        RECT 99.745 136.210 100.075 136.645 ;
        RECT 100.245 136.255 100.415 136.865 ;
        RECT 99.695 136.125 100.075 136.210 ;
        RECT 100.585 136.125 100.915 136.650 ;
        RECT 101.175 136.335 101.385 136.865 ;
        RECT 101.660 136.415 102.445 136.585 ;
        RECT 102.615 136.415 103.020 136.585 ;
        RECT 95.095 135.575 96.745 136.095 ;
        RECT 99.695 136.085 99.920 136.125 ;
        RECT 93.790 135.455 94.005 135.505 ;
        RECT 92.210 135.045 93.105 135.420 ;
        RECT 93.615 135.375 94.005 135.455 ;
        RECT 91.155 134.615 92.040 134.785 ;
        RECT 92.220 134.315 92.535 134.815 ;
        RECT 92.765 134.485 93.105 135.045 ;
        RECT 93.275 134.315 93.445 135.325 ;
        RECT 93.615 134.530 93.945 135.375 ;
        RECT 94.115 134.315 94.285 135.230 ;
        RECT 94.635 134.315 94.925 135.480 ;
        RECT 96.915 135.405 98.605 135.925 ;
        RECT 95.095 134.315 98.605 135.405 ;
        RECT 99.695 135.505 99.865 136.085 ;
        RECT 100.585 135.955 100.785 136.125 ;
        RECT 101.660 135.955 101.830 136.415 ;
        RECT 100.035 135.625 100.785 135.955 ;
        RECT 100.955 135.625 101.830 135.955 ;
        RECT 99.695 135.455 99.910 135.505 ;
        RECT 99.695 135.375 100.085 135.455 ;
        RECT 99.755 134.530 100.085 135.375 ;
        RECT 100.595 135.420 100.785 135.625 ;
        RECT 100.255 134.315 100.425 135.325 ;
        RECT 100.595 135.045 101.490 135.420 ;
        RECT 100.595 134.485 100.935 135.045 ;
        RECT 101.165 134.315 101.480 134.815 ;
        RECT 101.660 134.785 101.830 135.625 ;
        RECT 102.000 135.915 102.465 136.245 ;
        RECT 102.850 136.185 103.020 136.415 ;
        RECT 103.200 136.365 103.570 136.865 ;
        RECT 103.890 136.415 104.565 136.585 ;
        RECT 104.760 136.415 105.095 136.585 ;
        RECT 102.000 134.955 102.320 135.915 ;
        RECT 102.850 135.885 103.680 136.185 ;
        RECT 102.490 134.985 102.680 135.705 ;
        RECT 102.850 134.815 103.020 135.885 ;
        RECT 103.480 135.855 103.680 135.885 ;
        RECT 103.190 135.635 103.360 135.705 ;
        RECT 103.890 135.635 104.060 136.415 ;
        RECT 104.925 136.275 105.095 136.415 ;
        RECT 105.265 136.405 105.515 136.865 ;
        RECT 103.190 135.465 104.060 135.635 ;
        RECT 104.230 135.995 104.755 136.215 ;
        RECT 104.925 136.145 105.150 136.275 ;
        RECT 103.190 135.375 103.700 135.465 ;
        RECT 101.660 134.615 102.545 134.785 ;
        RECT 102.770 134.485 103.020 134.815 ;
        RECT 103.190 134.315 103.360 135.115 ;
        RECT 103.530 134.760 103.700 135.375 ;
        RECT 104.230 135.295 104.400 135.995 ;
        RECT 103.870 134.930 104.400 135.295 ;
        RECT 104.570 135.230 104.810 135.825 ;
        RECT 104.980 135.040 105.150 136.145 ;
        RECT 105.320 135.285 105.600 136.235 ;
        RECT 104.845 134.910 105.150 135.040 ;
        RECT 103.530 134.590 104.635 134.760 ;
        RECT 104.845 134.485 105.095 134.910 ;
        RECT 105.265 134.315 105.530 134.775 ;
        RECT 105.770 134.485 105.955 136.605 ;
        RECT 106.125 136.485 106.455 136.865 ;
        RECT 106.625 136.315 106.795 136.605 ;
        RECT 106.130 136.145 106.795 136.315 ;
        RECT 107.145 136.315 107.315 136.605 ;
        RECT 107.485 136.485 107.815 136.865 ;
        RECT 107.145 136.145 107.810 136.315 ;
        RECT 106.130 135.155 106.360 136.145 ;
        RECT 106.530 135.325 106.880 135.975 ;
        RECT 107.060 135.325 107.410 135.975 ;
        RECT 107.580 135.155 107.810 136.145 ;
        RECT 106.130 134.985 106.795 135.155 ;
        RECT 106.125 134.315 106.455 134.815 ;
        RECT 106.625 134.485 106.795 134.985 ;
        RECT 107.145 134.985 107.810 135.155 ;
        RECT 107.145 134.485 107.315 134.985 ;
        RECT 107.485 134.315 107.815 134.815 ;
        RECT 107.985 134.485 108.170 136.605 ;
        RECT 108.425 136.405 108.675 136.865 ;
        RECT 108.845 136.415 109.180 136.585 ;
        RECT 109.375 136.415 110.050 136.585 ;
        RECT 108.845 136.275 109.015 136.415 ;
        RECT 108.340 135.285 108.620 136.235 ;
        RECT 108.790 136.145 109.015 136.275 ;
        RECT 108.790 135.040 108.960 136.145 ;
        RECT 109.185 135.995 109.710 136.215 ;
        RECT 109.130 135.230 109.370 135.825 ;
        RECT 109.540 135.295 109.710 135.995 ;
        RECT 109.880 135.635 110.050 136.415 ;
        RECT 110.370 136.365 110.740 136.865 ;
        RECT 110.920 136.415 111.325 136.585 ;
        RECT 111.495 136.415 112.280 136.585 ;
        RECT 110.920 136.185 111.090 136.415 ;
        RECT 110.260 135.885 111.090 136.185 ;
        RECT 111.475 135.915 111.940 136.245 ;
        RECT 110.260 135.855 110.460 135.885 ;
        RECT 110.580 135.635 110.750 135.705 ;
        RECT 109.880 135.465 110.750 135.635 ;
        RECT 110.240 135.375 110.750 135.465 ;
        RECT 108.790 134.910 109.095 135.040 ;
        RECT 109.540 134.930 110.070 135.295 ;
        RECT 108.410 134.315 108.675 134.775 ;
        RECT 108.845 134.485 109.095 134.910 ;
        RECT 110.240 134.760 110.410 135.375 ;
        RECT 109.305 134.590 110.410 134.760 ;
        RECT 110.580 134.315 110.750 135.115 ;
        RECT 110.920 134.815 111.090 135.885 ;
        RECT 111.260 134.985 111.450 135.705 ;
        RECT 111.620 134.955 111.940 135.915 ;
        RECT 112.110 135.955 112.280 136.415 ;
        RECT 112.555 136.335 112.765 136.865 ;
        RECT 113.025 136.125 113.355 136.650 ;
        RECT 113.525 136.255 113.695 136.865 ;
        RECT 113.865 136.210 114.195 136.645 ;
        RECT 113.865 136.125 114.245 136.210 ;
        RECT 113.155 135.955 113.355 136.125 ;
        RECT 114.020 136.085 114.245 136.125 ;
        RECT 112.110 135.625 112.985 135.955 ;
        RECT 113.155 135.625 113.905 135.955 ;
        RECT 110.920 134.485 111.170 134.815 ;
        RECT 112.110 134.785 112.280 135.625 ;
        RECT 113.155 135.420 113.345 135.625 ;
        RECT 114.075 135.505 114.245 136.085 ;
        RECT 114.415 136.095 116.085 136.865 ;
        RECT 114.415 135.575 115.165 136.095 ;
        RECT 114.030 135.455 114.245 135.505 ;
        RECT 112.450 135.045 113.345 135.420 ;
        RECT 113.855 135.375 114.245 135.455 ;
        RECT 115.335 135.405 116.085 135.925 ;
        RECT 111.395 134.615 112.280 134.785 ;
        RECT 112.460 134.315 112.775 134.815 ;
        RECT 113.005 134.485 113.345 135.045 ;
        RECT 113.515 134.315 113.685 135.325 ;
        RECT 113.855 134.530 114.185 135.375 ;
        RECT 114.415 134.315 116.085 135.405 ;
        RECT 116.715 135.920 117.055 136.695 ;
        RECT 117.225 136.405 117.395 136.865 ;
        RECT 117.635 136.430 117.995 136.695 ;
        RECT 117.635 136.425 117.990 136.430 ;
        RECT 117.635 136.415 117.985 136.425 ;
        RECT 117.635 136.410 117.980 136.415 ;
        RECT 117.635 136.400 117.975 136.410 ;
        RECT 118.625 136.405 118.795 136.865 ;
        RECT 117.635 136.395 117.970 136.400 ;
        RECT 117.635 136.385 117.960 136.395 ;
        RECT 117.635 136.375 117.950 136.385 ;
        RECT 117.635 136.235 117.935 136.375 ;
        RECT 117.225 136.045 117.935 136.235 ;
        RECT 118.125 136.235 118.455 136.315 ;
        RECT 118.965 136.235 119.305 136.695 ;
        RECT 118.125 136.045 119.305 136.235 ;
        RECT 120.395 136.140 120.685 136.865 ;
        RECT 120.855 136.125 121.240 136.695 ;
        RECT 121.410 136.405 121.735 136.865 ;
        RECT 122.255 136.235 122.535 136.695 ;
        RECT 116.715 134.485 116.995 135.920 ;
        RECT 117.225 135.475 117.510 136.045 ;
        RECT 117.695 135.645 118.165 135.875 ;
        RECT 118.335 135.855 118.665 135.875 ;
        RECT 118.335 135.675 118.785 135.855 ;
        RECT 118.975 135.675 119.305 135.875 ;
        RECT 117.225 135.260 118.375 135.475 ;
        RECT 117.165 134.315 117.875 135.090 ;
        RECT 118.045 134.485 118.375 135.260 ;
        RECT 118.570 134.560 118.785 135.675 ;
        RECT 119.075 135.335 119.305 135.675 ;
        RECT 118.965 134.315 119.295 135.035 ;
        RECT 120.395 134.315 120.685 135.480 ;
        RECT 120.855 135.455 121.135 136.125 ;
        RECT 121.410 136.065 122.535 136.235 ;
        RECT 121.410 135.955 121.860 136.065 ;
        RECT 121.305 135.625 121.860 135.955 ;
        RECT 122.725 135.895 123.125 136.695 ;
        RECT 123.525 136.405 123.795 136.865 ;
        RECT 123.965 136.235 124.250 136.695 ;
        RECT 120.855 134.485 121.240 135.455 ;
        RECT 121.410 135.165 121.860 135.625 ;
        RECT 122.030 135.335 123.125 135.895 ;
        RECT 121.410 134.945 122.535 135.165 ;
        RECT 121.410 134.315 121.735 134.775 ;
        RECT 122.255 134.485 122.535 134.945 ;
        RECT 122.725 134.485 123.125 135.335 ;
        RECT 123.295 136.065 124.250 136.235 ;
        RECT 124.535 136.125 124.920 136.695 ;
        RECT 125.090 136.405 125.415 136.865 ;
        RECT 125.935 136.235 126.215 136.695 ;
        RECT 123.295 135.165 123.505 136.065 ;
        RECT 123.675 135.335 124.365 135.895 ;
        RECT 124.535 135.455 124.815 136.125 ;
        RECT 125.090 136.065 126.215 136.235 ;
        RECT 125.090 135.955 125.540 136.065 ;
        RECT 124.985 135.625 125.540 135.955 ;
        RECT 126.405 135.895 126.805 136.695 ;
        RECT 127.205 136.405 127.475 136.865 ;
        RECT 127.645 136.235 127.930 136.695 ;
        RECT 123.295 134.945 124.250 135.165 ;
        RECT 123.525 134.315 123.795 134.775 ;
        RECT 123.965 134.485 124.250 134.945 ;
        RECT 124.535 134.485 124.920 135.455 ;
        RECT 125.090 135.165 125.540 135.625 ;
        RECT 125.710 135.335 126.805 135.895 ;
        RECT 125.090 134.945 126.215 135.165 ;
        RECT 125.090 134.315 125.415 134.775 ;
        RECT 125.935 134.485 126.215 134.945 ;
        RECT 126.405 134.485 126.805 135.335 ;
        RECT 126.975 136.065 127.930 136.235 ;
        RECT 126.975 135.165 127.185 136.065 ;
        RECT 127.355 135.335 128.045 135.895 ;
        RECT 128.680 135.265 129.015 136.685 ;
        RECT 129.195 136.495 129.940 136.865 ;
        RECT 130.505 136.325 130.760 136.685 ;
        RECT 130.940 136.495 131.270 136.865 ;
        RECT 131.450 136.325 131.675 136.685 ;
        RECT 129.190 136.135 131.675 136.325 ;
        RECT 129.190 135.445 129.415 136.135 ;
        RECT 132.170 136.055 132.415 136.660 ;
        RECT 132.635 136.330 133.145 136.865 ;
        RECT 129.615 135.625 129.895 135.955 ;
        RECT 130.075 135.625 130.650 135.955 ;
        RECT 130.830 135.625 131.265 135.955 ;
        RECT 131.445 135.625 131.715 135.955 ;
        RECT 131.895 135.885 133.125 136.055 ;
        RECT 129.190 135.265 131.685 135.445 ;
        RECT 126.975 134.945 127.930 135.165 ;
        RECT 127.205 134.315 127.475 134.775 ;
        RECT 127.645 134.485 127.930 134.945 ;
        RECT 128.680 134.495 128.945 135.265 ;
        RECT 129.115 134.315 129.445 135.035 ;
        RECT 129.635 134.855 130.825 135.085 ;
        RECT 129.635 134.495 129.895 134.855 ;
        RECT 130.065 134.315 130.395 134.685 ;
        RECT 130.565 134.495 130.825 134.855 ;
        RECT 131.395 134.495 131.685 135.265 ;
        RECT 131.895 135.075 132.235 135.885 ;
        RECT 132.405 135.320 133.155 135.510 ;
        RECT 131.895 134.665 132.410 135.075 ;
        RECT 132.645 134.315 132.815 135.075 ;
        RECT 132.985 134.655 133.155 135.320 ;
        RECT 133.325 135.335 133.515 136.695 ;
        RECT 133.685 135.845 133.960 136.695 ;
        RECT 134.150 136.330 134.680 136.695 ;
        RECT 135.105 136.465 135.435 136.865 ;
        RECT 134.505 136.295 134.680 136.330 ;
        RECT 133.685 135.675 133.965 135.845 ;
        RECT 133.685 135.535 133.960 135.675 ;
        RECT 134.165 135.335 134.335 136.135 ;
        RECT 133.325 135.165 134.335 135.335 ;
        RECT 134.505 136.125 135.435 136.295 ;
        RECT 135.605 136.125 135.860 136.695 ;
        RECT 136.125 136.315 136.295 136.605 ;
        RECT 136.465 136.485 136.795 136.865 ;
        RECT 136.125 136.145 136.790 136.315 ;
        RECT 134.505 134.995 134.675 136.125 ;
        RECT 135.265 135.955 135.435 136.125 ;
        RECT 133.550 134.825 134.675 134.995 ;
        RECT 134.845 135.625 135.040 135.955 ;
        RECT 135.265 135.625 135.520 135.955 ;
        RECT 134.845 134.655 135.015 135.625 ;
        RECT 135.690 135.455 135.860 136.125 ;
        RECT 132.985 134.485 135.015 134.655 ;
        RECT 135.185 134.315 135.355 135.455 ;
        RECT 135.525 134.485 135.860 135.455 ;
        RECT 136.040 135.325 136.390 135.975 ;
        RECT 136.560 135.155 136.790 136.145 ;
        RECT 136.125 134.985 136.790 135.155 ;
        RECT 136.125 134.485 136.295 134.985 ;
        RECT 136.465 134.315 136.795 134.815 ;
        RECT 136.965 134.485 137.150 136.605 ;
        RECT 137.405 136.405 137.655 136.865 ;
        RECT 137.825 136.415 138.160 136.585 ;
        RECT 138.355 136.415 139.030 136.585 ;
        RECT 137.825 136.275 137.995 136.415 ;
        RECT 137.320 135.285 137.600 136.235 ;
        RECT 137.770 136.145 137.995 136.275 ;
        RECT 137.770 135.040 137.940 136.145 ;
        RECT 138.165 135.995 138.690 136.215 ;
        RECT 138.110 135.230 138.350 135.825 ;
        RECT 138.520 135.295 138.690 135.995 ;
        RECT 138.860 135.635 139.030 136.415 ;
        RECT 139.350 136.365 139.720 136.865 ;
        RECT 139.900 136.415 140.305 136.585 ;
        RECT 140.475 136.415 141.260 136.585 ;
        RECT 139.900 136.185 140.070 136.415 ;
        RECT 139.240 135.885 140.070 136.185 ;
        RECT 140.455 135.915 140.920 136.245 ;
        RECT 139.240 135.855 139.440 135.885 ;
        RECT 139.560 135.635 139.730 135.705 ;
        RECT 138.860 135.465 139.730 135.635 ;
        RECT 139.220 135.375 139.730 135.465 ;
        RECT 137.770 134.910 138.075 135.040 ;
        RECT 138.520 134.930 139.050 135.295 ;
        RECT 137.390 134.315 137.655 134.775 ;
        RECT 137.825 134.485 138.075 134.910 ;
        RECT 139.220 134.760 139.390 135.375 ;
        RECT 138.285 134.590 139.390 134.760 ;
        RECT 139.560 134.315 139.730 135.115 ;
        RECT 139.900 134.815 140.070 135.885 ;
        RECT 140.240 134.985 140.430 135.705 ;
        RECT 140.600 134.955 140.920 135.915 ;
        RECT 141.090 135.955 141.260 136.415 ;
        RECT 141.535 136.335 141.745 136.865 ;
        RECT 142.005 136.125 142.335 136.650 ;
        RECT 142.505 136.255 142.675 136.865 ;
        RECT 142.845 136.210 143.175 136.645 ;
        RECT 143.945 136.315 144.115 136.695 ;
        RECT 144.330 136.485 144.660 136.865 ;
        RECT 142.845 136.125 143.225 136.210 ;
        RECT 143.945 136.145 144.660 136.315 ;
        RECT 142.135 135.955 142.335 136.125 ;
        RECT 143.000 136.085 143.225 136.125 ;
        RECT 141.090 135.625 141.965 135.955 ;
        RECT 142.135 135.625 142.885 135.955 ;
        RECT 139.900 134.485 140.150 134.815 ;
        RECT 141.090 134.785 141.260 135.625 ;
        RECT 142.135 135.420 142.325 135.625 ;
        RECT 143.055 135.505 143.225 136.085 ;
        RECT 143.855 135.595 144.210 135.965 ;
        RECT 144.490 135.955 144.660 136.145 ;
        RECT 144.830 136.120 145.085 136.695 ;
        RECT 144.490 135.625 144.745 135.955 ;
        RECT 143.010 135.455 143.225 135.505 ;
        RECT 141.430 135.045 142.325 135.420 ;
        RECT 142.835 135.375 143.225 135.455 ;
        RECT 144.490 135.415 144.660 135.625 ;
        RECT 140.375 134.615 141.260 134.785 ;
        RECT 141.440 134.315 141.755 134.815 ;
        RECT 141.985 134.485 142.325 135.045 ;
        RECT 142.495 134.315 142.665 135.325 ;
        RECT 142.835 134.530 143.165 135.375 ;
        RECT 143.945 135.245 144.660 135.415 ;
        RECT 144.915 135.390 145.085 136.120 ;
        RECT 145.260 136.025 145.520 136.865 ;
        RECT 145.695 136.115 146.905 136.865 ;
        RECT 143.945 134.485 144.115 135.245 ;
        RECT 144.330 134.315 144.660 135.075 ;
        RECT 144.830 134.485 145.085 135.390 ;
        RECT 145.260 134.315 145.520 135.465 ;
        RECT 145.695 135.405 146.215 135.945 ;
        RECT 146.385 135.575 146.905 136.115 ;
        RECT 145.695 134.315 146.905 135.405 ;
        RECT 17.270 134.145 146.990 134.315 ;
        RECT 17.355 133.055 18.565 134.145 ;
        RECT 19.285 133.475 19.455 133.975 ;
        RECT 19.625 133.645 19.955 134.145 ;
        RECT 19.285 133.305 19.950 133.475 ;
        RECT 17.355 132.345 17.875 132.885 ;
        RECT 18.045 132.515 18.565 133.055 ;
        RECT 19.200 132.485 19.550 133.135 ;
        RECT 17.355 131.595 18.565 132.345 ;
        RECT 19.720 132.315 19.950 133.305 ;
        RECT 19.285 132.145 19.950 132.315 ;
        RECT 19.285 131.855 19.455 132.145 ;
        RECT 19.625 131.595 19.955 131.975 ;
        RECT 20.125 131.855 20.310 133.975 ;
        RECT 20.550 133.685 20.815 134.145 ;
        RECT 20.985 133.550 21.235 133.975 ;
        RECT 21.445 133.700 22.550 133.870 ;
        RECT 20.930 133.420 21.235 133.550 ;
        RECT 20.480 132.225 20.760 133.175 ;
        RECT 20.930 132.315 21.100 133.420 ;
        RECT 21.270 132.635 21.510 133.230 ;
        RECT 21.680 133.165 22.210 133.530 ;
        RECT 21.680 132.465 21.850 133.165 ;
        RECT 22.380 133.085 22.550 133.700 ;
        RECT 22.720 133.345 22.890 134.145 ;
        RECT 23.060 133.645 23.310 133.975 ;
        RECT 23.535 133.675 24.420 133.845 ;
        RECT 22.380 132.995 22.890 133.085 ;
        RECT 20.930 132.185 21.155 132.315 ;
        RECT 21.325 132.245 21.850 132.465 ;
        RECT 22.020 132.825 22.890 132.995 ;
        RECT 20.565 131.595 20.815 132.055 ;
        RECT 20.985 132.045 21.155 132.185 ;
        RECT 22.020 132.045 22.190 132.825 ;
        RECT 22.720 132.755 22.890 132.825 ;
        RECT 22.400 132.575 22.600 132.605 ;
        RECT 23.060 132.575 23.230 133.645 ;
        RECT 23.400 132.755 23.590 133.475 ;
        RECT 22.400 132.275 23.230 132.575 ;
        RECT 23.760 132.545 24.080 133.505 ;
        RECT 20.985 131.875 21.320 132.045 ;
        RECT 21.515 131.875 22.190 132.045 ;
        RECT 22.510 131.595 22.880 132.095 ;
        RECT 23.060 132.045 23.230 132.275 ;
        RECT 23.615 132.215 24.080 132.545 ;
        RECT 24.250 132.835 24.420 133.675 ;
        RECT 24.600 133.645 24.915 134.145 ;
        RECT 25.145 133.415 25.485 133.975 ;
        RECT 24.590 133.040 25.485 133.415 ;
        RECT 25.655 133.135 25.825 134.145 ;
        RECT 25.295 132.835 25.485 133.040 ;
        RECT 25.995 133.085 26.325 133.930 ;
        RECT 27.015 133.345 27.455 133.975 ;
        RECT 25.995 133.005 26.385 133.085 ;
        RECT 26.170 132.955 26.385 133.005 ;
        RECT 24.250 132.505 25.125 132.835 ;
        RECT 25.295 132.505 26.045 132.835 ;
        RECT 24.250 132.045 24.420 132.505 ;
        RECT 25.295 132.335 25.495 132.505 ;
        RECT 26.215 132.375 26.385 132.955 ;
        RECT 26.160 132.335 26.385 132.375 ;
        RECT 23.060 131.875 23.465 132.045 ;
        RECT 23.635 131.875 24.420 132.045 ;
        RECT 24.695 131.595 24.905 132.125 ;
        RECT 25.165 131.810 25.495 132.335 ;
        RECT 26.005 132.250 26.385 132.335 ;
        RECT 27.015 132.335 27.325 133.345 ;
        RECT 27.630 133.295 27.945 134.145 ;
        RECT 28.115 133.805 29.545 133.975 ;
        RECT 28.115 133.125 28.285 133.805 ;
        RECT 27.495 132.955 28.285 133.125 ;
        RECT 27.495 132.505 27.665 132.955 ;
        RECT 28.455 132.835 28.655 133.635 ;
        RECT 27.835 132.505 28.225 132.785 ;
        RECT 28.410 132.505 28.655 132.835 ;
        RECT 28.855 132.505 29.105 133.635 ;
        RECT 29.295 133.175 29.545 133.805 ;
        RECT 29.725 133.345 30.055 134.145 ;
        RECT 29.295 133.005 30.065 133.175 ;
        RECT 29.320 132.505 29.725 132.835 ;
        RECT 29.895 132.335 30.065 133.005 ;
        RECT 30.235 132.980 30.525 134.145 ;
        RECT 30.730 133.355 31.265 133.975 ;
        RECT 25.665 131.595 25.835 132.205 ;
        RECT 26.005 131.815 26.335 132.250 ;
        RECT 27.015 131.775 27.455 132.335 ;
        RECT 27.625 131.595 28.075 132.335 ;
        RECT 28.245 132.165 29.405 132.335 ;
        RECT 28.245 131.765 28.415 132.165 ;
        RECT 28.585 131.595 29.005 131.995 ;
        RECT 29.175 131.765 29.405 132.165 ;
        RECT 29.575 131.765 30.065 132.335 ;
        RECT 30.730 132.335 31.045 133.355 ;
        RECT 31.435 133.345 31.765 134.145 ;
        RECT 32.250 133.175 32.640 133.350 ;
        RECT 31.215 133.005 32.640 133.175 ;
        RECT 33.055 133.005 33.265 134.145 ;
        RECT 31.215 132.505 31.385 133.005 ;
        RECT 30.235 131.595 30.525 132.320 ;
        RECT 30.730 131.765 31.345 132.335 ;
        RECT 31.635 132.275 31.900 132.835 ;
        RECT 32.070 132.105 32.240 133.005 ;
        RECT 33.435 132.995 33.765 133.975 ;
        RECT 33.935 133.005 34.165 134.145 ;
        RECT 34.375 133.710 39.720 134.145 ;
        RECT 39.895 133.710 45.240 134.145 ;
        RECT 45.415 133.710 50.760 134.145 ;
        RECT 32.410 132.275 32.765 132.835 ;
        RECT 31.515 131.595 31.730 132.105 ;
        RECT 31.960 131.775 32.240 132.105 ;
        RECT 32.420 131.595 32.660 132.105 ;
        RECT 33.055 131.595 33.265 132.415 ;
        RECT 33.435 132.395 33.685 132.995 ;
        RECT 33.855 132.585 34.185 132.835 ;
        RECT 33.435 131.765 33.765 132.395 ;
        RECT 33.935 131.595 34.165 132.415 ;
        RECT 35.960 132.140 36.300 132.970 ;
        RECT 37.780 132.460 38.130 133.710 ;
        RECT 41.480 132.140 41.820 132.970 ;
        RECT 43.300 132.460 43.650 133.710 ;
        RECT 47.000 132.140 47.340 132.970 ;
        RECT 48.820 132.460 49.170 133.710 ;
        RECT 50.935 133.055 54.445 134.145 ;
        RECT 54.615 133.055 55.825 134.145 ;
        RECT 50.935 132.365 52.585 132.885 ;
        RECT 52.755 132.535 54.445 133.055 ;
        RECT 34.375 131.595 39.720 132.140 ;
        RECT 39.895 131.595 45.240 132.140 ;
        RECT 45.415 131.595 50.760 132.140 ;
        RECT 50.935 131.595 54.445 132.365 ;
        RECT 54.615 132.345 55.135 132.885 ;
        RECT 55.305 132.515 55.825 133.055 ;
        RECT 55.995 132.980 56.285 134.145 ;
        RECT 56.455 133.710 61.800 134.145 ;
        RECT 54.615 131.595 55.825 132.345 ;
        RECT 55.995 131.595 56.285 132.320 ;
        RECT 58.040 132.140 58.380 132.970 ;
        RECT 59.860 132.460 60.210 133.710 ;
        RECT 62.065 133.475 62.235 133.975 ;
        RECT 62.405 133.645 62.735 134.145 ;
        RECT 62.065 133.305 62.730 133.475 ;
        RECT 61.980 132.485 62.330 133.135 ;
        RECT 62.500 132.315 62.730 133.305 ;
        RECT 62.065 132.145 62.730 132.315 ;
        RECT 56.455 131.595 61.800 132.140 ;
        RECT 62.065 131.855 62.235 132.145 ;
        RECT 62.405 131.595 62.735 131.975 ;
        RECT 62.905 131.855 63.090 133.975 ;
        RECT 63.330 133.685 63.595 134.145 ;
        RECT 63.765 133.550 64.015 133.975 ;
        RECT 64.225 133.700 65.330 133.870 ;
        RECT 63.710 133.420 64.015 133.550 ;
        RECT 63.260 132.225 63.540 133.175 ;
        RECT 63.710 132.315 63.880 133.420 ;
        RECT 64.050 132.635 64.290 133.230 ;
        RECT 64.460 133.165 64.990 133.530 ;
        RECT 64.460 132.465 64.630 133.165 ;
        RECT 65.160 133.085 65.330 133.700 ;
        RECT 65.500 133.345 65.670 134.145 ;
        RECT 65.840 133.645 66.090 133.975 ;
        RECT 66.315 133.675 67.200 133.845 ;
        RECT 65.160 132.995 65.670 133.085 ;
        RECT 63.710 132.185 63.935 132.315 ;
        RECT 64.105 132.245 64.630 132.465 ;
        RECT 64.800 132.825 65.670 132.995 ;
        RECT 63.345 131.595 63.595 132.055 ;
        RECT 63.765 132.045 63.935 132.185 ;
        RECT 64.800 132.045 64.970 132.825 ;
        RECT 65.500 132.755 65.670 132.825 ;
        RECT 65.180 132.575 65.380 132.605 ;
        RECT 65.840 132.575 66.010 133.645 ;
        RECT 66.180 132.755 66.370 133.475 ;
        RECT 65.180 132.275 66.010 132.575 ;
        RECT 66.540 132.545 66.860 133.505 ;
        RECT 63.765 131.875 64.100 132.045 ;
        RECT 64.295 131.875 64.970 132.045 ;
        RECT 65.290 131.595 65.660 132.095 ;
        RECT 65.840 132.045 66.010 132.275 ;
        RECT 66.395 132.215 66.860 132.545 ;
        RECT 67.030 132.835 67.200 133.675 ;
        RECT 67.380 133.645 67.695 134.145 ;
        RECT 67.925 133.415 68.265 133.975 ;
        RECT 67.370 133.040 68.265 133.415 ;
        RECT 68.435 133.135 68.605 134.145 ;
        RECT 68.075 132.835 68.265 133.040 ;
        RECT 68.775 133.085 69.105 133.930 ;
        RECT 69.275 133.230 69.445 134.145 ;
        RECT 69.795 133.425 70.255 133.975 ;
        RECT 70.445 133.425 70.775 134.145 ;
        RECT 68.775 133.005 69.165 133.085 ;
        RECT 68.950 132.955 69.165 133.005 ;
        RECT 67.030 132.505 67.905 132.835 ;
        RECT 68.075 132.505 68.825 132.835 ;
        RECT 67.030 132.045 67.200 132.505 ;
        RECT 68.075 132.335 68.275 132.505 ;
        RECT 68.995 132.375 69.165 132.955 ;
        RECT 68.940 132.335 69.165 132.375 ;
        RECT 65.840 131.875 66.245 132.045 ;
        RECT 66.415 131.875 67.200 132.045 ;
        RECT 67.475 131.595 67.685 132.125 ;
        RECT 67.945 131.810 68.275 132.335 ;
        RECT 68.785 132.250 69.165 132.335 ;
        RECT 68.445 131.595 68.615 132.205 ;
        RECT 68.785 131.815 69.115 132.250 ;
        RECT 69.285 131.595 69.455 132.110 ;
        RECT 69.795 132.055 70.045 133.425 ;
        RECT 70.975 133.255 71.275 133.805 ;
        RECT 71.445 133.475 71.725 134.145 ;
        RECT 72.645 133.475 72.815 133.975 ;
        RECT 72.985 133.645 73.315 134.145 ;
        RECT 72.645 133.305 73.310 133.475 ;
        RECT 70.335 133.085 71.275 133.255 ;
        RECT 70.335 132.835 70.505 133.085 ;
        RECT 71.645 132.835 71.910 133.195 ;
        RECT 70.215 132.505 70.505 132.835 ;
        RECT 70.675 132.585 71.015 132.835 ;
        RECT 71.235 132.585 71.910 132.835 ;
        RECT 70.335 132.415 70.505 132.505 ;
        RECT 72.560 132.485 72.910 133.135 ;
        RECT 70.335 132.225 71.725 132.415 ;
        RECT 73.080 132.315 73.310 133.305 ;
        RECT 69.795 131.765 70.355 132.055 ;
        RECT 70.525 131.595 70.775 132.055 ;
        RECT 71.395 131.865 71.725 132.225 ;
        RECT 72.645 132.145 73.310 132.315 ;
        RECT 72.645 131.855 72.815 132.145 ;
        RECT 72.985 131.595 73.315 131.975 ;
        RECT 73.485 131.855 73.670 133.975 ;
        RECT 73.910 133.685 74.175 134.145 ;
        RECT 74.345 133.550 74.595 133.975 ;
        RECT 74.805 133.700 75.910 133.870 ;
        RECT 74.290 133.420 74.595 133.550 ;
        RECT 73.840 132.225 74.120 133.175 ;
        RECT 74.290 132.315 74.460 133.420 ;
        RECT 74.630 132.635 74.870 133.230 ;
        RECT 75.040 133.165 75.570 133.530 ;
        RECT 75.040 132.465 75.210 133.165 ;
        RECT 75.740 133.085 75.910 133.700 ;
        RECT 76.080 133.345 76.250 134.145 ;
        RECT 76.420 133.645 76.670 133.975 ;
        RECT 76.895 133.675 77.780 133.845 ;
        RECT 75.740 132.995 76.250 133.085 ;
        RECT 74.290 132.185 74.515 132.315 ;
        RECT 74.685 132.245 75.210 132.465 ;
        RECT 75.380 132.825 76.250 132.995 ;
        RECT 73.925 131.595 74.175 132.055 ;
        RECT 74.345 132.045 74.515 132.185 ;
        RECT 75.380 132.045 75.550 132.825 ;
        RECT 76.080 132.755 76.250 132.825 ;
        RECT 75.760 132.575 75.960 132.605 ;
        RECT 76.420 132.575 76.590 133.645 ;
        RECT 76.760 132.755 76.950 133.475 ;
        RECT 75.760 132.275 76.590 132.575 ;
        RECT 77.120 132.545 77.440 133.505 ;
        RECT 74.345 131.875 74.680 132.045 ;
        RECT 74.875 131.875 75.550 132.045 ;
        RECT 75.870 131.595 76.240 132.095 ;
        RECT 76.420 132.045 76.590 132.275 ;
        RECT 76.975 132.215 77.440 132.545 ;
        RECT 77.610 132.835 77.780 133.675 ;
        RECT 77.960 133.645 78.275 134.145 ;
        RECT 78.505 133.415 78.845 133.975 ;
        RECT 77.950 133.040 78.845 133.415 ;
        RECT 79.015 133.135 79.185 134.145 ;
        RECT 78.655 132.835 78.845 133.040 ;
        RECT 79.355 133.085 79.685 133.930 ;
        RECT 79.355 133.005 79.745 133.085 ;
        RECT 79.915 133.055 81.585 134.145 ;
        RECT 79.530 132.955 79.745 133.005 ;
        RECT 77.610 132.505 78.485 132.835 ;
        RECT 78.655 132.505 79.405 132.835 ;
        RECT 77.610 132.045 77.780 132.505 ;
        RECT 78.655 132.335 78.855 132.505 ;
        RECT 79.575 132.375 79.745 132.955 ;
        RECT 79.520 132.335 79.745 132.375 ;
        RECT 76.420 131.875 76.825 132.045 ;
        RECT 76.995 131.875 77.780 132.045 ;
        RECT 78.055 131.595 78.265 132.125 ;
        RECT 78.525 131.810 78.855 132.335 ;
        RECT 79.365 132.250 79.745 132.335 ;
        RECT 79.915 132.365 80.665 132.885 ;
        RECT 80.835 132.535 81.585 133.055 ;
        RECT 81.755 132.980 82.045 134.145 ;
        RECT 82.215 133.055 83.425 134.145 ;
        RECT 79.025 131.595 79.195 132.205 ;
        RECT 79.365 131.815 79.695 132.250 ;
        RECT 79.915 131.595 81.585 132.365 ;
        RECT 82.215 132.345 82.735 132.885 ;
        RECT 82.905 132.515 83.425 133.055 ;
        RECT 83.595 133.385 84.110 133.795 ;
        RECT 84.345 133.385 84.515 134.145 ;
        RECT 84.685 133.805 86.715 133.975 ;
        RECT 83.595 132.575 83.935 133.385 ;
        RECT 84.685 133.140 84.855 133.805 ;
        RECT 85.250 133.465 86.375 133.635 ;
        RECT 84.105 132.950 84.855 133.140 ;
        RECT 85.025 133.125 86.035 133.295 ;
        RECT 83.595 132.405 84.825 132.575 ;
        RECT 81.755 131.595 82.045 132.320 ;
        RECT 82.215 131.595 83.425 132.345 ;
        RECT 83.870 131.800 84.115 132.405 ;
        RECT 84.335 131.595 84.845 132.130 ;
        RECT 85.025 131.765 85.215 133.125 ;
        RECT 85.385 132.785 85.660 132.925 ;
        RECT 85.385 132.615 85.665 132.785 ;
        RECT 85.385 131.765 85.660 132.615 ;
        RECT 85.865 132.325 86.035 133.125 ;
        RECT 86.205 132.335 86.375 133.465 ;
        RECT 86.545 132.835 86.715 133.805 ;
        RECT 86.885 133.005 87.055 134.145 ;
        RECT 87.225 133.005 87.560 133.975 ;
        RECT 87.825 133.475 87.995 133.975 ;
        RECT 88.165 133.645 88.495 134.145 ;
        RECT 87.825 133.305 88.490 133.475 ;
        RECT 86.545 132.505 86.740 132.835 ;
        RECT 86.965 132.505 87.220 132.835 ;
        RECT 86.965 132.335 87.135 132.505 ;
        RECT 87.390 132.335 87.560 133.005 ;
        RECT 87.740 132.485 88.090 133.135 ;
        RECT 86.205 132.165 87.135 132.335 ;
        RECT 86.205 132.130 86.380 132.165 ;
        RECT 85.850 131.765 86.380 132.130 ;
        RECT 86.805 131.595 87.135 131.995 ;
        RECT 87.305 131.765 87.560 132.335 ;
        RECT 88.260 132.315 88.490 133.305 ;
        RECT 87.825 132.145 88.490 132.315 ;
        RECT 87.825 131.855 87.995 132.145 ;
        RECT 88.165 131.595 88.495 131.975 ;
        RECT 88.665 131.855 88.850 133.975 ;
        RECT 89.090 133.685 89.355 134.145 ;
        RECT 89.525 133.550 89.775 133.975 ;
        RECT 89.985 133.700 91.090 133.870 ;
        RECT 89.470 133.420 89.775 133.550 ;
        RECT 89.020 132.225 89.300 133.175 ;
        RECT 89.470 132.315 89.640 133.420 ;
        RECT 89.810 132.635 90.050 133.230 ;
        RECT 90.220 133.165 90.750 133.530 ;
        RECT 90.220 132.465 90.390 133.165 ;
        RECT 90.920 133.085 91.090 133.700 ;
        RECT 91.260 133.345 91.430 134.145 ;
        RECT 91.600 133.645 91.850 133.975 ;
        RECT 92.075 133.675 92.960 133.845 ;
        RECT 90.920 132.995 91.430 133.085 ;
        RECT 89.470 132.185 89.695 132.315 ;
        RECT 89.865 132.245 90.390 132.465 ;
        RECT 90.560 132.825 91.430 132.995 ;
        RECT 89.105 131.595 89.355 132.055 ;
        RECT 89.525 132.045 89.695 132.185 ;
        RECT 90.560 132.045 90.730 132.825 ;
        RECT 91.260 132.755 91.430 132.825 ;
        RECT 90.940 132.575 91.140 132.605 ;
        RECT 91.600 132.575 91.770 133.645 ;
        RECT 91.940 132.755 92.130 133.475 ;
        RECT 90.940 132.275 91.770 132.575 ;
        RECT 92.300 132.545 92.620 133.505 ;
        RECT 89.525 131.875 89.860 132.045 ;
        RECT 90.055 131.875 90.730 132.045 ;
        RECT 91.050 131.595 91.420 132.095 ;
        RECT 91.600 132.045 91.770 132.275 ;
        RECT 92.155 132.215 92.620 132.545 ;
        RECT 92.790 132.835 92.960 133.675 ;
        RECT 93.140 133.645 93.455 134.145 ;
        RECT 93.685 133.415 94.025 133.975 ;
        RECT 93.130 133.040 94.025 133.415 ;
        RECT 94.195 133.135 94.365 134.145 ;
        RECT 93.835 132.835 94.025 133.040 ;
        RECT 94.535 133.085 94.865 133.930 ;
        RECT 95.035 133.230 95.205 134.145 ;
        RECT 94.535 133.005 94.925 133.085 ;
        RECT 94.710 132.955 94.925 133.005 ;
        RECT 92.790 132.505 93.665 132.835 ;
        RECT 93.835 132.505 94.585 132.835 ;
        RECT 92.790 132.045 92.960 132.505 ;
        RECT 93.835 132.335 94.035 132.505 ;
        RECT 94.755 132.375 94.925 132.955 ;
        RECT 94.700 132.335 94.925 132.375 ;
        RECT 91.600 131.875 92.005 132.045 ;
        RECT 92.175 131.875 92.960 132.045 ;
        RECT 93.235 131.595 93.445 132.125 ;
        RECT 93.705 131.810 94.035 132.335 ;
        RECT 94.545 132.250 94.925 132.335 ;
        RECT 95.555 133.005 95.940 133.975 ;
        RECT 96.110 133.685 96.435 134.145 ;
        RECT 96.955 133.515 97.235 133.975 ;
        RECT 96.110 133.295 97.235 133.515 ;
        RECT 95.555 132.335 95.835 133.005 ;
        RECT 96.110 132.835 96.560 133.295 ;
        RECT 97.425 133.125 97.825 133.975 ;
        RECT 98.225 133.685 98.495 134.145 ;
        RECT 98.665 133.515 98.950 133.975 ;
        RECT 96.005 132.505 96.560 132.835 ;
        RECT 96.730 132.565 97.825 133.125 ;
        RECT 96.110 132.395 96.560 132.505 ;
        RECT 94.205 131.595 94.375 132.205 ;
        RECT 94.545 131.815 94.875 132.250 ;
        RECT 95.045 131.595 95.215 132.110 ;
        RECT 95.555 131.765 95.940 132.335 ;
        RECT 96.110 132.225 97.235 132.395 ;
        RECT 96.110 131.595 96.435 132.055 ;
        RECT 96.955 131.765 97.235 132.225 ;
        RECT 97.425 131.765 97.825 132.565 ;
        RECT 97.995 133.295 98.950 133.515 ;
        RECT 99.810 133.515 100.095 133.975 ;
        RECT 100.265 133.685 100.535 134.145 ;
        RECT 99.810 133.295 100.765 133.515 ;
        RECT 97.995 132.395 98.205 133.295 ;
        RECT 98.375 132.565 99.065 133.125 ;
        RECT 99.695 132.565 100.385 133.125 ;
        RECT 100.555 132.395 100.765 133.295 ;
        RECT 97.995 132.225 98.950 132.395 ;
        RECT 98.225 131.595 98.495 132.055 ;
        RECT 98.665 131.765 98.950 132.225 ;
        RECT 99.810 132.225 100.765 132.395 ;
        RECT 100.935 133.125 101.335 133.975 ;
        RECT 101.525 133.515 101.805 133.975 ;
        RECT 102.325 133.685 102.650 134.145 ;
        RECT 101.525 133.295 102.650 133.515 ;
        RECT 100.935 132.565 102.030 133.125 ;
        RECT 102.200 132.835 102.650 133.295 ;
        RECT 102.820 133.005 103.205 133.975 ;
        RECT 99.810 131.765 100.095 132.225 ;
        RECT 100.265 131.595 100.535 132.055 ;
        RECT 100.935 131.765 101.335 132.565 ;
        RECT 102.200 132.505 102.755 132.835 ;
        RECT 102.200 132.395 102.650 132.505 ;
        RECT 101.525 132.225 102.650 132.395 ;
        RECT 102.925 132.335 103.205 133.005 ;
        RECT 103.375 133.385 103.890 133.795 ;
        RECT 104.125 133.385 104.295 134.145 ;
        RECT 104.465 133.805 106.495 133.975 ;
        RECT 103.375 132.575 103.715 133.385 ;
        RECT 104.465 133.140 104.635 133.805 ;
        RECT 105.030 133.465 106.155 133.635 ;
        RECT 103.885 132.950 104.635 133.140 ;
        RECT 104.805 133.125 105.815 133.295 ;
        RECT 103.375 132.405 104.605 132.575 ;
        RECT 101.525 131.765 101.805 132.225 ;
        RECT 102.325 131.595 102.650 132.055 ;
        RECT 102.820 131.765 103.205 132.335 ;
        RECT 103.650 131.800 103.895 132.405 ;
        RECT 104.115 131.595 104.625 132.130 ;
        RECT 104.805 131.765 104.995 133.125 ;
        RECT 105.165 132.445 105.440 132.925 ;
        RECT 105.165 132.275 105.445 132.445 ;
        RECT 105.645 132.325 105.815 133.125 ;
        RECT 105.985 132.335 106.155 133.465 ;
        RECT 106.325 132.835 106.495 133.805 ;
        RECT 106.665 133.005 106.835 134.145 ;
        RECT 107.005 133.005 107.340 133.975 ;
        RECT 106.325 132.505 106.520 132.835 ;
        RECT 106.745 132.505 107.000 132.835 ;
        RECT 106.745 132.335 106.915 132.505 ;
        RECT 107.170 132.335 107.340 133.005 ;
        RECT 107.515 132.980 107.805 134.145 ;
        RECT 108.065 133.475 108.235 133.975 ;
        RECT 108.405 133.645 108.735 134.145 ;
        RECT 108.065 133.305 108.730 133.475 ;
        RECT 107.980 132.485 108.330 133.135 ;
        RECT 105.165 131.765 105.440 132.275 ;
        RECT 105.985 132.165 106.915 132.335 ;
        RECT 105.985 132.130 106.160 132.165 ;
        RECT 105.630 131.765 106.160 132.130 ;
        RECT 106.585 131.595 106.915 131.995 ;
        RECT 107.085 131.765 107.340 132.335 ;
        RECT 107.515 131.595 107.805 132.320 ;
        RECT 108.500 132.315 108.730 133.305 ;
        RECT 108.065 132.145 108.730 132.315 ;
        RECT 108.065 131.855 108.235 132.145 ;
        RECT 108.405 131.595 108.735 131.975 ;
        RECT 108.905 131.855 109.090 133.975 ;
        RECT 109.330 133.685 109.595 134.145 ;
        RECT 109.765 133.550 110.015 133.975 ;
        RECT 110.225 133.700 111.330 133.870 ;
        RECT 109.710 133.420 110.015 133.550 ;
        RECT 109.260 132.225 109.540 133.175 ;
        RECT 109.710 132.315 109.880 133.420 ;
        RECT 110.050 132.635 110.290 133.230 ;
        RECT 110.460 133.165 110.990 133.530 ;
        RECT 110.460 132.465 110.630 133.165 ;
        RECT 111.160 133.085 111.330 133.700 ;
        RECT 111.500 133.345 111.670 134.145 ;
        RECT 111.840 133.645 112.090 133.975 ;
        RECT 112.315 133.675 113.200 133.845 ;
        RECT 111.160 132.995 111.670 133.085 ;
        RECT 109.710 132.185 109.935 132.315 ;
        RECT 110.105 132.245 110.630 132.465 ;
        RECT 110.800 132.825 111.670 132.995 ;
        RECT 109.345 131.595 109.595 132.055 ;
        RECT 109.765 132.045 109.935 132.185 ;
        RECT 110.800 132.045 110.970 132.825 ;
        RECT 111.500 132.755 111.670 132.825 ;
        RECT 111.180 132.575 111.380 132.605 ;
        RECT 111.840 132.575 112.010 133.645 ;
        RECT 112.180 132.755 112.370 133.475 ;
        RECT 111.180 132.275 112.010 132.575 ;
        RECT 112.540 132.545 112.860 133.505 ;
        RECT 109.765 131.875 110.100 132.045 ;
        RECT 110.295 131.875 110.970 132.045 ;
        RECT 111.290 131.595 111.660 132.095 ;
        RECT 111.840 132.045 112.010 132.275 ;
        RECT 112.395 132.215 112.860 132.545 ;
        RECT 113.030 132.835 113.200 133.675 ;
        RECT 113.380 133.645 113.695 134.145 ;
        RECT 113.925 133.415 114.265 133.975 ;
        RECT 113.370 133.040 114.265 133.415 ;
        RECT 114.435 133.135 114.605 134.145 ;
        RECT 114.075 132.835 114.265 133.040 ;
        RECT 114.775 133.085 115.105 133.930 ;
        RECT 115.335 133.710 120.680 134.145 ;
        RECT 114.775 133.005 115.165 133.085 ;
        RECT 114.950 132.955 115.165 133.005 ;
        RECT 113.030 132.505 113.905 132.835 ;
        RECT 114.075 132.505 114.825 132.835 ;
        RECT 113.030 132.045 113.200 132.505 ;
        RECT 114.075 132.335 114.275 132.505 ;
        RECT 114.995 132.375 115.165 132.955 ;
        RECT 114.940 132.335 115.165 132.375 ;
        RECT 111.840 131.875 112.245 132.045 ;
        RECT 112.415 131.875 113.200 132.045 ;
        RECT 113.475 131.595 113.685 132.125 ;
        RECT 113.945 131.810 114.275 132.335 ;
        RECT 114.785 132.250 115.165 132.335 ;
        RECT 114.445 131.595 114.615 132.205 ;
        RECT 114.785 131.815 115.115 132.250 ;
        RECT 116.920 132.140 117.260 132.970 ;
        RECT 118.740 132.460 119.090 133.710 ;
        RECT 120.855 132.540 121.135 133.975 ;
        RECT 121.305 133.370 122.015 134.145 ;
        RECT 122.185 133.200 122.515 133.975 ;
        RECT 121.365 132.985 122.515 133.200 ;
        RECT 115.335 131.595 120.680 132.140 ;
        RECT 120.855 131.765 121.195 132.540 ;
        RECT 121.365 132.415 121.650 132.985 ;
        RECT 121.835 132.585 122.305 132.815 ;
        RECT 122.710 132.785 122.925 133.900 ;
        RECT 123.105 133.425 123.435 134.145 ;
        RECT 123.615 133.710 128.960 134.145 ;
        RECT 123.215 132.785 123.445 133.125 ;
        RECT 122.475 132.605 122.925 132.785 ;
        RECT 122.475 132.585 122.805 132.605 ;
        RECT 123.115 132.585 123.445 132.785 ;
        RECT 121.365 132.225 122.075 132.415 ;
        RECT 121.775 132.085 122.075 132.225 ;
        RECT 122.265 132.225 123.445 132.415 ;
        RECT 122.265 132.145 122.595 132.225 ;
        RECT 121.775 132.075 122.090 132.085 ;
        RECT 121.775 132.065 122.100 132.075 ;
        RECT 121.775 132.060 122.110 132.065 ;
        RECT 121.365 131.595 121.535 132.055 ;
        RECT 121.775 132.050 122.115 132.060 ;
        RECT 121.775 132.045 122.120 132.050 ;
        RECT 121.775 132.035 122.125 132.045 ;
        RECT 121.775 132.030 122.130 132.035 ;
        RECT 121.775 131.765 122.135 132.030 ;
        RECT 122.765 131.595 122.935 132.055 ;
        RECT 123.105 131.765 123.445 132.225 ;
        RECT 125.200 132.140 125.540 132.970 ;
        RECT 127.020 132.460 127.370 133.710 ;
        RECT 129.135 133.055 132.645 134.145 ;
        RECT 129.135 132.365 130.785 132.885 ;
        RECT 130.955 132.535 132.645 133.055 ;
        RECT 133.275 132.980 133.565 134.145 ;
        RECT 133.825 133.525 133.995 133.955 ;
        RECT 134.165 133.695 134.495 134.145 ;
        RECT 133.825 133.295 134.500 133.525 ;
        RECT 123.615 131.595 128.960 132.140 ;
        RECT 129.135 131.595 132.645 132.365 ;
        RECT 133.275 131.595 133.565 132.320 ;
        RECT 133.795 132.275 134.095 133.125 ;
        RECT 134.265 132.645 134.500 133.295 ;
        RECT 134.670 132.985 134.955 133.930 ;
        RECT 135.135 133.675 135.820 134.145 ;
        RECT 135.130 133.155 135.825 133.465 ;
        RECT 136.000 133.090 136.305 133.875 ;
        RECT 136.495 133.710 141.840 134.145 ;
        RECT 134.670 132.835 135.530 132.985 ;
        RECT 134.670 132.815 135.955 132.835 ;
        RECT 134.265 132.315 134.800 132.645 ;
        RECT 134.970 132.455 135.955 132.815 ;
        RECT 134.265 132.165 134.485 132.315 ;
        RECT 133.740 131.595 134.075 132.100 ;
        RECT 134.245 131.790 134.485 132.165 ;
        RECT 134.970 132.120 135.140 132.455 ;
        RECT 136.130 132.285 136.305 133.090 ;
        RECT 134.765 131.925 135.140 132.120 ;
        RECT 134.765 131.780 134.935 131.925 ;
        RECT 135.500 131.595 135.895 132.090 ;
        RECT 136.065 131.765 136.305 132.285 ;
        RECT 138.080 132.140 138.420 132.970 ;
        RECT 139.900 132.460 140.250 133.710 ;
        RECT 142.105 133.215 142.275 133.975 ;
        RECT 142.490 133.385 142.820 134.145 ;
        RECT 142.105 133.045 142.820 133.215 ;
        RECT 142.990 133.070 143.245 133.975 ;
        RECT 142.015 132.495 142.370 132.865 ;
        RECT 142.650 132.835 142.820 133.045 ;
        RECT 142.650 132.505 142.905 132.835 ;
        RECT 142.650 132.315 142.820 132.505 ;
        RECT 143.075 132.340 143.245 133.070 ;
        RECT 143.420 132.995 143.680 134.145 ;
        RECT 143.945 133.215 144.115 133.975 ;
        RECT 144.330 133.385 144.660 134.145 ;
        RECT 143.945 133.045 144.660 133.215 ;
        RECT 144.830 133.070 145.085 133.975 ;
        RECT 143.855 132.495 144.210 132.865 ;
        RECT 144.490 132.835 144.660 133.045 ;
        RECT 144.490 132.505 144.745 132.835 ;
        RECT 142.105 132.145 142.820 132.315 ;
        RECT 136.495 131.595 141.840 132.140 ;
        RECT 142.105 131.765 142.275 132.145 ;
        RECT 142.490 131.595 142.820 131.975 ;
        RECT 142.990 131.765 143.245 132.340 ;
        RECT 143.420 131.595 143.680 132.435 ;
        RECT 144.490 132.315 144.660 132.505 ;
        RECT 144.915 132.340 145.085 133.070 ;
        RECT 145.260 132.995 145.520 134.145 ;
        RECT 145.695 133.055 146.905 134.145 ;
        RECT 145.695 132.515 146.215 133.055 ;
        RECT 143.945 132.145 144.660 132.315 ;
        RECT 143.945 131.765 144.115 132.145 ;
        RECT 144.330 131.595 144.660 131.975 ;
        RECT 144.830 131.765 145.085 132.340 ;
        RECT 145.260 131.595 145.520 132.435 ;
        RECT 146.385 132.345 146.905 132.885 ;
        RECT 145.695 131.595 146.905 132.345 ;
        RECT 17.270 131.425 146.990 131.595 ;
        RECT 17.355 130.675 18.565 131.425 ;
        RECT 17.355 130.135 17.875 130.675 ;
        RECT 18.740 130.585 19.000 131.425 ;
        RECT 19.175 130.680 19.430 131.255 ;
        RECT 19.600 131.045 19.930 131.425 ;
        RECT 20.145 130.875 20.315 131.255 ;
        RECT 19.600 130.705 20.315 130.875 ;
        RECT 18.045 129.965 18.565 130.505 ;
        RECT 17.355 128.875 18.565 129.965 ;
        RECT 18.740 128.875 19.000 130.025 ;
        RECT 19.175 129.950 19.345 130.680 ;
        RECT 19.600 130.515 19.770 130.705 ;
        RECT 20.575 130.675 21.785 131.425 ;
        RECT 21.960 130.685 22.215 131.255 ;
        RECT 22.385 131.025 22.715 131.425 ;
        RECT 23.140 130.890 23.670 131.255 ;
        RECT 23.140 130.855 23.315 130.890 ;
        RECT 22.385 130.685 23.315 130.855 ;
        RECT 23.860 130.745 24.135 131.255 ;
        RECT 19.515 130.185 19.770 130.515 ;
        RECT 19.600 129.975 19.770 130.185 ;
        RECT 20.050 130.155 20.405 130.525 ;
        RECT 20.575 130.135 21.095 130.675 ;
        RECT 19.175 129.045 19.430 129.950 ;
        RECT 19.600 129.805 20.315 129.975 ;
        RECT 21.265 129.965 21.785 130.505 ;
        RECT 19.600 128.875 19.930 129.635 ;
        RECT 20.145 129.045 20.315 129.805 ;
        RECT 20.575 128.875 21.785 129.965 ;
        RECT 21.960 130.015 22.130 130.685 ;
        RECT 22.385 130.515 22.555 130.685 ;
        RECT 22.300 130.185 22.555 130.515 ;
        RECT 22.780 130.185 22.975 130.515 ;
        RECT 21.960 129.045 22.295 130.015 ;
        RECT 22.465 128.875 22.635 130.015 ;
        RECT 22.805 129.215 22.975 130.185 ;
        RECT 23.145 129.555 23.315 130.685 ;
        RECT 23.485 129.895 23.655 130.695 ;
        RECT 23.855 130.575 24.135 130.745 ;
        RECT 23.860 130.095 24.135 130.575 ;
        RECT 24.305 129.895 24.495 131.255 ;
        RECT 24.675 130.890 25.185 131.425 ;
        RECT 25.405 130.615 25.650 131.220 ;
        RECT 26.095 130.880 31.440 131.425 ;
        RECT 31.615 130.880 36.960 131.425 ;
        RECT 37.135 130.880 42.480 131.425 ;
        RECT 24.695 130.445 25.925 130.615 ;
        RECT 23.485 129.725 24.495 129.895 ;
        RECT 24.665 129.880 25.415 130.070 ;
        RECT 23.145 129.385 24.270 129.555 ;
        RECT 24.665 129.215 24.835 129.880 ;
        RECT 25.585 129.635 25.925 130.445 ;
        RECT 27.680 130.050 28.020 130.880 ;
        RECT 22.805 129.045 24.835 129.215 ;
        RECT 25.005 128.875 25.175 129.635 ;
        RECT 25.410 129.225 25.925 129.635 ;
        RECT 29.500 129.310 29.850 130.560 ;
        RECT 33.200 130.050 33.540 130.880 ;
        RECT 35.020 129.310 35.370 130.560 ;
        RECT 38.720 130.050 39.060 130.880 ;
        RECT 43.115 130.700 43.405 131.425 ;
        RECT 43.575 130.880 48.920 131.425 ;
        RECT 49.095 130.880 54.440 131.425 ;
        RECT 54.615 130.880 59.960 131.425 ;
        RECT 60.640 130.965 60.905 131.425 ;
        RECT 40.540 129.310 40.890 130.560 ;
        RECT 45.160 130.050 45.500 130.880 ;
        RECT 26.095 128.875 31.440 129.310 ;
        RECT 31.615 128.875 36.960 129.310 ;
        RECT 37.135 128.875 42.480 129.310 ;
        RECT 43.115 128.875 43.405 130.040 ;
        RECT 46.980 129.310 47.330 130.560 ;
        RECT 50.680 130.050 51.020 130.880 ;
        RECT 52.500 129.310 52.850 130.560 ;
        RECT 56.200 130.050 56.540 130.880 ;
        RECT 61.275 130.785 61.445 131.255 ;
        RECT 61.695 130.965 61.865 131.425 ;
        RECT 62.115 130.785 62.285 131.255 ;
        RECT 62.535 130.965 62.705 131.425 ;
        RECT 62.955 130.785 63.125 131.255 ;
        RECT 63.295 130.960 63.545 131.425 ;
        RECT 63.875 130.965 64.120 131.425 ;
        RECT 61.275 130.605 63.645 130.785 ;
        RECT 58.020 129.310 58.370 130.560 ;
        RECT 60.615 130.185 63.125 130.435 ;
        RECT 63.295 130.015 63.645 130.605 ;
        RECT 63.815 130.185 64.130 130.795 ;
        RECT 64.300 130.435 64.550 131.245 ;
        RECT 64.720 130.900 64.980 131.425 ;
        RECT 65.150 130.775 65.410 131.230 ;
        RECT 65.580 130.945 65.840 131.425 ;
        RECT 66.010 130.775 66.270 131.230 ;
        RECT 66.440 130.945 66.700 131.425 ;
        RECT 66.870 130.775 67.130 131.230 ;
        RECT 67.300 130.945 67.560 131.425 ;
        RECT 67.730 130.775 67.990 131.230 ;
        RECT 68.160 130.945 68.460 131.425 ;
        RECT 65.150 130.605 68.460 130.775 ;
        RECT 68.875 130.700 69.165 131.425 ;
        RECT 69.425 130.875 69.595 131.165 ;
        RECT 69.765 131.045 70.095 131.425 ;
        RECT 69.425 130.705 70.090 130.875 ;
        RECT 64.300 130.185 67.320 130.435 ;
        RECT 43.575 128.875 48.920 129.310 ;
        RECT 49.095 128.875 54.440 129.310 ;
        RECT 54.615 128.875 59.960 129.310 ;
        RECT 60.640 128.875 60.935 130.015 ;
        RECT 61.195 129.845 63.645 130.015 ;
        RECT 61.195 129.045 61.525 129.845 ;
        RECT 61.695 128.875 61.865 129.675 ;
        RECT 62.035 129.045 62.365 129.845 ;
        RECT 62.875 129.825 63.645 129.845 ;
        RECT 62.535 128.875 62.705 129.675 ;
        RECT 62.875 129.045 63.205 129.825 ;
        RECT 63.375 128.875 63.545 129.335 ;
        RECT 63.825 128.875 64.120 129.985 ;
        RECT 64.300 129.050 64.550 130.185 ;
        RECT 67.490 130.015 68.460 130.605 ;
        RECT 64.720 128.875 64.980 129.985 ;
        RECT 65.150 129.775 68.460 130.015 ;
        RECT 65.150 129.050 65.410 129.775 ;
        RECT 65.580 128.875 65.840 129.605 ;
        RECT 66.010 129.050 66.270 129.775 ;
        RECT 66.440 128.875 66.700 129.605 ;
        RECT 66.870 129.050 67.130 129.775 ;
        RECT 67.300 128.875 67.560 129.605 ;
        RECT 67.730 129.050 67.990 129.775 ;
        RECT 68.160 128.875 68.455 129.605 ;
        RECT 68.875 128.875 69.165 130.040 ;
        RECT 69.340 129.885 69.690 130.535 ;
        RECT 69.860 129.715 70.090 130.705 ;
        RECT 69.425 129.545 70.090 129.715 ;
        RECT 69.425 129.045 69.595 129.545 ;
        RECT 69.765 128.875 70.095 129.375 ;
        RECT 70.265 129.045 70.450 131.165 ;
        RECT 70.705 130.965 70.955 131.425 ;
        RECT 71.125 130.975 71.460 131.145 ;
        RECT 71.655 130.975 72.330 131.145 ;
        RECT 71.125 130.835 71.295 130.975 ;
        RECT 70.620 129.845 70.900 130.795 ;
        RECT 71.070 130.705 71.295 130.835 ;
        RECT 71.070 129.600 71.240 130.705 ;
        RECT 71.465 130.555 71.990 130.775 ;
        RECT 71.410 129.790 71.650 130.385 ;
        RECT 71.820 129.855 71.990 130.555 ;
        RECT 72.160 130.195 72.330 130.975 ;
        RECT 72.650 130.925 73.020 131.425 ;
        RECT 73.200 130.975 73.605 131.145 ;
        RECT 73.775 130.975 74.560 131.145 ;
        RECT 73.200 130.745 73.370 130.975 ;
        RECT 72.540 130.445 73.370 130.745 ;
        RECT 73.755 130.475 74.220 130.805 ;
        RECT 72.540 130.415 72.740 130.445 ;
        RECT 72.860 130.195 73.030 130.265 ;
        RECT 72.160 130.025 73.030 130.195 ;
        RECT 72.520 129.935 73.030 130.025 ;
        RECT 71.070 129.470 71.375 129.600 ;
        RECT 71.820 129.490 72.350 129.855 ;
        RECT 70.690 128.875 70.955 129.335 ;
        RECT 71.125 129.045 71.375 129.470 ;
        RECT 72.520 129.320 72.690 129.935 ;
        RECT 71.585 129.150 72.690 129.320 ;
        RECT 72.860 128.875 73.030 129.675 ;
        RECT 73.200 129.375 73.370 130.445 ;
        RECT 73.540 129.545 73.730 130.265 ;
        RECT 73.900 129.515 74.220 130.475 ;
        RECT 74.390 130.515 74.560 130.975 ;
        RECT 74.835 130.895 75.045 131.425 ;
        RECT 75.305 130.685 75.635 131.210 ;
        RECT 75.805 130.815 75.975 131.425 ;
        RECT 76.145 130.770 76.475 131.205 ;
        RECT 76.645 130.910 76.815 131.425 ;
        RECT 77.205 130.770 77.535 131.205 ;
        RECT 77.705 130.815 77.875 131.425 ;
        RECT 76.145 130.685 76.525 130.770 ;
        RECT 75.435 130.515 75.635 130.685 ;
        RECT 76.300 130.645 76.525 130.685 ;
        RECT 74.390 130.185 75.265 130.515 ;
        RECT 75.435 130.185 76.185 130.515 ;
        RECT 73.200 129.045 73.450 129.375 ;
        RECT 74.390 129.345 74.560 130.185 ;
        RECT 75.435 129.980 75.625 130.185 ;
        RECT 76.355 130.065 76.525 130.645 ;
        RECT 76.310 130.015 76.525 130.065 ;
        RECT 74.730 129.605 75.625 129.980 ;
        RECT 76.135 129.935 76.525 130.015 ;
        RECT 77.155 130.685 77.535 130.770 ;
        RECT 78.045 130.685 78.375 131.210 ;
        RECT 78.635 130.895 78.845 131.425 ;
        RECT 79.120 130.975 79.905 131.145 ;
        RECT 80.075 130.975 80.480 131.145 ;
        RECT 77.155 130.645 77.380 130.685 ;
        RECT 77.155 130.065 77.325 130.645 ;
        RECT 78.045 130.515 78.245 130.685 ;
        RECT 79.120 130.515 79.290 130.975 ;
        RECT 77.495 130.185 78.245 130.515 ;
        RECT 78.415 130.185 79.290 130.515 ;
        RECT 77.155 130.015 77.370 130.065 ;
        RECT 77.155 129.935 77.545 130.015 ;
        RECT 73.675 129.175 74.560 129.345 ;
        RECT 74.740 128.875 75.055 129.375 ;
        RECT 75.285 129.045 75.625 129.605 ;
        RECT 75.795 128.875 75.965 129.885 ;
        RECT 76.135 129.090 76.465 129.935 ;
        RECT 76.635 128.875 76.805 129.790 ;
        RECT 77.215 129.090 77.545 129.935 ;
        RECT 78.055 129.980 78.245 130.185 ;
        RECT 77.715 128.875 77.885 129.885 ;
        RECT 78.055 129.605 78.950 129.980 ;
        RECT 78.055 129.045 78.395 129.605 ;
        RECT 78.625 128.875 78.940 129.375 ;
        RECT 79.120 129.345 79.290 130.185 ;
        RECT 79.460 130.475 79.925 130.805 ;
        RECT 80.310 130.745 80.480 130.975 ;
        RECT 80.660 130.925 81.030 131.425 ;
        RECT 81.350 130.975 82.025 131.145 ;
        RECT 82.220 130.975 82.555 131.145 ;
        RECT 79.460 129.515 79.780 130.475 ;
        RECT 80.310 130.445 81.140 130.745 ;
        RECT 79.950 129.545 80.140 130.265 ;
        RECT 80.310 129.375 80.480 130.445 ;
        RECT 80.940 130.415 81.140 130.445 ;
        RECT 80.650 130.195 80.820 130.265 ;
        RECT 81.350 130.195 81.520 130.975 ;
        RECT 82.385 130.835 82.555 130.975 ;
        RECT 82.725 130.965 82.975 131.425 ;
        RECT 80.650 130.025 81.520 130.195 ;
        RECT 81.690 130.555 82.215 130.775 ;
        RECT 82.385 130.705 82.610 130.835 ;
        RECT 80.650 129.935 81.160 130.025 ;
        RECT 79.120 129.175 80.005 129.345 ;
        RECT 80.230 129.045 80.480 129.375 ;
        RECT 80.650 128.875 80.820 129.675 ;
        RECT 80.990 129.320 81.160 129.935 ;
        RECT 81.690 129.855 81.860 130.555 ;
        RECT 81.330 129.490 81.860 129.855 ;
        RECT 82.030 129.790 82.270 130.385 ;
        RECT 82.440 129.600 82.610 130.705 ;
        RECT 82.780 129.845 83.060 130.795 ;
        RECT 82.305 129.470 82.610 129.600 ;
        RECT 80.990 129.150 82.095 129.320 ;
        RECT 82.305 129.045 82.555 129.470 ;
        RECT 82.725 128.875 82.990 129.335 ;
        RECT 83.230 129.045 83.415 131.165 ;
        RECT 83.585 131.045 83.915 131.425 ;
        RECT 84.085 130.875 84.255 131.165 ;
        RECT 83.590 130.705 84.255 130.875 ;
        RECT 85.525 130.875 85.695 131.165 ;
        RECT 85.865 131.045 86.195 131.425 ;
        RECT 85.525 130.705 86.190 130.875 ;
        RECT 83.590 129.715 83.820 130.705 ;
        RECT 83.990 129.885 84.340 130.535 ;
        RECT 85.440 129.885 85.790 130.535 ;
        RECT 85.960 129.715 86.190 130.705 ;
        RECT 83.590 129.545 84.255 129.715 ;
        RECT 83.585 128.875 83.915 129.375 ;
        RECT 84.085 129.045 84.255 129.545 ;
        RECT 85.525 129.545 86.190 129.715 ;
        RECT 85.525 129.045 85.695 129.545 ;
        RECT 85.865 128.875 86.195 129.375 ;
        RECT 86.365 129.045 86.550 131.165 ;
        RECT 86.805 130.965 87.055 131.425 ;
        RECT 87.225 130.975 87.560 131.145 ;
        RECT 87.755 130.975 88.430 131.145 ;
        RECT 87.225 130.835 87.395 130.975 ;
        RECT 86.720 129.845 87.000 130.795 ;
        RECT 87.170 130.705 87.395 130.835 ;
        RECT 87.170 129.600 87.340 130.705 ;
        RECT 87.565 130.555 88.090 130.775 ;
        RECT 87.510 129.790 87.750 130.385 ;
        RECT 87.920 129.855 88.090 130.555 ;
        RECT 88.260 130.195 88.430 130.975 ;
        RECT 88.750 130.925 89.120 131.425 ;
        RECT 89.300 130.975 89.705 131.145 ;
        RECT 89.875 130.975 90.660 131.145 ;
        RECT 89.300 130.745 89.470 130.975 ;
        RECT 88.640 130.445 89.470 130.745 ;
        RECT 89.855 130.475 90.320 130.805 ;
        RECT 88.640 130.415 88.840 130.445 ;
        RECT 88.960 130.195 89.130 130.265 ;
        RECT 88.260 130.025 89.130 130.195 ;
        RECT 88.620 129.935 89.130 130.025 ;
        RECT 87.170 129.470 87.475 129.600 ;
        RECT 87.920 129.490 88.450 129.855 ;
        RECT 86.790 128.875 87.055 129.335 ;
        RECT 87.225 129.045 87.475 129.470 ;
        RECT 88.620 129.320 88.790 129.935 ;
        RECT 87.685 129.150 88.790 129.320 ;
        RECT 88.960 128.875 89.130 129.675 ;
        RECT 89.300 129.375 89.470 130.445 ;
        RECT 89.640 129.545 89.830 130.265 ;
        RECT 90.000 129.515 90.320 130.475 ;
        RECT 90.490 130.515 90.660 130.975 ;
        RECT 90.935 130.895 91.145 131.425 ;
        RECT 91.405 130.685 91.735 131.210 ;
        RECT 91.905 130.815 92.075 131.425 ;
        RECT 92.245 130.770 92.575 131.205 ;
        RECT 92.745 130.910 92.915 131.425 ;
        RECT 92.245 130.685 92.625 130.770 ;
        RECT 91.535 130.515 91.735 130.685 ;
        RECT 92.400 130.645 92.625 130.685 ;
        RECT 90.490 130.185 91.365 130.515 ;
        RECT 91.535 130.185 92.285 130.515 ;
        RECT 89.300 129.045 89.550 129.375 ;
        RECT 90.490 129.345 90.660 130.185 ;
        RECT 91.535 129.980 91.725 130.185 ;
        RECT 92.455 130.065 92.625 130.645 ;
        RECT 93.255 130.675 94.465 131.425 ;
        RECT 94.635 130.700 94.925 131.425 ;
        RECT 93.255 130.135 93.775 130.675 ;
        RECT 95.095 130.655 97.685 131.425 ;
        RECT 97.970 130.795 98.255 131.255 ;
        RECT 98.425 130.965 98.695 131.425 ;
        RECT 92.410 130.015 92.625 130.065 ;
        RECT 90.830 129.605 91.725 129.980 ;
        RECT 92.235 129.935 92.625 130.015 ;
        RECT 93.945 129.965 94.465 130.505 ;
        RECT 95.095 130.135 96.305 130.655 ;
        RECT 97.970 130.625 98.925 130.795 ;
        RECT 89.775 129.175 90.660 129.345 ;
        RECT 90.840 128.875 91.155 129.375 ;
        RECT 91.385 129.045 91.725 129.605 ;
        RECT 91.895 128.875 92.065 129.885 ;
        RECT 92.235 129.090 92.565 129.935 ;
        RECT 92.735 128.875 92.905 129.790 ;
        RECT 93.255 128.875 94.465 129.965 ;
        RECT 94.635 128.875 94.925 130.040 ;
        RECT 96.475 129.965 97.685 130.485 ;
        RECT 95.095 128.875 97.685 129.965 ;
        RECT 97.855 129.895 98.545 130.455 ;
        RECT 98.715 129.725 98.925 130.625 ;
        RECT 97.970 129.505 98.925 129.725 ;
        RECT 99.095 130.455 99.495 131.255 ;
        RECT 99.685 130.795 99.965 131.255 ;
        RECT 100.485 130.965 100.810 131.425 ;
        RECT 99.685 130.625 100.810 130.795 ;
        RECT 100.980 130.685 101.365 131.255 ;
        RECT 100.360 130.515 100.810 130.625 ;
        RECT 99.095 129.895 100.190 130.455 ;
        RECT 100.360 130.185 100.915 130.515 ;
        RECT 97.970 129.045 98.255 129.505 ;
        RECT 98.425 128.875 98.695 129.335 ;
        RECT 99.095 129.045 99.495 129.895 ;
        RECT 100.360 129.725 100.810 130.185 ;
        RECT 101.085 130.015 101.365 130.685 ;
        RECT 101.535 130.655 105.045 131.425 ;
        RECT 105.215 130.675 106.425 131.425 ;
        RECT 106.645 130.885 106.870 131.245 ;
        RECT 107.050 131.055 107.380 131.425 ;
        RECT 107.560 130.885 107.815 131.245 ;
        RECT 108.380 131.055 109.125 131.425 ;
        RECT 106.645 130.695 109.130 130.885 ;
        RECT 101.535 130.135 103.185 130.655 ;
        RECT 99.685 129.505 100.810 129.725 ;
        RECT 99.685 129.045 99.965 129.505 ;
        RECT 100.485 128.875 100.810 129.335 ;
        RECT 100.980 129.045 101.365 130.015 ;
        RECT 103.355 129.965 105.045 130.485 ;
        RECT 105.215 130.135 105.735 130.675 ;
        RECT 105.905 129.965 106.425 130.505 ;
        RECT 106.605 130.185 106.875 130.515 ;
        RECT 107.055 130.185 107.490 130.515 ;
        RECT 107.670 130.185 108.245 130.515 ;
        RECT 108.425 130.185 108.705 130.515 ;
        RECT 108.905 130.005 109.130 130.695 ;
        RECT 101.535 128.875 105.045 129.965 ;
        RECT 105.215 128.875 106.425 129.965 ;
        RECT 106.635 129.825 109.130 130.005 ;
        RECT 109.305 129.825 109.640 131.245 ;
        RECT 109.815 130.655 111.485 131.425 ;
        RECT 111.745 130.875 111.915 131.165 ;
        RECT 112.085 131.045 112.415 131.425 ;
        RECT 111.745 130.705 112.410 130.875 ;
        RECT 109.815 130.135 110.565 130.655 ;
        RECT 110.735 129.965 111.485 130.485 ;
        RECT 106.635 129.055 106.925 129.825 ;
        RECT 107.495 129.415 108.685 129.645 ;
        RECT 107.495 129.055 107.755 129.415 ;
        RECT 107.925 128.875 108.255 129.245 ;
        RECT 108.425 129.055 108.685 129.415 ;
        RECT 108.875 128.875 109.205 129.595 ;
        RECT 109.375 129.055 109.640 129.825 ;
        RECT 109.815 128.875 111.485 129.965 ;
        RECT 111.660 129.885 112.010 130.535 ;
        RECT 112.180 129.715 112.410 130.705 ;
        RECT 111.745 129.545 112.410 129.715 ;
        RECT 111.745 129.045 111.915 129.545 ;
        RECT 112.085 128.875 112.415 129.375 ;
        RECT 112.585 129.045 112.770 131.165 ;
        RECT 113.025 130.965 113.275 131.425 ;
        RECT 113.445 130.975 113.780 131.145 ;
        RECT 113.975 130.975 114.650 131.145 ;
        RECT 113.445 130.835 113.615 130.975 ;
        RECT 112.940 129.845 113.220 130.795 ;
        RECT 113.390 130.705 113.615 130.835 ;
        RECT 113.390 129.600 113.560 130.705 ;
        RECT 113.785 130.555 114.310 130.775 ;
        RECT 113.730 129.790 113.970 130.385 ;
        RECT 114.140 129.855 114.310 130.555 ;
        RECT 114.480 130.195 114.650 130.975 ;
        RECT 114.970 130.925 115.340 131.425 ;
        RECT 115.520 130.975 115.925 131.145 ;
        RECT 116.095 130.975 116.880 131.145 ;
        RECT 115.520 130.745 115.690 130.975 ;
        RECT 114.860 130.445 115.690 130.745 ;
        RECT 116.075 130.475 116.540 130.805 ;
        RECT 114.860 130.415 115.060 130.445 ;
        RECT 115.180 130.195 115.350 130.265 ;
        RECT 114.480 130.025 115.350 130.195 ;
        RECT 114.840 129.935 115.350 130.025 ;
        RECT 113.390 129.470 113.695 129.600 ;
        RECT 114.140 129.490 114.670 129.855 ;
        RECT 113.010 128.875 113.275 129.335 ;
        RECT 113.445 129.045 113.695 129.470 ;
        RECT 114.840 129.320 115.010 129.935 ;
        RECT 113.905 129.150 115.010 129.320 ;
        RECT 115.180 128.875 115.350 129.675 ;
        RECT 115.520 129.375 115.690 130.445 ;
        RECT 115.860 129.545 116.050 130.265 ;
        RECT 116.220 129.515 116.540 130.475 ;
        RECT 116.710 130.515 116.880 130.975 ;
        RECT 117.155 130.895 117.365 131.425 ;
        RECT 117.625 130.685 117.955 131.210 ;
        RECT 118.125 130.815 118.295 131.425 ;
        RECT 118.465 130.770 118.795 131.205 ;
        RECT 118.465 130.685 118.845 130.770 ;
        RECT 117.755 130.515 117.955 130.685 ;
        RECT 118.620 130.645 118.845 130.685 ;
        RECT 116.710 130.185 117.585 130.515 ;
        RECT 117.755 130.185 118.505 130.515 ;
        RECT 115.520 129.045 115.770 129.375 ;
        RECT 116.710 129.345 116.880 130.185 ;
        RECT 117.755 129.980 117.945 130.185 ;
        RECT 118.675 130.065 118.845 130.645 ;
        RECT 119.015 130.675 120.225 131.425 ;
        RECT 120.395 130.700 120.685 131.425 ;
        RECT 120.875 130.735 121.115 131.255 ;
        RECT 121.285 130.930 121.680 131.425 ;
        RECT 122.245 131.095 122.415 131.240 ;
        RECT 122.040 130.900 122.415 131.095 ;
        RECT 119.015 130.135 119.535 130.675 ;
        RECT 118.630 130.015 118.845 130.065 ;
        RECT 117.050 129.605 117.945 129.980 ;
        RECT 118.455 129.935 118.845 130.015 ;
        RECT 119.705 129.965 120.225 130.505 ;
        RECT 115.995 129.175 116.880 129.345 ;
        RECT 117.060 128.875 117.375 129.375 ;
        RECT 117.605 129.045 117.945 129.605 ;
        RECT 118.115 128.875 118.285 129.885 ;
        RECT 118.455 129.090 118.785 129.935 ;
        RECT 119.015 128.875 120.225 129.965 ;
        RECT 120.395 128.875 120.685 130.040 ;
        RECT 120.875 129.930 121.050 130.735 ;
        RECT 122.040 130.565 122.210 130.900 ;
        RECT 122.695 130.855 122.935 131.230 ;
        RECT 123.105 130.920 123.440 131.425 ;
        RECT 123.615 130.880 128.960 131.425 ;
        RECT 129.600 130.920 129.935 131.425 ;
        RECT 122.695 130.705 122.915 130.855 ;
        RECT 121.225 130.205 122.210 130.565 ;
        RECT 122.380 130.375 122.915 130.705 ;
        RECT 121.225 130.185 122.510 130.205 ;
        RECT 121.650 130.035 122.510 130.185 ;
        RECT 120.875 129.145 121.180 129.930 ;
        RECT 121.355 129.555 122.050 129.865 ;
        RECT 121.360 128.875 122.045 129.345 ;
        RECT 122.225 129.090 122.510 130.035 ;
        RECT 122.680 129.725 122.915 130.375 ;
        RECT 123.085 129.895 123.385 130.745 ;
        RECT 125.200 130.050 125.540 130.880 ;
        RECT 130.105 130.855 130.345 131.230 ;
        RECT 130.625 131.095 130.795 131.240 ;
        RECT 130.625 130.900 131.000 131.095 ;
        RECT 131.360 130.930 131.755 131.425 ;
        RECT 122.680 129.495 123.355 129.725 ;
        RECT 122.685 128.875 123.015 129.325 ;
        RECT 123.185 129.065 123.355 129.495 ;
        RECT 127.020 129.310 127.370 130.560 ;
        RECT 129.655 129.895 129.955 130.745 ;
        RECT 130.125 130.705 130.345 130.855 ;
        RECT 130.125 130.375 130.660 130.705 ;
        RECT 130.830 130.565 131.000 130.900 ;
        RECT 131.925 130.735 132.165 131.255 ;
        RECT 130.125 129.725 130.360 130.375 ;
        RECT 130.830 130.205 131.815 130.565 ;
        RECT 129.685 129.495 130.360 129.725 ;
        RECT 130.530 130.185 131.815 130.205 ;
        RECT 130.530 130.035 131.390 130.185 ;
        RECT 123.615 128.875 128.960 129.310 ;
        RECT 129.685 129.065 129.855 129.495 ;
        RECT 130.025 128.875 130.355 129.325 ;
        RECT 130.530 129.090 130.815 130.035 ;
        RECT 131.990 129.930 132.165 130.735 ;
        RECT 132.355 130.655 134.945 131.425 ;
        RECT 135.580 130.685 135.835 131.255 ;
        RECT 136.005 131.025 136.335 131.425 ;
        RECT 136.760 130.890 137.290 131.255 ;
        RECT 137.480 131.085 137.755 131.255 ;
        RECT 137.475 130.915 137.755 131.085 ;
        RECT 136.760 130.855 136.935 130.890 ;
        RECT 136.005 130.685 136.935 130.855 ;
        RECT 132.355 130.135 133.565 130.655 ;
        RECT 133.735 129.965 134.945 130.485 ;
        RECT 130.990 129.555 131.685 129.865 ;
        RECT 130.995 128.875 131.680 129.345 ;
        RECT 131.860 129.145 132.165 129.930 ;
        RECT 132.355 128.875 134.945 129.965 ;
        RECT 135.580 130.015 135.750 130.685 ;
        RECT 136.005 130.515 136.175 130.685 ;
        RECT 135.920 130.185 136.175 130.515 ;
        RECT 136.400 130.185 136.595 130.515 ;
        RECT 135.580 129.045 135.915 130.015 ;
        RECT 136.085 128.875 136.255 130.015 ;
        RECT 136.425 129.215 136.595 130.185 ;
        RECT 136.765 129.555 136.935 130.685 ;
        RECT 137.105 129.895 137.275 130.695 ;
        RECT 137.480 130.095 137.755 130.915 ;
        RECT 137.925 129.895 138.115 131.255 ;
        RECT 138.295 130.890 138.805 131.425 ;
        RECT 139.025 130.615 139.270 131.220 ;
        RECT 139.715 130.880 145.060 131.425 ;
        RECT 138.315 130.445 139.545 130.615 ;
        RECT 137.105 129.725 138.115 129.895 ;
        RECT 138.285 129.880 139.035 130.070 ;
        RECT 136.765 129.385 137.890 129.555 ;
        RECT 138.285 129.215 138.455 129.880 ;
        RECT 139.205 129.635 139.545 130.445 ;
        RECT 141.300 130.050 141.640 130.880 ;
        RECT 145.695 130.675 146.905 131.425 ;
        RECT 136.425 129.045 138.455 129.215 ;
        RECT 138.625 128.875 138.795 129.635 ;
        RECT 139.030 129.225 139.545 129.635 ;
        RECT 143.120 129.310 143.470 130.560 ;
        RECT 145.695 129.965 146.215 130.505 ;
        RECT 146.385 130.135 146.905 130.675 ;
        RECT 139.715 128.875 145.060 129.310 ;
        RECT 145.695 128.875 146.905 129.965 ;
        RECT 17.270 128.705 146.990 128.875 ;
        RECT 17.355 127.615 18.565 128.705 ;
        RECT 17.355 126.905 17.875 127.445 ;
        RECT 18.045 127.075 18.565 127.615 ;
        RECT 18.740 127.555 19.000 128.705 ;
        RECT 19.175 127.630 19.430 128.535 ;
        RECT 19.600 127.945 19.930 128.705 ;
        RECT 20.145 127.775 20.315 128.535 ;
        RECT 17.355 126.155 18.565 126.905 ;
        RECT 18.740 126.155 19.000 126.995 ;
        RECT 19.175 126.900 19.345 127.630 ;
        RECT 19.600 127.605 20.315 127.775 ;
        RECT 19.600 127.395 19.770 127.605 ;
        RECT 20.580 127.555 20.840 128.705 ;
        RECT 21.015 127.630 21.270 128.535 ;
        RECT 21.440 127.945 21.770 128.705 ;
        RECT 21.985 127.775 22.155 128.535 ;
        RECT 19.515 127.065 19.770 127.395 ;
        RECT 19.175 126.325 19.430 126.900 ;
        RECT 19.600 126.875 19.770 127.065 ;
        RECT 20.050 127.055 20.405 127.425 ;
        RECT 19.600 126.705 20.315 126.875 ;
        RECT 19.600 126.155 19.930 126.535 ;
        RECT 20.145 126.325 20.315 126.705 ;
        RECT 20.580 126.155 20.840 126.995 ;
        RECT 21.015 126.900 21.185 127.630 ;
        RECT 21.440 127.605 22.155 127.775 ;
        RECT 22.415 127.615 25.925 128.705 ;
        RECT 21.440 127.395 21.610 127.605 ;
        RECT 21.355 127.065 21.610 127.395 ;
        RECT 21.015 126.325 21.270 126.900 ;
        RECT 21.440 126.875 21.610 127.065 ;
        RECT 21.890 127.055 22.245 127.425 ;
        RECT 22.415 126.925 24.065 127.445 ;
        RECT 24.235 127.095 25.925 127.615 ;
        RECT 26.280 127.735 26.670 127.910 ;
        RECT 27.155 127.905 27.485 128.705 ;
        RECT 27.655 127.915 28.190 128.535 ;
        RECT 26.280 127.565 27.705 127.735 ;
        RECT 21.440 126.705 22.155 126.875 ;
        RECT 21.440 126.155 21.770 126.535 ;
        RECT 21.985 126.325 22.155 126.705 ;
        RECT 22.415 126.155 25.925 126.925 ;
        RECT 26.155 126.835 26.510 127.395 ;
        RECT 26.680 126.665 26.850 127.565 ;
        RECT 27.020 126.835 27.285 127.395 ;
        RECT 27.535 127.065 27.705 127.565 ;
        RECT 27.875 126.895 28.190 127.915 ;
        RECT 28.395 127.615 30.065 128.705 ;
        RECT 26.260 126.155 26.500 126.665 ;
        RECT 26.680 126.335 26.960 126.665 ;
        RECT 27.190 126.155 27.405 126.665 ;
        RECT 27.575 126.325 28.190 126.895 ;
        RECT 28.395 126.925 29.145 127.445 ;
        RECT 29.315 127.095 30.065 127.615 ;
        RECT 30.235 127.540 30.525 128.705 ;
        RECT 30.695 128.270 36.040 128.705 ;
        RECT 36.215 128.270 41.560 128.705 ;
        RECT 41.735 128.270 47.080 128.705 ;
        RECT 47.255 128.270 52.600 128.705 ;
        RECT 28.395 126.155 30.065 126.925 ;
        RECT 30.235 126.155 30.525 126.880 ;
        RECT 32.280 126.700 32.620 127.530 ;
        RECT 34.100 127.020 34.450 128.270 ;
        RECT 37.800 126.700 38.140 127.530 ;
        RECT 39.620 127.020 39.970 128.270 ;
        RECT 43.320 126.700 43.660 127.530 ;
        RECT 45.140 127.020 45.490 128.270 ;
        RECT 48.840 126.700 49.180 127.530 ;
        RECT 50.660 127.020 51.010 128.270 ;
        RECT 52.775 127.615 55.365 128.705 ;
        RECT 52.775 126.925 53.985 127.445 ;
        RECT 54.155 127.095 55.365 127.615 ;
        RECT 55.995 127.540 56.285 128.705 ;
        RECT 56.455 128.270 61.800 128.705 ;
        RECT 30.695 126.155 36.040 126.700 ;
        RECT 36.215 126.155 41.560 126.700 ;
        RECT 41.735 126.155 47.080 126.700 ;
        RECT 47.255 126.155 52.600 126.700 ;
        RECT 52.775 126.155 55.365 126.925 ;
        RECT 55.995 126.155 56.285 126.880 ;
        RECT 58.040 126.700 58.380 127.530 ;
        RECT 59.860 127.020 60.210 128.270 ;
        RECT 61.975 127.615 64.565 128.705 ;
        RECT 61.975 126.925 63.185 127.445 ;
        RECT 63.355 127.095 64.565 127.615 ;
        RECT 64.740 127.565 65.075 128.535 ;
        RECT 65.245 127.565 65.415 128.705 ;
        RECT 65.585 128.365 67.615 128.535 ;
        RECT 56.455 126.155 61.800 126.700 ;
        RECT 61.975 126.155 64.565 126.925 ;
        RECT 64.740 126.895 64.910 127.565 ;
        RECT 65.585 127.395 65.755 128.365 ;
        RECT 65.080 127.065 65.335 127.395 ;
        RECT 65.560 127.065 65.755 127.395 ;
        RECT 65.925 128.025 67.050 128.195 ;
        RECT 65.165 126.895 65.335 127.065 ;
        RECT 65.925 126.895 66.095 128.025 ;
        RECT 64.740 126.325 64.995 126.895 ;
        RECT 65.165 126.725 66.095 126.895 ;
        RECT 66.265 127.685 67.275 127.855 ;
        RECT 66.265 126.885 66.435 127.685 ;
        RECT 65.920 126.690 66.095 126.725 ;
        RECT 65.165 126.155 65.495 126.555 ;
        RECT 65.920 126.325 66.450 126.690 ;
        RECT 66.640 126.665 66.915 127.485 ;
        RECT 66.635 126.495 66.915 126.665 ;
        RECT 66.640 126.325 66.915 126.495 ;
        RECT 67.085 126.325 67.275 127.685 ;
        RECT 67.445 127.700 67.615 128.365 ;
        RECT 67.785 127.945 67.955 128.705 ;
        RECT 68.190 127.945 68.705 128.355 ;
        RECT 67.445 127.510 68.195 127.700 ;
        RECT 68.365 127.135 68.705 127.945 ;
        RECT 68.875 127.615 71.465 128.705 ;
        RECT 67.475 126.965 68.705 127.135 ;
        RECT 67.455 126.155 67.965 126.690 ;
        RECT 68.185 126.360 68.430 126.965 ;
        RECT 68.875 126.925 70.085 127.445 ;
        RECT 70.255 127.095 71.465 127.615 ;
        RECT 71.640 127.565 71.975 128.535 ;
        RECT 72.145 127.565 72.315 128.705 ;
        RECT 72.485 128.365 74.515 128.535 ;
        RECT 68.875 126.155 71.465 126.925 ;
        RECT 71.640 126.895 71.810 127.565 ;
        RECT 72.485 127.395 72.655 128.365 ;
        RECT 71.980 127.065 72.235 127.395 ;
        RECT 72.460 127.065 72.655 127.395 ;
        RECT 72.825 128.025 73.950 128.195 ;
        RECT 72.065 126.895 72.235 127.065 ;
        RECT 72.825 126.895 72.995 128.025 ;
        RECT 71.640 126.325 71.895 126.895 ;
        RECT 72.065 126.725 72.995 126.895 ;
        RECT 73.165 127.685 74.175 127.855 ;
        RECT 73.165 126.885 73.335 127.685 ;
        RECT 73.540 127.005 73.815 127.485 ;
        RECT 73.535 126.835 73.815 127.005 ;
        RECT 72.820 126.690 72.995 126.725 ;
        RECT 72.065 126.155 72.395 126.555 ;
        RECT 72.820 126.325 73.350 126.690 ;
        RECT 73.540 126.325 73.815 126.835 ;
        RECT 73.985 126.325 74.175 127.685 ;
        RECT 74.345 127.700 74.515 128.365 ;
        RECT 74.685 127.945 74.855 128.705 ;
        RECT 75.090 127.945 75.605 128.355 ;
        RECT 75.775 128.270 81.120 128.705 ;
        RECT 74.345 127.510 75.095 127.700 ;
        RECT 75.265 127.135 75.605 127.945 ;
        RECT 74.375 126.965 75.605 127.135 ;
        RECT 74.355 126.155 74.865 126.690 ;
        RECT 75.085 126.360 75.330 126.965 ;
        RECT 77.360 126.700 77.700 127.530 ;
        RECT 79.180 127.020 79.530 128.270 ;
        RECT 81.755 127.540 82.045 128.705 ;
        RECT 82.220 127.565 82.555 128.535 ;
        RECT 82.725 127.565 82.895 128.705 ;
        RECT 83.065 128.365 85.095 128.535 ;
        RECT 82.220 126.895 82.390 127.565 ;
        RECT 83.065 127.395 83.235 128.365 ;
        RECT 82.560 127.065 82.815 127.395 ;
        RECT 83.040 127.065 83.235 127.395 ;
        RECT 83.405 128.025 84.530 128.195 ;
        RECT 82.645 126.895 82.815 127.065 ;
        RECT 83.405 126.895 83.575 128.025 ;
        RECT 75.775 126.155 81.120 126.700 ;
        RECT 81.755 126.155 82.045 126.880 ;
        RECT 82.220 126.325 82.475 126.895 ;
        RECT 82.645 126.725 83.575 126.895 ;
        RECT 83.745 127.685 84.755 127.855 ;
        RECT 83.745 126.885 83.915 127.685 ;
        RECT 84.120 127.345 84.395 127.485 ;
        RECT 84.115 127.175 84.395 127.345 ;
        RECT 83.400 126.690 83.575 126.725 ;
        RECT 82.645 126.155 82.975 126.555 ;
        RECT 83.400 126.325 83.930 126.690 ;
        RECT 84.120 126.325 84.395 127.175 ;
        RECT 84.565 126.325 84.755 127.685 ;
        RECT 84.925 127.700 85.095 128.365 ;
        RECT 85.265 127.945 85.435 128.705 ;
        RECT 85.670 127.945 86.185 128.355 ;
        RECT 84.925 127.510 85.675 127.700 ;
        RECT 85.845 127.135 86.185 127.945 ;
        RECT 86.355 127.615 89.865 128.705 ;
        RECT 90.035 127.615 91.245 128.705 ;
        RECT 91.665 127.975 91.960 128.705 ;
        RECT 92.130 127.805 92.390 128.530 ;
        RECT 92.560 127.975 92.820 128.705 ;
        RECT 92.990 127.805 93.250 128.530 ;
        RECT 93.420 127.975 93.680 128.705 ;
        RECT 93.850 127.805 94.110 128.530 ;
        RECT 94.280 127.975 94.540 128.705 ;
        RECT 94.710 127.805 94.970 128.530 ;
        RECT 84.955 126.965 86.185 127.135 ;
        RECT 84.935 126.155 85.445 126.690 ;
        RECT 85.665 126.360 85.910 126.965 ;
        RECT 86.355 126.925 88.005 127.445 ;
        RECT 88.175 127.095 89.865 127.615 ;
        RECT 86.355 126.155 89.865 126.925 ;
        RECT 90.035 126.905 90.555 127.445 ;
        RECT 90.725 127.075 91.245 127.615 ;
        RECT 91.660 127.565 94.970 127.805 ;
        RECT 95.140 127.595 95.400 128.705 ;
        RECT 91.660 126.975 92.630 127.565 ;
        RECT 95.570 127.395 95.820 128.530 ;
        RECT 96.000 127.595 96.295 128.705 ;
        RECT 96.480 127.565 96.815 128.535 ;
        RECT 96.985 127.565 97.155 128.705 ;
        RECT 97.325 128.365 99.355 128.535 ;
        RECT 92.800 127.145 95.820 127.395 ;
        RECT 90.035 126.155 91.245 126.905 ;
        RECT 91.660 126.805 94.970 126.975 ;
        RECT 91.660 126.155 91.960 126.635 ;
        RECT 92.130 126.350 92.390 126.805 ;
        RECT 92.560 126.155 92.820 126.635 ;
        RECT 92.990 126.350 93.250 126.805 ;
        RECT 93.420 126.155 93.680 126.635 ;
        RECT 93.850 126.350 94.110 126.805 ;
        RECT 94.280 126.155 94.540 126.635 ;
        RECT 94.710 126.350 94.970 126.805 ;
        RECT 95.140 126.155 95.400 126.680 ;
        RECT 95.570 126.335 95.820 127.145 ;
        RECT 95.990 126.785 96.305 127.395 ;
        RECT 96.480 126.895 96.650 127.565 ;
        RECT 97.325 127.395 97.495 128.365 ;
        RECT 96.820 127.065 97.075 127.395 ;
        RECT 97.300 127.065 97.495 127.395 ;
        RECT 97.665 128.025 98.790 128.195 ;
        RECT 96.905 126.895 97.075 127.065 ;
        RECT 97.665 126.895 97.835 128.025 ;
        RECT 96.000 126.155 96.245 126.615 ;
        RECT 96.480 126.325 96.735 126.895 ;
        RECT 96.905 126.725 97.835 126.895 ;
        RECT 98.005 127.685 99.015 127.855 ;
        RECT 98.005 126.885 98.175 127.685 ;
        RECT 98.380 127.005 98.655 127.485 ;
        RECT 98.375 126.835 98.655 127.005 ;
        RECT 97.660 126.690 97.835 126.725 ;
        RECT 96.905 126.155 97.235 126.555 ;
        RECT 97.660 126.325 98.190 126.690 ;
        RECT 98.380 126.325 98.655 126.835 ;
        RECT 98.825 126.325 99.015 127.685 ;
        RECT 99.185 127.700 99.355 128.365 ;
        RECT 99.525 127.945 99.695 128.705 ;
        RECT 99.930 127.945 100.445 128.355 ;
        RECT 99.185 127.510 99.935 127.700 ;
        RECT 100.105 127.135 100.445 127.945 ;
        RECT 99.215 126.965 100.445 127.135 ;
        RECT 100.620 127.565 100.955 128.535 ;
        RECT 101.125 127.565 101.295 128.705 ;
        RECT 101.465 128.365 103.495 128.535 ;
        RECT 99.195 126.155 99.705 126.690 ;
        RECT 99.925 126.360 100.170 126.965 ;
        RECT 100.620 126.895 100.790 127.565 ;
        RECT 101.465 127.395 101.635 128.365 ;
        RECT 100.960 127.065 101.215 127.395 ;
        RECT 101.440 127.065 101.635 127.395 ;
        RECT 101.805 128.025 102.930 128.195 ;
        RECT 101.045 126.895 101.215 127.065 ;
        RECT 101.805 126.895 101.975 128.025 ;
        RECT 100.620 126.325 100.875 126.895 ;
        RECT 101.045 126.725 101.975 126.895 ;
        RECT 102.145 127.685 103.155 127.855 ;
        RECT 102.145 126.885 102.315 127.685 ;
        RECT 102.520 127.005 102.795 127.485 ;
        RECT 102.515 126.835 102.795 127.005 ;
        RECT 101.800 126.690 101.975 126.725 ;
        RECT 101.045 126.155 101.375 126.555 ;
        RECT 101.800 126.325 102.330 126.690 ;
        RECT 102.520 126.325 102.795 126.835 ;
        RECT 102.965 126.325 103.155 127.685 ;
        RECT 103.325 127.700 103.495 128.365 ;
        RECT 103.665 127.945 103.835 128.705 ;
        RECT 104.070 127.945 104.585 128.355 ;
        RECT 103.325 127.510 104.075 127.700 ;
        RECT 104.245 127.135 104.585 127.945 ;
        RECT 104.755 127.615 107.345 128.705 ;
        RECT 103.355 126.965 104.585 127.135 ;
        RECT 103.335 126.155 103.845 126.690 ;
        RECT 104.065 126.360 104.310 126.965 ;
        RECT 104.755 126.925 105.965 127.445 ;
        RECT 106.135 127.095 107.345 127.615 ;
        RECT 107.515 127.540 107.805 128.705 ;
        RECT 108.985 128.085 109.155 128.515 ;
        RECT 109.325 128.255 109.655 128.705 ;
        RECT 108.985 127.855 109.660 128.085 ;
        RECT 104.755 126.155 107.345 126.925 ;
        RECT 107.515 126.155 107.805 126.880 ;
        RECT 108.955 126.835 109.255 127.685 ;
        RECT 109.425 127.205 109.660 127.855 ;
        RECT 109.830 127.545 110.115 128.490 ;
        RECT 110.295 128.235 110.980 128.705 ;
        RECT 110.290 127.715 110.985 128.025 ;
        RECT 111.160 127.650 111.465 128.435 ;
        RECT 109.830 127.395 110.690 127.545 ;
        RECT 109.830 127.375 111.115 127.395 ;
        RECT 109.425 126.875 109.960 127.205 ;
        RECT 110.130 127.015 111.115 127.375 ;
        RECT 109.425 126.725 109.645 126.875 ;
        RECT 108.900 126.155 109.235 126.660 ;
        RECT 109.405 126.350 109.645 126.725 ;
        RECT 110.130 126.680 110.300 127.015 ;
        RECT 111.290 126.845 111.465 127.650 ;
        RECT 109.925 126.485 110.300 126.680 ;
        RECT 109.925 126.340 110.095 126.485 ;
        RECT 110.660 126.155 111.055 126.650 ;
        RECT 111.225 126.325 111.465 126.845 ;
        RECT 111.660 127.565 111.995 128.535 ;
        RECT 112.165 127.565 112.335 128.705 ;
        RECT 112.505 128.365 114.535 128.535 ;
        RECT 111.660 126.895 111.830 127.565 ;
        RECT 112.505 127.395 112.675 128.365 ;
        RECT 112.000 127.065 112.255 127.395 ;
        RECT 112.480 127.065 112.675 127.395 ;
        RECT 112.845 128.025 113.970 128.195 ;
        RECT 112.085 126.895 112.255 127.065 ;
        RECT 112.845 126.895 113.015 128.025 ;
        RECT 111.660 126.325 111.915 126.895 ;
        RECT 112.085 126.725 113.015 126.895 ;
        RECT 113.185 127.685 114.195 127.855 ;
        RECT 113.185 126.885 113.355 127.685 ;
        RECT 113.560 127.005 113.835 127.485 ;
        RECT 113.555 126.835 113.835 127.005 ;
        RECT 112.840 126.690 113.015 126.725 ;
        RECT 112.085 126.155 112.415 126.555 ;
        RECT 112.840 126.325 113.370 126.690 ;
        RECT 113.560 126.325 113.835 126.835 ;
        RECT 114.005 126.325 114.195 127.685 ;
        RECT 114.365 127.700 114.535 128.365 ;
        RECT 114.705 127.945 114.875 128.705 ;
        RECT 115.110 127.945 115.625 128.355 ;
        RECT 114.365 127.510 115.115 127.700 ;
        RECT 115.285 127.135 115.625 127.945 ;
        RECT 115.795 127.615 117.465 128.705 ;
        RECT 114.395 126.965 115.625 127.135 ;
        RECT 114.375 126.155 114.885 126.690 ;
        RECT 115.105 126.360 115.350 126.965 ;
        RECT 115.795 126.925 116.545 127.445 ;
        RECT 116.715 127.095 117.465 127.615 ;
        RECT 117.640 127.755 117.905 128.525 ;
        RECT 118.075 127.985 118.405 128.705 ;
        RECT 118.595 128.165 118.855 128.525 ;
        RECT 119.025 128.335 119.355 128.705 ;
        RECT 119.525 128.165 119.785 128.525 ;
        RECT 118.595 127.935 119.785 128.165 ;
        RECT 120.355 127.755 120.645 128.525 ;
        RECT 120.945 128.035 121.115 128.535 ;
        RECT 121.285 128.205 121.615 128.705 ;
        RECT 120.945 127.865 121.610 128.035 ;
        RECT 115.795 126.155 117.465 126.925 ;
        RECT 117.640 126.335 117.975 127.755 ;
        RECT 118.150 127.575 120.645 127.755 ;
        RECT 118.150 126.885 118.375 127.575 ;
        RECT 118.575 127.065 118.855 127.395 ;
        RECT 119.035 127.065 119.610 127.395 ;
        RECT 119.790 127.065 120.225 127.395 ;
        RECT 120.405 127.065 120.675 127.395 ;
        RECT 120.860 127.045 121.210 127.695 ;
        RECT 118.150 126.695 120.635 126.885 ;
        RECT 121.380 126.875 121.610 127.865 ;
        RECT 118.155 126.155 118.900 126.525 ;
        RECT 119.465 126.335 119.720 126.695 ;
        RECT 119.900 126.155 120.230 126.525 ;
        RECT 120.410 126.335 120.635 126.695 ;
        RECT 120.945 126.705 121.610 126.875 ;
        RECT 120.945 126.415 121.115 126.705 ;
        RECT 121.285 126.155 121.615 126.535 ;
        RECT 121.785 126.415 121.970 128.535 ;
        RECT 122.210 128.245 122.475 128.705 ;
        RECT 122.645 128.110 122.895 128.535 ;
        RECT 123.105 128.260 124.210 128.430 ;
        RECT 122.590 127.980 122.895 128.110 ;
        RECT 122.140 126.785 122.420 127.735 ;
        RECT 122.590 126.875 122.760 127.980 ;
        RECT 122.930 127.195 123.170 127.790 ;
        RECT 123.340 127.725 123.870 128.090 ;
        RECT 123.340 127.025 123.510 127.725 ;
        RECT 124.040 127.645 124.210 128.260 ;
        RECT 124.380 127.905 124.550 128.705 ;
        RECT 124.720 128.205 124.970 128.535 ;
        RECT 125.195 128.235 126.080 128.405 ;
        RECT 124.040 127.555 124.550 127.645 ;
        RECT 122.590 126.745 122.815 126.875 ;
        RECT 122.985 126.805 123.510 127.025 ;
        RECT 123.680 127.385 124.550 127.555 ;
        RECT 122.225 126.155 122.475 126.615 ;
        RECT 122.645 126.605 122.815 126.745 ;
        RECT 123.680 126.605 123.850 127.385 ;
        RECT 124.380 127.315 124.550 127.385 ;
        RECT 124.060 127.135 124.260 127.165 ;
        RECT 124.720 127.135 124.890 128.205 ;
        RECT 125.060 127.315 125.250 128.035 ;
        RECT 124.060 126.835 124.890 127.135 ;
        RECT 125.420 127.105 125.740 128.065 ;
        RECT 122.645 126.435 122.980 126.605 ;
        RECT 123.175 126.435 123.850 126.605 ;
        RECT 124.170 126.155 124.540 126.655 ;
        RECT 124.720 126.605 124.890 126.835 ;
        RECT 125.275 126.775 125.740 127.105 ;
        RECT 125.910 127.395 126.080 128.235 ;
        RECT 126.260 128.205 126.575 128.705 ;
        RECT 126.805 127.975 127.145 128.535 ;
        RECT 126.250 127.600 127.145 127.975 ;
        RECT 127.315 127.695 127.485 128.705 ;
        RECT 126.955 127.395 127.145 127.600 ;
        RECT 127.655 127.645 127.985 128.490 ;
        RECT 127.655 127.565 128.045 127.645 ;
        RECT 128.215 127.615 129.885 128.705 ;
        RECT 130.605 128.085 130.775 128.515 ;
        RECT 130.945 128.255 131.275 128.705 ;
        RECT 130.605 127.855 131.280 128.085 ;
        RECT 127.830 127.515 128.045 127.565 ;
        RECT 125.910 127.065 126.785 127.395 ;
        RECT 126.955 127.065 127.705 127.395 ;
        RECT 125.910 126.605 126.080 127.065 ;
        RECT 126.955 126.895 127.155 127.065 ;
        RECT 127.875 126.935 128.045 127.515 ;
        RECT 127.820 126.895 128.045 126.935 ;
        RECT 124.720 126.435 125.125 126.605 ;
        RECT 125.295 126.435 126.080 126.605 ;
        RECT 126.355 126.155 126.565 126.685 ;
        RECT 126.825 126.370 127.155 126.895 ;
        RECT 127.665 126.810 128.045 126.895 ;
        RECT 128.215 126.925 128.965 127.445 ;
        RECT 129.135 127.095 129.885 127.615 ;
        RECT 127.325 126.155 127.495 126.765 ;
        RECT 127.665 126.375 127.995 126.810 ;
        RECT 128.215 126.155 129.885 126.925 ;
        RECT 130.575 126.835 130.875 127.685 ;
        RECT 131.045 127.205 131.280 127.855 ;
        RECT 131.450 127.545 131.735 128.490 ;
        RECT 131.915 128.235 132.600 128.705 ;
        RECT 131.910 127.715 132.605 128.025 ;
        RECT 132.780 127.650 133.085 128.435 ;
        RECT 131.450 127.395 132.310 127.545 ;
        RECT 131.450 127.375 132.735 127.395 ;
        RECT 131.045 126.875 131.580 127.205 ;
        RECT 131.750 127.015 132.735 127.375 ;
        RECT 131.045 126.725 131.265 126.875 ;
        RECT 130.520 126.155 130.855 126.660 ;
        RECT 131.025 126.350 131.265 126.725 ;
        RECT 131.750 126.680 131.920 127.015 ;
        RECT 132.910 126.845 133.085 127.650 ;
        RECT 133.275 127.540 133.565 128.705 ;
        RECT 133.740 127.755 134.005 128.525 ;
        RECT 134.175 127.985 134.505 128.705 ;
        RECT 134.695 128.165 134.955 128.525 ;
        RECT 135.125 128.335 135.455 128.705 ;
        RECT 135.625 128.165 135.885 128.525 ;
        RECT 134.695 127.935 135.885 128.165 ;
        RECT 136.455 127.755 136.745 128.525 ;
        RECT 137.505 128.035 137.675 128.535 ;
        RECT 137.845 128.205 138.175 128.705 ;
        RECT 137.505 127.865 138.170 128.035 ;
        RECT 131.545 126.485 131.920 126.680 ;
        RECT 131.545 126.340 131.715 126.485 ;
        RECT 132.280 126.155 132.675 126.650 ;
        RECT 132.845 126.325 133.085 126.845 ;
        RECT 133.275 126.155 133.565 126.880 ;
        RECT 133.740 126.335 134.075 127.755 ;
        RECT 134.250 127.575 136.745 127.755 ;
        RECT 134.250 126.885 134.475 127.575 ;
        RECT 134.675 127.065 134.955 127.395 ;
        RECT 135.135 127.065 135.710 127.395 ;
        RECT 135.890 127.065 136.325 127.395 ;
        RECT 136.505 127.065 136.775 127.395 ;
        RECT 137.420 127.045 137.770 127.695 ;
        RECT 134.250 126.695 136.735 126.885 ;
        RECT 137.940 126.875 138.170 127.865 ;
        RECT 134.255 126.155 135.000 126.525 ;
        RECT 135.565 126.335 135.820 126.695 ;
        RECT 136.000 126.155 136.330 126.525 ;
        RECT 136.510 126.335 136.735 126.695 ;
        RECT 137.505 126.705 138.170 126.875 ;
        RECT 137.505 126.415 137.675 126.705 ;
        RECT 137.845 126.155 138.175 126.535 ;
        RECT 138.345 126.415 138.530 128.535 ;
        RECT 138.770 128.245 139.035 128.705 ;
        RECT 139.205 128.110 139.455 128.535 ;
        RECT 139.665 128.260 140.770 128.430 ;
        RECT 139.150 127.980 139.455 128.110 ;
        RECT 138.700 126.785 138.980 127.735 ;
        RECT 139.150 126.875 139.320 127.980 ;
        RECT 139.490 127.195 139.730 127.790 ;
        RECT 139.900 127.725 140.430 128.090 ;
        RECT 139.900 127.025 140.070 127.725 ;
        RECT 140.600 127.645 140.770 128.260 ;
        RECT 140.940 127.905 141.110 128.705 ;
        RECT 141.280 128.205 141.530 128.535 ;
        RECT 141.755 128.235 142.640 128.405 ;
        RECT 140.600 127.555 141.110 127.645 ;
        RECT 139.150 126.745 139.375 126.875 ;
        RECT 139.545 126.805 140.070 127.025 ;
        RECT 140.240 127.385 141.110 127.555 ;
        RECT 138.785 126.155 139.035 126.615 ;
        RECT 139.205 126.605 139.375 126.745 ;
        RECT 140.240 126.605 140.410 127.385 ;
        RECT 140.940 127.315 141.110 127.385 ;
        RECT 140.620 127.135 140.820 127.165 ;
        RECT 141.280 127.135 141.450 128.205 ;
        RECT 141.620 127.315 141.810 128.035 ;
        RECT 140.620 126.835 141.450 127.135 ;
        RECT 141.980 127.105 142.300 128.065 ;
        RECT 139.205 126.435 139.540 126.605 ;
        RECT 139.735 126.435 140.410 126.605 ;
        RECT 140.730 126.155 141.100 126.655 ;
        RECT 141.280 126.605 141.450 126.835 ;
        RECT 141.835 126.775 142.300 127.105 ;
        RECT 142.470 127.395 142.640 128.235 ;
        RECT 142.820 128.205 143.135 128.705 ;
        RECT 143.365 127.975 143.705 128.535 ;
        RECT 142.810 127.600 143.705 127.975 ;
        RECT 143.875 127.695 144.045 128.705 ;
        RECT 143.515 127.395 143.705 127.600 ;
        RECT 144.215 127.645 144.545 128.490 ;
        RECT 144.215 127.565 144.605 127.645 ;
        RECT 144.390 127.515 144.605 127.565 ;
        RECT 142.470 127.065 143.345 127.395 ;
        RECT 143.515 127.065 144.265 127.395 ;
        RECT 142.470 126.605 142.640 127.065 ;
        RECT 143.515 126.895 143.715 127.065 ;
        RECT 144.435 126.935 144.605 127.515 ;
        RECT 145.695 127.615 146.905 128.705 ;
        RECT 145.695 127.075 146.215 127.615 ;
        RECT 144.380 126.895 144.605 126.935 ;
        RECT 146.385 126.905 146.905 127.445 ;
        RECT 141.280 126.435 141.685 126.605 ;
        RECT 141.855 126.435 142.640 126.605 ;
        RECT 142.915 126.155 143.125 126.685 ;
        RECT 143.385 126.370 143.715 126.895 ;
        RECT 144.225 126.810 144.605 126.895 ;
        RECT 143.885 126.155 144.055 126.765 ;
        RECT 144.225 126.375 144.555 126.810 ;
        RECT 145.695 126.155 146.905 126.905 ;
        RECT 17.270 125.985 146.990 126.155 ;
        RECT 17.355 125.235 18.565 125.985 ;
        RECT 19.655 125.485 19.915 125.815 ;
        RECT 20.125 125.505 20.400 125.985 ;
        RECT 17.355 124.695 17.875 125.235 ;
        RECT 18.045 124.525 18.565 125.065 ;
        RECT 17.355 123.435 18.565 124.525 ;
        RECT 19.655 124.575 19.825 125.485 ;
        RECT 20.610 125.415 20.815 125.815 ;
        RECT 20.985 125.585 21.320 125.985 ;
        RECT 19.995 124.745 20.355 125.325 ;
        RECT 20.610 125.245 21.295 125.415 ;
        RECT 20.535 124.575 20.785 125.075 ;
        RECT 19.655 124.405 20.785 124.575 ;
        RECT 19.655 123.635 19.925 124.405 ;
        RECT 20.955 124.215 21.295 125.245 ;
        RECT 21.495 125.235 22.705 125.985 ;
        RECT 22.925 125.330 23.255 125.765 ;
        RECT 23.425 125.375 23.595 125.985 ;
        RECT 22.875 125.245 23.255 125.330 ;
        RECT 23.765 125.245 24.095 125.770 ;
        RECT 24.355 125.455 24.565 125.985 ;
        RECT 24.840 125.535 25.625 125.705 ;
        RECT 25.795 125.535 26.200 125.705 ;
        RECT 21.495 124.695 22.015 125.235 ;
        RECT 22.875 125.205 23.100 125.245 ;
        RECT 22.185 124.525 22.705 125.065 ;
        RECT 20.095 123.435 20.425 124.215 ;
        RECT 20.630 124.040 21.295 124.215 ;
        RECT 20.630 123.635 20.815 124.040 ;
        RECT 20.985 123.435 21.320 123.860 ;
        RECT 21.495 123.435 22.705 124.525 ;
        RECT 22.875 124.625 23.045 125.205 ;
        RECT 23.765 125.075 23.965 125.245 ;
        RECT 24.840 125.075 25.010 125.535 ;
        RECT 23.215 124.745 23.965 125.075 ;
        RECT 24.135 124.745 25.010 125.075 ;
        RECT 22.875 124.575 23.090 124.625 ;
        RECT 22.875 124.495 23.265 124.575 ;
        RECT 22.935 123.650 23.265 124.495 ;
        RECT 23.775 124.540 23.965 124.745 ;
        RECT 23.435 123.435 23.605 124.445 ;
        RECT 23.775 124.165 24.670 124.540 ;
        RECT 23.775 123.605 24.115 124.165 ;
        RECT 24.345 123.435 24.660 123.935 ;
        RECT 24.840 123.905 25.010 124.745 ;
        RECT 25.180 125.035 25.645 125.365 ;
        RECT 26.030 125.305 26.200 125.535 ;
        RECT 26.380 125.485 26.750 125.985 ;
        RECT 27.070 125.535 27.745 125.705 ;
        RECT 27.940 125.535 28.275 125.705 ;
        RECT 25.180 124.075 25.500 125.035 ;
        RECT 26.030 125.005 26.860 125.305 ;
        RECT 25.670 124.105 25.860 124.825 ;
        RECT 26.030 123.935 26.200 125.005 ;
        RECT 26.660 124.975 26.860 125.005 ;
        RECT 26.370 124.755 26.540 124.825 ;
        RECT 27.070 124.755 27.240 125.535 ;
        RECT 28.105 125.395 28.275 125.535 ;
        RECT 28.445 125.525 28.695 125.985 ;
        RECT 26.370 124.585 27.240 124.755 ;
        RECT 27.410 125.115 27.935 125.335 ;
        RECT 28.105 125.265 28.330 125.395 ;
        RECT 26.370 124.495 26.880 124.585 ;
        RECT 24.840 123.735 25.725 123.905 ;
        RECT 25.950 123.605 26.200 123.935 ;
        RECT 26.370 123.435 26.540 124.235 ;
        RECT 26.710 123.880 26.880 124.495 ;
        RECT 27.410 124.415 27.580 125.115 ;
        RECT 27.050 124.050 27.580 124.415 ;
        RECT 27.750 124.350 27.990 124.945 ;
        RECT 28.160 124.160 28.330 125.265 ;
        RECT 28.500 124.405 28.780 125.355 ;
        RECT 28.025 124.030 28.330 124.160 ;
        RECT 26.710 123.710 27.815 123.880 ;
        RECT 28.025 123.605 28.275 124.030 ;
        RECT 28.445 123.435 28.710 123.895 ;
        RECT 28.950 123.605 29.135 125.725 ;
        RECT 29.305 125.605 29.635 125.985 ;
        RECT 29.805 125.435 29.975 125.725 ;
        RECT 29.310 125.265 29.975 125.435 ;
        RECT 29.310 124.275 29.540 125.265 ;
        RECT 30.235 125.185 30.575 125.815 ;
        RECT 30.865 125.525 31.035 125.985 ;
        RECT 31.305 125.355 31.635 125.800 ;
        RECT 29.710 124.445 30.060 125.095 ;
        RECT 30.235 124.615 30.505 125.185 ;
        RECT 30.885 125.165 31.635 125.355 ;
        RECT 31.805 125.335 31.975 125.655 ;
        RECT 32.200 125.525 32.530 125.985 ;
        RECT 32.730 125.335 33.060 125.815 ;
        RECT 33.275 125.525 33.605 125.985 ;
        RECT 33.775 125.335 34.105 125.815 ;
        RECT 34.375 125.440 39.720 125.985 ;
        RECT 31.805 125.165 34.105 125.335 ;
        RECT 30.885 124.995 31.255 125.165 ;
        RECT 30.675 124.785 31.255 124.995 ;
        RECT 31.425 124.785 31.845 124.995 ;
        RECT 30.995 124.615 31.255 124.785 ;
        RECT 29.310 124.105 29.975 124.275 ;
        RECT 29.305 123.435 29.635 123.935 ;
        RECT 29.805 123.605 29.975 124.105 ;
        RECT 30.235 123.605 30.760 124.615 ;
        RECT 30.995 124.325 31.745 124.615 ;
        RECT 30.995 123.435 31.325 124.155 ;
        RECT 31.495 123.605 31.745 124.325 ;
        RECT 32.015 123.680 32.345 124.995 ;
        RECT 32.555 123.680 32.885 124.995 ;
        RECT 33.055 123.680 33.425 124.995 ;
        RECT 33.635 124.745 34.145 124.995 ;
        RECT 35.960 124.610 36.300 125.440 ;
        RECT 39.895 125.215 42.485 125.985 ;
        RECT 43.115 125.260 43.405 125.985 ;
        RECT 43.575 125.440 48.920 125.985 ;
        RECT 49.095 125.440 54.440 125.985 ;
        RECT 54.615 125.440 59.960 125.985 ;
        RECT 60.135 125.440 65.480 125.985 ;
        RECT 33.755 123.435 34.085 124.555 ;
        RECT 37.780 123.870 38.130 125.120 ;
        RECT 39.895 124.695 41.105 125.215 ;
        RECT 41.275 124.525 42.485 125.045 ;
        RECT 45.160 124.610 45.500 125.440 ;
        RECT 34.375 123.435 39.720 123.870 ;
        RECT 39.895 123.435 42.485 124.525 ;
        RECT 43.115 123.435 43.405 124.600 ;
        RECT 46.980 123.870 47.330 125.120 ;
        RECT 50.680 124.610 51.020 125.440 ;
        RECT 52.500 123.870 52.850 125.120 ;
        RECT 56.200 124.610 56.540 125.440 ;
        RECT 58.020 123.870 58.370 125.120 ;
        RECT 61.720 124.610 62.060 125.440 ;
        RECT 65.655 125.215 68.245 125.985 ;
        RECT 68.875 125.260 69.165 125.985 ;
        RECT 69.335 125.440 74.680 125.985 ;
        RECT 74.855 125.440 80.200 125.985 ;
        RECT 80.375 125.440 85.720 125.985 ;
        RECT 86.825 125.495 87.155 125.985 ;
        RECT 63.540 123.870 63.890 125.120 ;
        RECT 65.655 124.695 66.865 125.215 ;
        RECT 67.035 124.525 68.245 125.045 ;
        RECT 70.920 124.610 71.260 125.440 ;
        RECT 43.575 123.435 48.920 123.870 ;
        RECT 49.095 123.435 54.440 123.870 ;
        RECT 54.615 123.435 59.960 123.870 ;
        RECT 60.135 123.435 65.480 123.870 ;
        RECT 65.655 123.435 68.245 124.525 ;
        RECT 68.875 123.435 69.165 124.600 ;
        RECT 72.740 123.870 73.090 125.120 ;
        RECT 76.440 124.610 76.780 125.440 ;
        RECT 78.260 123.870 78.610 125.120 ;
        RECT 81.960 124.610 82.300 125.440 ;
        RECT 87.325 125.390 87.945 125.815 ;
        RECT 83.780 123.870 84.130 125.120 ;
        RECT 86.815 124.745 87.155 125.325 ;
        RECT 87.325 125.055 87.685 125.390 ;
        RECT 88.405 125.295 88.735 125.985 ;
        RECT 89.635 125.525 89.880 125.985 ;
        RECT 87.325 124.775 88.745 125.055 ;
        RECT 69.335 123.435 74.680 123.870 ;
        RECT 74.855 123.435 80.200 123.870 ;
        RECT 80.375 123.435 85.720 123.870 ;
        RECT 86.825 123.435 87.155 124.575 ;
        RECT 87.325 123.605 87.685 124.775 ;
        RECT 87.885 123.435 88.215 124.605 ;
        RECT 88.415 123.605 88.745 124.775 ;
        RECT 89.575 124.745 89.890 125.355 ;
        RECT 90.060 124.995 90.310 125.805 ;
        RECT 90.480 125.460 90.740 125.985 ;
        RECT 90.910 125.335 91.170 125.790 ;
        RECT 91.340 125.505 91.600 125.985 ;
        RECT 91.770 125.335 92.030 125.790 ;
        RECT 92.200 125.505 92.460 125.985 ;
        RECT 92.630 125.335 92.890 125.790 ;
        RECT 93.060 125.505 93.320 125.985 ;
        RECT 93.490 125.335 93.750 125.790 ;
        RECT 93.920 125.505 94.220 125.985 ;
        RECT 90.910 125.165 94.220 125.335 ;
        RECT 94.635 125.260 94.925 125.985 ;
        RECT 95.185 125.435 95.355 125.725 ;
        RECT 95.525 125.605 95.855 125.985 ;
        RECT 95.185 125.265 95.850 125.435 ;
        RECT 90.060 124.745 93.080 124.995 ;
        RECT 88.945 123.435 89.275 124.605 ;
        RECT 89.585 123.435 89.880 124.545 ;
        RECT 90.060 123.610 90.310 124.745 ;
        RECT 93.250 124.575 94.220 125.165 ;
        RECT 90.480 123.435 90.740 124.545 ;
        RECT 90.910 124.335 94.220 124.575 ;
        RECT 90.910 123.610 91.170 124.335 ;
        RECT 91.340 123.435 91.600 124.165 ;
        RECT 91.770 123.610 92.030 124.335 ;
        RECT 92.200 123.435 92.460 124.165 ;
        RECT 92.630 123.610 92.890 124.335 ;
        RECT 93.060 123.435 93.320 124.165 ;
        RECT 93.490 123.610 93.750 124.335 ;
        RECT 93.920 123.435 94.215 124.165 ;
        RECT 94.635 123.435 94.925 124.600 ;
        RECT 95.100 124.445 95.450 125.095 ;
        RECT 95.620 124.275 95.850 125.265 ;
        RECT 95.185 124.105 95.850 124.275 ;
        RECT 95.185 123.605 95.355 124.105 ;
        RECT 95.525 123.435 95.855 123.935 ;
        RECT 96.025 123.605 96.210 125.725 ;
        RECT 96.465 125.525 96.715 125.985 ;
        RECT 96.885 125.535 97.220 125.705 ;
        RECT 97.415 125.535 98.090 125.705 ;
        RECT 96.885 125.395 97.055 125.535 ;
        RECT 96.380 124.405 96.660 125.355 ;
        RECT 96.830 125.265 97.055 125.395 ;
        RECT 96.830 124.160 97.000 125.265 ;
        RECT 97.225 125.115 97.750 125.335 ;
        RECT 97.170 124.350 97.410 124.945 ;
        RECT 97.580 124.415 97.750 125.115 ;
        RECT 97.920 124.755 98.090 125.535 ;
        RECT 98.410 125.485 98.780 125.985 ;
        RECT 98.960 125.535 99.365 125.705 ;
        RECT 99.535 125.535 100.320 125.705 ;
        RECT 98.960 125.305 99.130 125.535 ;
        RECT 98.300 125.005 99.130 125.305 ;
        RECT 99.515 125.035 99.980 125.365 ;
        RECT 98.300 124.975 98.500 125.005 ;
        RECT 98.620 124.755 98.790 124.825 ;
        RECT 97.920 124.585 98.790 124.755 ;
        RECT 98.280 124.495 98.790 124.585 ;
        RECT 96.830 124.030 97.135 124.160 ;
        RECT 97.580 124.050 98.110 124.415 ;
        RECT 96.450 123.435 96.715 123.895 ;
        RECT 96.885 123.605 97.135 124.030 ;
        RECT 98.280 123.880 98.450 124.495 ;
        RECT 97.345 123.710 98.450 123.880 ;
        RECT 98.620 123.435 98.790 124.235 ;
        RECT 98.960 123.935 99.130 125.005 ;
        RECT 99.300 124.105 99.490 124.825 ;
        RECT 99.660 124.075 99.980 125.035 ;
        RECT 100.150 125.075 100.320 125.535 ;
        RECT 100.595 125.455 100.805 125.985 ;
        RECT 101.065 125.245 101.395 125.770 ;
        RECT 101.565 125.375 101.735 125.985 ;
        RECT 101.905 125.330 102.235 125.765 ;
        RECT 102.525 125.585 102.855 125.985 ;
        RECT 103.025 125.415 103.195 125.685 ;
        RECT 103.365 125.585 103.695 125.985 ;
        RECT 103.865 125.415 104.120 125.685 ;
        RECT 104.295 125.440 109.640 125.985 ;
        RECT 101.905 125.245 102.285 125.330 ;
        RECT 101.195 125.075 101.395 125.245 ;
        RECT 102.060 125.205 102.285 125.245 ;
        RECT 100.150 124.745 101.025 125.075 ;
        RECT 101.195 124.745 101.945 125.075 ;
        RECT 98.960 123.605 99.210 123.935 ;
        RECT 100.150 123.905 100.320 124.745 ;
        RECT 101.195 124.540 101.385 124.745 ;
        RECT 102.115 124.625 102.285 125.205 ;
        RECT 102.070 124.575 102.285 124.625 ;
        RECT 100.490 124.165 101.385 124.540 ;
        RECT 101.895 124.495 102.285 124.575 ;
        RECT 99.435 123.735 100.320 123.905 ;
        RECT 100.500 123.435 100.815 123.935 ;
        RECT 101.045 123.605 101.385 124.165 ;
        RECT 101.555 123.435 101.725 124.445 ;
        RECT 101.895 123.650 102.225 124.495 ;
        RECT 102.455 124.405 102.725 125.415 ;
        RECT 102.895 125.245 104.120 125.415 ;
        RECT 102.895 124.575 103.065 125.245 ;
        RECT 103.235 124.745 103.615 125.075 ;
        RECT 103.785 124.745 104.120 125.075 ;
        RECT 102.895 124.405 103.210 124.575 ;
        RECT 102.460 123.435 102.775 124.235 ;
        RECT 103.040 123.790 103.210 124.405 ;
        RECT 103.380 124.065 103.615 124.745 ;
        RECT 105.880 124.610 106.220 125.440 ;
        RECT 109.815 125.215 113.325 125.985 ;
        RECT 113.960 125.245 114.215 125.815 ;
        RECT 114.385 125.585 114.715 125.985 ;
        RECT 115.140 125.450 115.670 125.815 ;
        RECT 115.860 125.645 116.135 125.815 ;
        RECT 115.855 125.475 116.135 125.645 ;
        RECT 115.140 125.415 115.315 125.450 ;
        RECT 114.385 125.245 115.315 125.415 ;
        RECT 103.785 123.790 104.120 124.575 ;
        RECT 107.700 123.870 108.050 125.120 ;
        RECT 109.815 124.695 111.465 125.215 ;
        RECT 111.635 124.525 113.325 125.045 ;
        RECT 103.040 123.620 104.120 123.790 ;
        RECT 104.295 123.435 109.640 123.870 ;
        RECT 109.815 123.435 113.325 124.525 ;
        RECT 113.960 124.575 114.130 125.245 ;
        RECT 114.385 125.075 114.555 125.245 ;
        RECT 114.300 124.745 114.555 125.075 ;
        RECT 114.780 124.745 114.975 125.075 ;
        RECT 113.960 123.605 114.295 124.575 ;
        RECT 114.465 123.435 114.635 124.575 ;
        RECT 114.805 123.775 114.975 124.745 ;
        RECT 115.145 124.115 115.315 125.245 ;
        RECT 115.485 124.455 115.655 125.255 ;
        RECT 115.860 124.655 116.135 125.475 ;
        RECT 116.305 124.455 116.495 125.815 ;
        RECT 116.675 125.450 117.185 125.985 ;
        RECT 117.405 125.175 117.650 125.780 ;
        RECT 118.095 125.215 119.765 125.985 ;
        RECT 120.395 125.260 120.685 125.985 ;
        RECT 121.835 125.525 122.080 125.985 ;
        RECT 116.695 125.005 117.925 125.175 ;
        RECT 115.485 124.285 116.495 124.455 ;
        RECT 116.665 124.440 117.415 124.630 ;
        RECT 115.145 123.945 116.270 124.115 ;
        RECT 116.665 123.775 116.835 124.440 ;
        RECT 117.585 124.195 117.925 125.005 ;
        RECT 118.095 124.695 118.845 125.215 ;
        RECT 119.015 124.525 119.765 125.045 ;
        RECT 121.775 124.745 122.090 125.355 ;
        RECT 122.260 124.995 122.510 125.805 ;
        RECT 122.680 125.460 122.940 125.985 ;
        RECT 123.110 125.335 123.370 125.790 ;
        RECT 123.540 125.505 123.800 125.985 ;
        RECT 123.970 125.335 124.230 125.790 ;
        RECT 124.400 125.505 124.660 125.985 ;
        RECT 124.830 125.335 125.090 125.790 ;
        RECT 125.260 125.505 125.520 125.985 ;
        RECT 125.690 125.335 125.950 125.790 ;
        RECT 126.120 125.505 126.420 125.985 ;
        RECT 123.110 125.165 126.420 125.335 ;
        RECT 122.260 124.745 125.280 124.995 ;
        RECT 114.805 123.605 116.835 123.775 ;
        RECT 117.005 123.435 117.175 124.195 ;
        RECT 117.410 123.785 117.925 124.195 ;
        RECT 118.095 123.435 119.765 124.525 ;
        RECT 120.395 123.435 120.685 124.600 ;
        RECT 121.785 123.435 122.080 124.545 ;
        RECT 122.260 123.610 122.510 124.745 ;
        RECT 125.450 124.575 126.420 125.165 ;
        RECT 122.680 123.435 122.940 124.545 ;
        RECT 123.110 124.335 126.420 124.575 ;
        RECT 126.840 125.245 127.095 125.815 ;
        RECT 127.265 125.585 127.595 125.985 ;
        RECT 128.020 125.450 128.550 125.815 ;
        RECT 128.740 125.645 129.015 125.815 ;
        RECT 128.735 125.475 129.015 125.645 ;
        RECT 128.020 125.415 128.195 125.450 ;
        RECT 127.265 125.245 128.195 125.415 ;
        RECT 126.840 124.575 127.010 125.245 ;
        RECT 127.265 125.075 127.435 125.245 ;
        RECT 127.180 124.745 127.435 125.075 ;
        RECT 127.660 124.745 127.855 125.075 ;
        RECT 123.110 123.610 123.370 124.335 ;
        RECT 123.540 123.435 123.800 124.165 ;
        RECT 123.970 123.610 124.230 124.335 ;
        RECT 124.400 123.435 124.660 124.165 ;
        RECT 124.830 123.610 125.090 124.335 ;
        RECT 125.260 123.435 125.520 124.165 ;
        RECT 125.690 123.610 125.950 124.335 ;
        RECT 126.120 123.435 126.415 124.165 ;
        RECT 126.840 123.605 127.175 124.575 ;
        RECT 127.345 123.435 127.515 124.575 ;
        RECT 127.685 123.775 127.855 124.745 ;
        RECT 128.025 124.115 128.195 125.245 ;
        RECT 128.365 124.455 128.535 125.255 ;
        RECT 128.740 124.655 129.015 125.475 ;
        RECT 129.185 124.455 129.375 125.815 ;
        RECT 129.555 125.450 130.065 125.985 ;
        RECT 130.285 125.175 130.530 125.780 ;
        RECT 130.975 125.235 132.185 125.985 ;
        RECT 132.445 125.435 132.615 125.725 ;
        RECT 132.785 125.605 133.115 125.985 ;
        RECT 132.445 125.265 133.110 125.435 ;
        RECT 129.575 125.005 130.805 125.175 ;
        RECT 128.365 124.285 129.375 124.455 ;
        RECT 129.545 124.440 130.295 124.630 ;
        RECT 128.025 123.945 129.150 124.115 ;
        RECT 129.545 123.775 129.715 124.440 ;
        RECT 130.465 124.195 130.805 125.005 ;
        RECT 130.975 124.695 131.495 125.235 ;
        RECT 131.665 124.525 132.185 125.065 ;
        RECT 127.685 123.605 129.715 123.775 ;
        RECT 129.885 123.435 130.055 124.195 ;
        RECT 130.290 123.785 130.805 124.195 ;
        RECT 130.975 123.435 132.185 124.525 ;
        RECT 132.360 124.445 132.710 125.095 ;
        RECT 132.880 124.275 133.110 125.265 ;
        RECT 132.445 124.105 133.110 124.275 ;
        RECT 132.445 123.605 132.615 124.105 ;
        RECT 132.785 123.435 133.115 123.935 ;
        RECT 133.285 123.605 133.470 125.725 ;
        RECT 133.725 125.525 133.975 125.985 ;
        RECT 134.145 125.535 134.480 125.705 ;
        RECT 134.675 125.535 135.350 125.705 ;
        RECT 134.145 125.395 134.315 125.535 ;
        RECT 133.640 124.405 133.920 125.355 ;
        RECT 134.090 125.265 134.315 125.395 ;
        RECT 134.090 124.160 134.260 125.265 ;
        RECT 134.485 125.115 135.010 125.335 ;
        RECT 134.430 124.350 134.670 124.945 ;
        RECT 134.840 124.415 135.010 125.115 ;
        RECT 135.180 124.755 135.350 125.535 ;
        RECT 135.670 125.485 136.040 125.985 ;
        RECT 136.220 125.535 136.625 125.705 ;
        RECT 136.795 125.535 137.580 125.705 ;
        RECT 136.220 125.305 136.390 125.535 ;
        RECT 135.560 125.005 136.390 125.305 ;
        RECT 136.775 125.035 137.240 125.365 ;
        RECT 135.560 124.975 135.760 125.005 ;
        RECT 135.880 124.755 136.050 124.825 ;
        RECT 135.180 124.585 136.050 124.755 ;
        RECT 135.540 124.495 136.050 124.585 ;
        RECT 134.090 124.030 134.395 124.160 ;
        RECT 134.840 124.050 135.370 124.415 ;
        RECT 133.710 123.435 133.975 123.895 ;
        RECT 134.145 123.605 134.395 124.030 ;
        RECT 135.540 123.880 135.710 124.495 ;
        RECT 134.605 123.710 135.710 123.880 ;
        RECT 135.880 123.435 136.050 124.235 ;
        RECT 136.220 123.935 136.390 125.005 ;
        RECT 136.560 124.105 136.750 124.825 ;
        RECT 136.920 124.075 137.240 125.035 ;
        RECT 137.410 125.075 137.580 125.535 ;
        RECT 137.855 125.455 138.065 125.985 ;
        RECT 138.325 125.245 138.655 125.770 ;
        RECT 138.825 125.375 138.995 125.985 ;
        RECT 139.165 125.330 139.495 125.765 ;
        RECT 139.165 125.245 139.545 125.330 ;
        RECT 138.455 125.075 138.655 125.245 ;
        RECT 139.320 125.205 139.545 125.245 ;
        RECT 137.410 124.745 138.285 125.075 ;
        RECT 138.455 124.745 139.205 125.075 ;
        RECT 136.220 123.605 136.470 123.935 ;
        RECT 137.410 123.905 137.580 124.745 ;
        RECT 138.455 124.540 138.645 124.745 ;
        RECT 139.375 124.625 139.545 125.205 ;
        RECT 139.715 125.215 141.385 125.985 ;
        RECT 142.105 125.435 142.275 125.815 ;
        RECT 142.490 125.605 142.820 125.985 ;
        RECT 142.105 125.265 142.820 125.435 ;
        RECT 139.715 124.695 140.465 125.215 ;
        RECT 139.330 124.575 139.545 124.625 ;
        RECT 137.750 124.165 138.645 124.540 ;
        RECT 139.155 124.495 139.545 124.575 ;
        RECT 140.635 124.525 141.385 125.045 ;
        RECT 142.015 124.715 142.370 125.085 ;
        RECT 142.650 125.075 142.820 125.265 ;
        RECT 142.990 125.240 143.245 125.815 ;
        RECT 142.650 124.745 142.905 125.075 ;
        RECT 142.650 124.535 142.820 124.745 ;
        RECT 136.695 123.735 137.580 123.905 ;
        RECT 137.760 123.435 138.075 123.935 ;
        RECT 138.305 123.605 138.645 124.165 ;
        RECT 138.815 123.435 138.985 124.445 ;
        RECT 139.155 123.650 139.485 124.495 ;
        RECT 139.715 123.435 141.385 124.525 ;
        RECT 142.105 124.365 142.820 124.535 ;
        RECT 143.075 124.510 143.245 125.240 ;
        RECT 143.420 125.145 143.680 125.985 ;
        RECT 143.945 125.435 144.115 125.815 ;
        RECT 144.330 125.605 144.660 125.985 ;
        RECT 143.945 125.265 144.660 125.435 ;
        RECT 143.855 124.715 144.210 125.085 ;
        RECT 144.490 125.075 144.660 125.265 ;
        RECT 144.830 125.240 145.085 125.815 ;
        RECT 144.490 124.745 144.745 125.075 ;
        RECT 142.105 123.605 142.275 124.365 ;
        RECT 142.490 123.435 142.820 124.195 ;
        RECT 142.990 123.605 143.245 124.510 ;
        RECT 143.420 123.435 143.680 124.585 ;
        RECT 144.490 124.535 144.660 124.745 ;
        RECT 143.945 124.365 144.660 124.535 ;
        RECT 144.915 124.510 145.085 125.240 ;
        RECT 145.260 125.145 145.520 125.985 ;
        RECT 145.695 125.235 146.905 125.985 ;
        RECT 143.945 123.605 144.115 124.365 ;
        RECT 144.330 123.435 144.660 124.195 ;
        RECT 144.830 123.605 145.085 124.510 ;
        RECT 145.260 123.435 145.520 124.585 ;
        RECT 145.695 124.525 146.215 125.065 ;
        RECT 146.385 124.695 146.905 125.235 ;
        RECT 145.695 123.435 146.905 124.525 ;
        RECT 17.270 123.265 146.990 123.435 ;
        RECT 17.355 122.175 18.565 123.265 ;
        RECT 19.285 122.595 19.455 123.095 ;
        RECT 19.625 122.765 19.955 123.265 ;
        RECT 19.285 122.425 19.950 122.595 ;
        RECT 17.355 121.465 17.875 122.005 ;
        RECT 18.045 121.635 18.565 122.175 ;
        RECT 19.200 121.605 19.550 122.255 ;
        RECT 17.355 120.715 18.565 121.465 ;
        RECT 19.720 121.435 19.950 122.425 ;
        RECT 19.285 121.265 19.950 121.435 ;
        RECT 19.285 120.975 19.455 121.265 ;
        RECT 19.625 120.715 19.955 121.095 ;
        RECT 20.125 120.975 20.310 123.095 ;
        RECT 20.550 122.805 20.815 123.265 ;
        RECT 20.985 122.670 21.235 123.095 ;
        RECT 21.445 122.820 22.550 122.990 ;
        RECT 20.930 122.540 21.235 122.670 ;
        RECT 20.480 121.345 20.760 122.295 ;
        RECT 20.930 121.435 21.100 122.540 ;
        RECT 21.270 121.755 21.510 122.350 ;
        RECT 21.680 122.285 22.210 122.650 ;
        RECT 21.680 121.585 21.850 122.285 ;
        RECT 22.380 122.205 22.550 122.820 ;
        RECT 22.720 122.465 22.890 123.265 ;
        RECT 23.060 122.765 23.310 123.095 ;
        RECT 23.535 122.795 24.420 122.965 ;
        RECT 22.380 122.115 22.890 122.205 ;
        RECT 20.930 121.305 21.155 121.435 ;
        RECT 21.325 121.365 21.850 121.585 ;
        RECT 22.020 121.945 22.890 122.115 ;
        RECT 20.565 120.715 20.815 121.175 ;
        RECT 20.985 121.165 21.155 121.305 ;
        RECT 22.020 121.165 22.190 121.945 ;
        RECT 22.720 121.875 22.890 121.945 ;
        RECT 22.400 121.695 22.600 121.725 ;
        RECT 23.060 121.695 23.230 122.765 ;
        RECT 23.400 121.875 23.590 122.595 ;
        RECT 22.400 121.395 23.230 121.695 ;
        RECT 23.760 121.665 24.080 122.625 ;
        RECT 20.985 120.995 21.320 121.165 ;
        RECT 21.515 120.995 22.190 121.165 ;
        RECT 22.510 120.715 22.880 121.215 ;
        RECT 23.060 121.165 23.230 121.395 ;
        RECT 23.615 121.335 24.080 121.665 ;
        RECT 24.250 121.955 24.420 122.795 ;
        RECT 24.600 122.765 24.915 123.265 ;
        RECT 25.145 122.535 25.485 123.095 ;
        RECT 24.590 122.160 25.485 122.535 ;
        RECT 25.655 122.255 25.825 123.265 ;
        RECT 25.295 121.955 25.485 122.160 ;
        RECT 25.995 122.205 26.325 123.050 ;
        RECT 27.015 122.310 27.285 123.265 ;
        RECT 27.470 122.210 27.775 122.995 ;
        RECT 27.955 122.795 28.640 123.265 ;
        RECT 27.950 122.275 28.645 122.585 ;
        RECT 25.995 122.125 26.385 122.205 ;
        RECT 26.170 122.075 26.385 122.125 ;
        RECT 24.250 121.625 25.125 121.955 ;
        RECT 25.295 121.625 26.045 121.955 ;
        RECT 24.250 121.165 24.420 121.625 ;
        RECT 25.295 121.455 25.495 121.625 ;
        RECT 26.215 121.495 26.385 122.075 ;
        RECT 26.160 121.455 26.385 121.495 ;
        RECT 23.060 120.995 23.465 121.165 ;
        RECT 23.635 120.995 24.420 121.165 ;
        RECT 24.695 120.715 24.905 121.245 ;
        RECT 25.165 120.930 25.495 121.455 ;
        RECT 26.005 121.370 26.385 121.455 ;
        RECT 27.470 121.405 27.645 122.210 ;
        RECT 28.820 122.105 29.105 123.050 ;
        RECT 29.305 122.815 29.635 123.265 ;
        RECT 29.805 122.645 29.975 123.075 ;
        RECT 28.245 121.955 29.105 122.105 ;
        RECT 27.815 121.935 29.105 121.955 ;
        RECT 29.295 122.415 29.975 122.645 ;
        RECT 27.815 121.575 28.805 121.935 ;
        RECT 29.295 121.765 29.530 122.415 ;
        RECT 25.665 120.715 25.835 121.325 ;
        RECT 26.005 120.935 26.335 121.370 ;
        RECT 27.015 120.715 27.285 121.350 ;
        RECT 27.470 120.885 27.705 121.405 ;
        RECT 28.635 121.240 28.805 121.575 ;
        RECT 28.975 121.435 29.530 121.765 ;
        RECT 29.315 121.285 29.530 121.435 ;
        RECT 29.700 121.565 30.000 122.245 ;
        RECT 30.235 122.100 30.525 123.265 ;
        RECT 30.785 122.595 30.955 123.095 ;
        RECT 31.125 122.765 31.455 123.265 ;
        RECT 30.785 122.425 31.450 122.595 ;
        RECT 30.700 121.605 31.050 122.255 ;
        RECT 29.700 121.395 30.005 121.565 ;
        RECT 27.875 120.715 28.275 121.210 ;
        RECT 28.635 121.045 29.035 121.240 ;
        RECT 28.865 120.900 29.035 121.045 ;
        RECT 29.315 120.910 29.555 121.285 ;
        RECT 29.725 120.715 30.055 121.220 ;
        RECT 30.235 120.715 30.525 121.440 ;
        RECT 31.220 121.435 31.450 122.425 ;
        RECT 30.785 121.265 31.450 121.435 ;
        RECT 30.785 120.975 30.955 121.265 ;
        RECT 31.125 120.715 31.455 121.095 ;
        RECT 31.625 120.975 31.810 123.095 ;
        RECT 32.050 122.805 32.315 123.265 ;
        RECT 32.485 122.670 32.735 123.095 ;
        RECT 32.945 122.820 34.050 122.990 ;
        RECT 32.430 122.540 32.735 122.670 ;
        RECT 31.980 121.345 32.260 122.295 ;
        RECT 32.430 121.435 32.600 122.540 ;
        RECT 32.770 121.755 33.010 122.350 ;
        RECT 33.180 122.285 33.710 122.650 ;
        RECT 33.180 121.585 33.350 122.285 ;
        RECT 33.880 122.205 34.050 122.820 ;
        RECT 34.220 122.465 34.390 123.265 ;
        RECT 34.560 122.765 34.810 123.095 ;
        RECT 35.035 122.795 35.920 122.965 ;
        RECT 33.880 122.115 34.390 122.205 ;
        RECT 32.430 121.305 32.655 121.435 ;
        RECT 32.825 121.365 33.350 121.585 ;
        RECT 33.520 121.945 34.390 122.115 ;
        RECT 32.065 120.715 32.315 121.175 ;
        RECT 32.485 121.165 32.655 121.305 ;
        RECT 33.520 121.165 33.690 121.945 ;
        RECT 34.220 121.875 34.390 121.945 ;
        RECT 33.900 121.695 34.100 121.725 ;
        RECT 34.560 121.695 34.730 122.765 ;
        RECT 34.900 121.875 35.090 122.595 ;
        RECT 33.900 121.395 34.730 121.695 ;
        RECT 35.260 121.665 35.580 122.625 ;
        RECT 32.485 120.995 32.820 121.165 ;
        RECT 33.015 120.995 33.690 121.165 ;
        RECT 34.010 120.715 34.380 121.215 ;
        RECT 34.560 121.165 34.730 121.395 ;
        RECT 35.115 121.335 35.580 121.665 ;
        RECT 35.750 121.955 35.920 122.795 ;
        RECT 36.100 122.765 36.415 123.265 ;
        RECT 36.645 122.535 36.985 123.095 ;
        RECT 36.090 122.160 36.985 122.535 ;
        RECT 37.155 122.255 37.325 123.265 ;
        RECT 36.795 121.955 36.985 122.160 ;
        RECT 37.495 122.205 37.825 123.050 ;
        RECT 38.055 122.830 43.400 123.265 ;
        RECT 43.575 122.830 48.920 123.265 ;
        RECT 49.095 122.830 54.440 123.265 ;
        RECT 37.495 122.125 37.885 122.205 ;
        RECT 37.670 122.075 37.885 122.125 ;
        RECT 35.750 121.625 36.625 121.955 ;
        RECT 36.795 121.625 37.545 121.955 ;
        RECT 35.750 121.165 35.920 121.625 ;
        RECT 36.795 121.455 36.995 121.625 ;
        RECT 37.715 121.495 37.885 122.075 ;
        RECT 37.660 121.455 37.885 121.495 ;
        RECT 34.560 120.995 34.965 121.165 ;
        RECT 35.135 120.995 35.920 121.165 ;
        RECT 36.195 120.715 36.405 121.245 ;
        RECT 36.665 120.930 36.995 121.455 ;
        RECT 37.505 121.370 37.885 121.455 ;
        RECT 37.165 120.715 37.335 121.325 ;
        RECT 37.505 120.935 37.835 121.370 ;
        RECT 39.640 121.260 39.980 122.090 ;
        RECT 41.460 121.580 41.810 122.830 ;
        RECT 45.160 121.260 45.500 122.090 ;
        RECT 46.980 121.580 47.330 122.830 ;
        RECT 50.680 121.260 51.020 122.090 ;
        RECT 52.500 121.580 52.850 122.830 ;
        RECT 54.615 122.175 55.825 123.265 ;
        RECT 54.615 121.465 55.135 122.005 ;
        RECT 55.305 121.635 55.825 122.175 ;
        RECT 55.995 122.100 56.285 123.265 ;
        RECT 56.455 122.830 61.800 123.265 ;
        RECT 61.975 122.830 67.320 123.265 ;
        RECT 67.495 122.830 72.840 123.265 ;
        RECT 73.015 122.830 78.360 123.265 ;
        RECT 38.055 120.715 43.400 121.260 ;
        RECT 43.575 120.715 48.920 121.260 ;
        RECT 49.095 120.715 54.440 121.260 ;
        RECT 54.615 120.715 55.825 121.465 ;
        RECT 55.995 120.715 56.285 121.440 ;
        RECT 58.040 121.260 58.380 122.090 ;
        RECT 59.860 121.580 60.210 122.830 ;
        RECT 63.560 121.260 63.900 122.090 ;
        RECT 65.380 121.580 65.730 122.830 ;
        RECT 69.080 121.260 69.420 122.090 ;
        RECT 70.900 121.580 71.250 122.830 ;
        RECT 74.600 121.260 74.940 122.090 ;
        RECT 76.420 121.580 76.770 122.830 ;
        RECT 78.535 122.175 81.125 123.265 ;
        RECT 78.535 121.485 79.745 122.005 ;
        RECT 79.915 121.655 81.125 122.175 ;
        RECT 81.755 122.100 82.045 123.265 ;
        RECT 82.215 122.175 85.725 123.265 ;
        RECT 86.905 122.645 87.075 123.075 ;
        RECT 87.245 122.815 87.575 123.265 ;
        RECT 86.905 122.415 87.580 122.645 ;
        RECT 82.215 121.485 83.865 122.005 ;
        RECT 84.035 121.655 85.725 122.175 ;
        RECT 56.455 120.715 61.800 121.260 ;
        RECT 61.975 120.715 67.320 121.260 ;
        RECT 67.495 120.715 72.840 121.260 ;
        RECT 73.015 120.715 78.360 121.260 ;
        RECT 78.535 120.715 81.125 121.485 ;
        RECT 81.755 120.715 82.045 121.440 ;
        RECT 82.215 120.715 85.725 121.485 ;
        RECT 86.875 121.395 87.175 122.245 ;
        RECT 87.345 121.765 87.580 122.415 ;
        RECT 87.750 122.105 88.035 123.050 ;
        RECT 88.215 122.795 88.900 123.265 ;
        RECT 88.210 122.275 88.905 122.585 ;
        RECT 89.080 122.210 89.385 122.995 ;
        RECT 87.750 121.955 88.610 122.105 ;
        RECT 87.750 121.935 89.035 121.955 ;
        RECT 87.345 121.435 87.880 121.765 ;
        RECT 88.050 121.575 89.035 121.935 ;
        RECT 87.345 121.285 87.565 121.435 ;
        RECT 86.820 120.715 87.155 121.220 ;
        RECT 87.325 120.910 87.565 121.285 ;
        RECT 88.050 121.240 88.220 121.575 ;
        RECT 89.210 121.405 89.385 122.210 ;
        RECT 90.165 122.095 90.495 123.265 ;
        RECT 90.695 121.925 91.025 123.095 ;
        RECT 91.225 122.095 91.555 123.265 ;
        RECT 91.755 121.925 92.115 123.095 ;
        RECT 92.285 122.125 92.615 123.265 ;
        RECT 93.345 122.595 93.515 123.095 ;
        RECT 93.685 122.765 94.015 123.265 ;
        RECT 93.345 122.425 94.010 122.595 ;
        RECT 90.695 121.645 92.115 121.925 ;
        RECT 87.845 121.045 88.220 121.240 ;
        RECT 87.845 120.900 88.015 121.045 ;
        RECT 88.580 120.715 88.975 121.210 ;
        RECT 89.145 120.885 89.385 121.405 ;
        RECT 90.705 120.715 91.035 121.405 ;
        RECT 91.755 121.310 92.115 121.645 ;
        RECT 92.285 121.375 92.625 121.955 ;
        RECT 93.260 121.605 93.610 122.255 ;
        RECT 93.780 121.435 94.010 122.425 ;
        RECT 91.495 120.885 92.115 121.310 ;
        RECT 93.345 121.265 94.010 121.435 ;
        RECT 92.285 120.715 92.615 121.205 ;
        RECT 93.345 120.975 93.515 121.265 ;
        RECT 93.685 120.715 94.015 121.095 ;
        RECT 94.185 120.975 94.370 123.095 ;
        RECT 94.610 122.805 94.875 123.265 ;
        RECT 95.045 122.670 95.295 123.095 ;
        RECT 95.505 122.820 96.610 122.990 ;
        RECT 94.990 122.540 95.295 122.670 ;
        RECT 94.540 121.345 94.820 122.295 ;
        RECT 94.990 121.435 95.160 122.540 ;
        RECT 95.330 121.755 95.570 122.350 ;
        RECT 95.740 122.285 96.270 122.650 ;
        RECT 95.740 121.585 95.910 122.285 ;
        RECT 96.440 122.205 96.610 122.820 ;
        RECT 96.780 122.465 96.950 123.265 ;
        RECT 97.120 122.765 97.370 123.095 ;
        RECT 97.595 122.795 98.480 122.965 ;
        RECT 96.440 122.115 96.950 122.205 ;
        RECT 94.990 121.305 95.215 121.435 ;
        RECT 95.385 121.365 95.910 121.585 ;
        RECT 96.080 121.945 96.950 122.115 ;
        RECT 94.625 120.715 94.875 121.175 ;
        RECT 95.045 121.165 95.215 121.305 ;
        RECT 96.080 121.165 96.250 121.945 ;
        RECT 96.780 121.875 96.950 121.945 ;
        RECT 96.460 121.695 96.660 121.725 ;
        RECT 97.120 121.695 97.290 122.765 ;
        RECT 97.460 121.875 97.650 122.595 ;
        RECT 96.460 121.395 97.290 121.695 ;
        RECT 97.820 121.665 98.140 122.625 ;
        RECT 95.045 120.995 95.380 121.165 ;
        RECT 95.575 120.995 96.250 121.165 ;
        RECT 96.570 120.715 96.940 121.215 ;
        RECT 97.120 121.165 97.290 121.395 ;
        RECT 97.675 121.335 98.140 121.665 ;
        RECT 98.310 121.955 98.480 122.795 ;
        RECT 98.660 122.765 98.975 123.265 ;
        RECT 99.205 122.535 99.545 123.095 ;
        RECT 98.650 122.160 99.545 122.535 ;
        RECT 99.715 122.255 99.885 123.265 ;
        RECT 99.355 121.955 99.545 122.160 ;
        RECT 100.055 122.205 100.385 123.050 ;
        RECT 100.055 122.125 100.445 122.205 ;
        RECT 100.665 122.170 100.915 123.265 ;
        RECT 101.650 122.925 103.715 123.095 ;
        RECT 100.230 122.075 100.445 122.125 ;
        RECT 101.085 122.085 101.440 122.500 ;
        RECT 101.650 122.085 101.895 122.925 ;
        RECT 98.310 121.625 99.185 121.955 ;
        RECT 99.355 121.625 100.105 121.955 ;
        RECT 98.310 121.165 98.480 121.625 ;
        RECT 99.355 121.455 99.555 121.625 ;
        RECT 100.275 121.495 100.445 122.075 ;
        RECT 101.270 121.915 101.440 122.085 ;
        RECT 100.615 121.705 101.100 121.915 ;
        RECT 101.270 121.705 101.895 121.915 ;
        RECT 101.270 121.535 101.440 121.705 ;
        RECT 102.065 121.535 102.315 122.755 ;
        RECT 102.485 122.085 102.755 122.925 ;
        RECT 103.045 122.255 103.295 122.755 ;
        RECT 103.465 122.425 103.715 122.925 ;
        RECT 103.885 122.255 104.135 123.095 ;
        RECT 104.305 122.425 104.555 123.265 ;
        RECT 104.725 122.255 105.040 123.095 ;
        RECT 105.220 122.840 105.555 123.265 ;
        RECT 105.725 122.660 105.910 123.065 ;
        RECT 103.045 122.085 105.040 122.255 ;
        RECT 105.245 122.485 105.910 122.660 ;
        RECT 106.115 122.485 106.445 123.265 ;
        RECT 102.490 121.705 103.995 121.915 ;
        RECT 104.165 121.705 105.020 121.915 ;
        RECT 100.220 121.455 100.445 121.495 ;
        RECT 97.120 120.995 97.525 121.165 ;
        RECT 97.695 120.995 98.480 121.165 ;
        RECT 98.755 120.715 98.965 121.245 ;
        RECT 99.225 120.930 99.555 121.455 ;
        RECT 100.065 121.370 100.445 121.455 ;
        RECT 99.725 120.715 99.895 121.325 ;
        RECT 100.065 120.935 100.395 121.370 ;
        RECT 100.625 120.715 100.915 121.455 ;
        RECT 101.085 121.010 101.440 121.535 ;
        RECT 101.650 120.715 101.855 121.525 ;
        RECT 102.025 121.355 104.595 121.535 ;
        RECT 102.025 120.885 102.355 121.355 ;
        RECT 102.525 120.715 103.255 121.185 ;
        RECT 103.425 120.885 103.755 121.355 ;
        RECT 103.925 120.715 104.095 121.185 ;
        RECT 104.265 120.885 104.595 121.355 ;
        RECT 104.765 120.715 105.040 121.535 ;
        RECT 105.245 121.455 105.585 122.485 ;
        RECT 106.615 122.295 106.885 123.065 ;
        RECT 105.755 122.125 106.885 122.295 ;
        RECT 105.755 121.625 106.005 122.125 ;
        RECT 105.245 121.285 105.930 121.455 ;
        RECT 106.185 121.375 106.545 121.955 ;
        RECT 105.220 120.715 105.555 121.115 ;
        RECT 105.725 120.885 105.930 121.285 ;
        RECT 106.715 121.215 106.885 122.125 ;
        RECT 107.515 122.100 107.805 123.265 ;
        RECT 107.980 122.315 108.245 123.085 ;
        RECT 108.415 122.545 108.745 123.265 ;
        RECT 108.935 122.725 109.195 123.085 ;
        RECT 109.365 122.895 109.695 123.265 ;
        RECT 109.865 122.725 110.125 123.085 ;
        RECT 108.935 122.495 110.125 122.725 ;
        RECT 110.695 122.315 110.985 123.085 ;
        RECT 106.140 120.715 106.415 121.195 ;
        RECT 106.625 120.885 106.885 121.215 ;
        RECT 107.515 120.715 107.805 121.440 ;
        RECT 107.980 120.895 108.315 122.315 ;
        RECT 108.490 122.135 110.985 122.315 ;
        RECT 111.195 122.175 112.865 123.265 ;
        RECT 113.585 122.595 113.755 123.095 ;
        RECT 113.925 122.765 114.255 123.265 ;
        RECT 113.585 122.425 114.250 122.595 ;
        RECT 108.490 121.445 108.715 122.135 ;
        RECT 108.915 121.625 109.195 121.955 ;
        RECT 109.375 121.625 109.950 121.955 ;
        RECT 110.130 121.625 110.565 121.955 ;
        RECT 110.745 121.625 111.015 121.955 ;
        RECT 111.195 121.485 111.945 122.005 ;
        RECT 112.115 121.655 112.865 122.175 ;
        RECT 113.500 121.605 113.850 122.255 ;
        RECT 108.490 121.255 110.975 121.445 ;
        RECT 108.495 120.715 109.240 121.085 ;
        RECT 109.805 120.895 110.060 121.255 ;
        RECT 110.240 120.715 110.570 121.085 ;
        RECT 110.750 120.895 110.975 121.255 ;
        RECT 111.195 120.715 112.865 121.485 ;
        RECT 114.020 121.435 114.250 122.425 ;
        RECT 113.585 121.265 114.250 121.435 ;
        RECT 113.585 120.975 113.755 121.265 ;
        RECT 113.925 120.715 114.255 121.095 ;
        RECT 114.425 120.975 114.610 123.095 ;
        RECT 114.850 122.805 115.115 123.265 ;
        RECT 115.285 122.670 115.535 123.095 ;
        RECT 115.745 122.820 116.850 122.990 ;
        RECT 115.230 122.540 115.535 122.670 ;
        RECT 114.780 121.345 115.060 122.295 ;
        RECT 115.230 121.435 115.400 122.540 ;
        RECT 115.570 121.755 115.810 122.350 ;
        RECT 115.980 122.285 116.510 122.650 ;
        RECT 115.980 121.585 116.150 122.285 ;
        RECT 116.680 122.205 116.850 122.820 ;
        RECT 117.020 122.465 117.190 123.265 ;
        RECT 117.360 122.765 117.610 123.095 ;
        RECT 117.835 122.795 118.720 122.965 ;
        RECT 116.680 122.115 117.190 122.205 ;
        RECT 115.230 121.305 115.455 121.435 ;
        RECT 115.625 121.365 116.150 121.585 ;
        RECT 116.320 121.945 117.190 122.115 ;
        RECT 114.865 120.715 115.115 121.175 ;
        RECT 115.285 121.165 115.455 121.305 ;
        RECT 116.320 121.165 116.490 121.945 ;
        RECT 117.020 121.875 117.190 121.945 ;
        RECT 116.700 121.695 116.900 121.725 ;
        RECT 117.360 121.695 117.530 122.765 ;
        RECT 117.700 121.875 117.890 122.595 ;
        RECT 116.700 121.395 117.530 121.695 ;
        RECT 118.060 121.665 118.380 122.625 ;
        RECT 115.285 120.995 115.620 121.165 ;
        RECT 115.815 120.995 116.490 121.165 ;
        RECT 116.810 120.715 117.180 121.215 ;
        RECT 117.360 121.165 117.530 121.395 ;
        RECT 117.915 121.335 118.380 121.665 ;
        RECT 118.550 121.955 118.720 122.795 ;
        RECT 118.900 122.765 119.215 123.265 ;
        RECT 119.445 122.535 119.785 123.095 ;
        RECT 118.890 122.160 119.785 122.535 ;
        RECT 119.955 122.255 120.125 123.265 ;
        RECT 119.595 121.955 119.785 122.160 ;
        RECT 120.295 122.205 120.625 123.050 ;
        RECT 120.295 122.125 120.685 122.205 ;
        RECT 120.865 122.155 121.160 123.265 ;
        RECT 120.470 122.075 120.685 122.125 ;
        RECT 118.550 121.625 119.425 121.955 ;
        RECT 119.595 121.625 120.345 121.955 ;
        RECT 118.550 121.165 118.720 121.625 ;
        RECT 119.595 121.455 119.795 121.625 ;
        RECT 120.515 121.495 120.685 122.075 ;
        RECT 121.340 121.955 121.590 123.090 ;
        RECT 121.760 122.155 122.020 123.265 ;
        RECT 122.190 122.365 122.450 123.090 ;
        RECT 122.620 122.535 122.880 123.265 ;
        RECT 123.050 122.365 123.310 123.090 ;
        RECT 123.480 122.535 123.740 123.265 ;
        RECT 123.910 122.365 124.170 123.090 ;
        RECT 124.340 122.535 124.600 123.265 ;
        RECT 124.770 122.365 125.030 123.090 ;
        RECT 125.200 122.535 125.495 123.265 ;
        RECT 122.190 122.125 125.500 122.365 ;
        RECT 125.915 122.175 129.425 123.265 ;
        RECT 120.460 121.455 120.685 121.495 ;
        RECT 117.360 120.995 117.765 121.165 ;
        RECT 117.935 120.995 118.720 121.165 ;
        RECT 118.995 120.715 119.205 121.245 ;
        RECT 119.465 120.930 119.795 121.455 ;
        RECT 120.305 121.370 120.685 121.455 ;
        RECT 119.965 120.715 120.135 121.325 ;
        RECT 120.305 120.935 120.635 121.370 ;
        RECT 120.855 121.345 121.170 121.955 ;
        RECT 121.340 121.705 124.360 121.955 ;
        RECT 120.915 120.715 121.160 121.175 ;
        RECT 121.340 120.895 121.590 121.705 ;
        RECT 124.530 121.535 125.500 122.125 ;
        RECT 122.190 121.365 125.500 121.535 ;
        RECT 125.915 121.485 127.565 122.005 ;
        RECT 127.735 121.655 129.425 122.175 ;
        RECT 129.685 122.255 129.855 123.095 ;
        RECT 130.025 122.925 131.195 123.095 ;
        RECT 130.025 122.425 130.355 122.925 ;
        RECT 130.865 122.885 131.195 122.925 ;
        RECT 131.385 122.845 131.740 123.265 ;
        RECT 130.525 122.665 130.755 122.755 ;
        RECT 131.910 122.665 132.160 123.095 ;
        RECT 130.525 122.425 132.160 122.665 ;
        RECT 132.330 122.505 132.660 123.265 ;
        RECT 132.830 122.425 133.085 123.095 ;
        RECT 129.685 122.085 132.745 122.255 ;
        RECT 129.600 121.705 129.950 121.915 ;
        RECT 130.120 121.705 130.565 121.905 ;
        RECT 130.735 121.705 131.210 121.905 ;
        RECT 121.760 120.715 122.020 121.240 ;
        RECT 122.190 120.910 122.450 121.365 ;
        RECT 122.620 120.715 122.880 121.195 ;
        RECT 123.050 120.910 123.310 121.365 ;
        RECT 123.480 120.715 123.740 121.195 ;
        RECT 123.910 120.910 124.170 121.365 ;
        RECT 124.340 120.715 124.600 121.195 ;
        RECT 124.770 120.910 125.030 121.365 ;
        RECT 125.200 120.715 125.500 121.195 ;
        RECT 125.915 120.715 129.425 121.485 ;
        RECT 129.685 121.365 130.750 121.535 ;
        RECT 129.685 120.885 129.855 121.365 ;
        RECT 130.025 120.715 130.355 121.195 ;
        RECT 130.580 121.135 130.750 121.365 ;
        RECT 130.930 121.305 131.210 121.705 ;
        RECT 131.480 121.705 131.810 121.905 ;
        RECT 131.980 121.705 132.345 121.905 ;
        RECT 131.480 121.305 131.765 121.705 ;
        RECT 132.575 121.535 132.745 122.085 ;
        RECT 131.945 121.365 132.745 121.535 ;
        RECT 131.945 121.135 132.115 121.365 ;
        RECT 132.915 121.295 133.085 122.425 ;
        RECT 133.275 122.100 133.565 123.265 ;
        RECT 133.740 122.125 134.075 123.095 ;
        RECT 134.245 122.125 134.415 123.265 ;
        RECT 134.585 122.925 136.615 123.095 ;
        RECT 133.740 121.455 133.910 122.125 ;
        RECT 134.585 121.955 134.755 122.925 ;
        RECT 134.080 121.625 134.335 121.955 ;
        RECT 134.560 121.625 134.755 121.955 ;
        RECT 134.925 122.585 136.050 122.755 ;
        RECT 134.165 121.455 134.335 121.625 ;
        RECT 134.925 121.455 135.095 122.585 ;
        RECT 132.900 121.215 133.085 121.295 ;
        RECT 130.580 120.885 132.115 121.135 ;
        RECT 132.285 120.715 132.615 121.195 ;
        RECT 132.830 120.885 133.085 121.215 ;
        RECT 133.275 120.715 133.565 121.440 ;
        RECT 133.740 120.885 133.995 121.455 ;
        RECT 134.165 121.285 135.095 121.455 ;
        RECT 135.265 122.245 136.275 122.415 ;
        RECT 135.265 121.445 135.435 122.245 ;
        RECT 135.640 121.905 135.915 122.045 ;
        RECT 135.635 121.735 135.915 121.905 ;
        RECT 134.920 121.250 135.095 121.285 ;
        RECT 134.165 120.715 134.495 121.115 ;
        RECT 134.920 120.885 135.450 121.250 ;
        RECT 135.640 120.885 135.915 121.735 ;
        RECT 136.085 120.885 136.275 122.245 ;
        RECT 136.445 122.260 136.615 122.925 ;
        RECT 136.785 122.505 136.955 123.265 ;
        RECT 137.190 122.505 137.705 122.915 ;
        RECT 136.445 122.070 137.195 122.260 ;
        RECT 137.365 121.695 137.705 122.505 ;
        RECT 137.875 122.175 141.385 123.265 ;
        RECT 136.475 121.525 137.705 121.695 ;
        RECT 136.455 120.715 136.965 121.250 ;
        RECT 137.185 120.920 137.430 121.525 ;
        RECT 137.875 121.485 139.525 122.005 ;
        RECT 139.695 121.655 141.385 122.175 ;
        RECT 142.105 122.335 142.275 123.095 ;
        RECT 142.490 122.505 142.820 123.265 ;
        RECT 142.105 122.165 142.820 122.335 ;
        RECT 142.990 122.190 143.245 123.095 ;
        RECT 142.015 121.615 142.370 121.985 ;
        RECT 142.650 121.955 142.820 122.165 ;
        RECT 142.650 121.625 142.905 121.955 ;
        RECT 137.875 120.715 141.385 121.485 ;
        RECT 142.650 121.435 142.820 121.625 ;
        RECT 143.075 121.460 143.245 122.190 ;
        RECT 143.420 122.115 143.680 123.265 ;
        RECT 143.945 122.335 144.115 123.095 ;
        RECT 144.330 122.505 144.660 123.265 ;
        RECT 143.945 122.165 144.660 122.335 ;
        RECT 144.830 122.190 145.085 123.095 ;
        RECT 143.855 121.615 144.210 121.985 ;
        RECT 144.490 121.955 144.660 122.165 ;
        RECT 144.490 121.625 144.745 121.955 ;
        RECT 142.105 121.265 142.820 121.435 ;
        RECT 142.105 120.885 142.275 121.265 ;
        RECT 142.490 120.715 142.820 121.095 ;
        RECT 142.990 120.885 143.245 121.460 ;
        RECT 143.420 120.715 143.680 121.555 ;
        RECT 144.490 121.435 144.660 121.625 ;
        RECT 144.915 121.460 145.085 122.190 ;
        RECT 145.260 122.115 145.520 123.265 ;
        RECT 145.695 122.175 146.905 123.265 ;
        RECT 145.695 121.635 146.215 122.175 ;
        RECT 143.945 121.265 144.660 121.435 ;
        RECT 143.945 120.885 144.115 121.265 ;
        RECT 144.330 120.715 144.660 121.095 ;
        RECT 144.830 120.885 145.085 121.460 ;
        RECT 145.260 120.715 145.520 121.555 ;
        RECT 146.385 121.465 146.905 122.005 ;
        RECT 145.695 120.715 146.905 121.465 ;
        RECT 17.270 120.545 146.990 120.715 ;
        RECT 17.355 119.795 18.565 120.545 ;
        RECT 18.825 119.995 18.995 120.375 ;
        RECT 19.175 120.165 19.505 120.545 ;
        RECT 18.825 119.825 19.490 119.995 ;
        RECT 19.685 119.870 19.945 120.375 ;
        RECT 17.355 119.255 17.875 119.795 ;
        RECT 18.045 119.085 18.565 119.625 ;
        RECT 18.755 119.275 19.095 119.645 ;
        RECT 19.320 119.570 19.490 119.825 ;
        RECT 19.320 119.240 19.595 119.570 ;
        RECT 19.320 119.095 19.490 119.240 ;
        RECT 17.355 117.995 18.565 119.085 ;
        RECT 18.815 118.925 19.490 119.095 ;
        RECT 19.765 119.070 19.945 119.870 ;
        RECT 20.205 119.995 20.375 120.375 ;
        RECT 20.555 120.165 20.885 120.545 ;
        RECT 20.205 119.825 20.870 119.995 ;
        RECT 21.065 119.870 21.325 120.375 ;
        RECT 20.135 119.275 20.475 119.645 ;
        RECT 20.700 119.570 20.870 119.825 ;
        RECT 20.700 119.240 20.975 119.570 ;
        RECT 20.700 119.095 20.870 119.240 ;
        RECT 18.815 118.165 18.995 118.925 ;
        RECT 19.175 117.995 19.505 118.755 ;
        RECT 19.675 118.165 19.945 119.070 ;
        RECT 20.195 118.925 20.870 119.095 ;
        RECT 21.145 119.070 21.325 119.870 ;
        RECT 20.195 118.165 20.375 118.925 ;
        RECT 20.555 117.995 20.885 118.755 ;
        RECT 21.055 118.165 21.325 119.070 ;
        RECT 21.500 119.805 21.755 120.375 ;
        RECT 21.925 120.145 22.255 120.545 ;
        RECT 22.680 120.010 23.210 120.375 ;
        RECT 23.400 120.205 23.675 120.375 ;
        RECT 23.395 120.035 23.675 120.205 ;
        RECT 22.680 119.975 22.855 120.010 ;
        RECT 21.925 119.805 22.855 119.975 ;
        RECT 21.500 119.135 21.670 119.805 ;
        RECT 21.925 119.635 22.095 119.805 ;
        RECT 21.840 119.305 22.095 119.635 ;
        RECT 22.320 119.305 22.515 119.635 ;
        RECT 21.500 118.165 21.835 119.135 ;
        RECT 22.005 117.995 22.175 119.135 ;
        RECT 22.345 118.335 22.515 119.305 ;
        RECT 22.685 118.675 22.855 119.805 ;
        RECT 23.025 119.015 23.195 119.815 ;
        RECT 23.400 119.215 23.675 120.035 ;
        RECT 23.845 119.015 24.035 120.375 ;
        RECT 24.215 120.010 24.725 120.545 ;
        RECT 24.945 119.735 25.190 120.340 ;
        RECT 26.185 119.995 26.355 120.285 ;
        RECT 26.525 120.165 26.855 120.545 ;
        RECT 26.185 119.825 26.850 119.995 ;
        RECT 24.235 119.565 25.465 119.735 ;
        RECT 23.025 118.845 24.035 119.015 ;
        RECT 24.205 119.000 24.955 119.190 ;
        RECT 22.685 118.505 23.810 118.675 ;
        RECT 24.205 118.335 24.375 119.000 ;
        RECT 25.125 118.755 25.465 119.565 ;
        RECT 26.100 119.005 26.450 119.655 ;
        RECT 26.620 118.835 26.850 119.825 ;
        RECT 22.345 118.165 24.375 118.335 ;
        RECT 24.545 117.995 24.715 118.755 ;
        RECT 24.950 118.345 25.465 118.755 ;
        RECT 26.185 118.665 26.850 118.835 ;
        RECT 26.185 118.165 26.355 118.665 ;
        RECT 26.525 117.995 26.855 118.495 ;
        RECT 27.025 118.165 27.210 120.285 ;
        RECT 27.465 120.085 27.715 120.545 ;
        RECT 27.885 120.095 28.220 120.265 ;
        RECT 28.415 120.095 29.090 120.265 ;
        RECT 27.885 119.955 28.055 120.095 ;
        RECT 27.380 118.965 27.660 119.915 ;
        RECT 27.830 119.825 28.055 119.955 ;
        RECT 27.830 118.720 28.000 119.825 ;
        RECT 28.225 119.675 28.750 119.895 ;
        RECT 28.170 118.910 28.410 119.505 ;
        RECT 28.580 118.975 28.750 119.675 ;
        RECT 28.920 119.315 29.090 120.095 ;
        RECT 29.410 120.045 29.780 120.545 ;
        RECT 29.960 120.095 30.365 120.265 ;
        RECT 30.535 120.095 31.320 120.265 ;
        RECT 29.960 119.865 30.130 120.095 ;
        RECT 29.300 119.565 30.130 119.865 ;
        RECT 30.515 119.595 30.980 119.925 ;
        RECT 29.300 119.535 29.500 119.565 ;
        RECT 29.620 119.315 29.790 119.385 ;
        RECT 28.920 119.145 29.790 119.315 ;
        RECT 29.280 119.055 29.790 119.145 ;
        RECT 27.830 118.590 28.135 118.720 ;
        RECT 28.580 118.610 29.110 118.975 ;
        RECT 27.450 117.995 27.715 118.455 ;
        RECT 27.885 118.165 28.135 118.590 ;
        RECT 29.280 118.440 29.450 119.055 ;
        RECT 28.345 118.270 29.450 118.440 ;
        RECT 29.620 117.995 29.790 118.795 ;
        RECT 29.960 118.495 30.130 119.565 ;
        RECT 30.300 118.665 30.490 119.385 ;
        RECT 30.660 118.635 30.980 119.595 ;
        RECT 31.150 119.635 31.320 120.095 ;
        RECT 31.595 120.015 31.805 120.545 ;
        RECT 32.065 119.805 32.395 120.330 ;
        RECT 32.565 119.935 32.735 120.545 ;
        RECT 32.905 119.890 33.235 120.325 ;
        RECT 33.465 120.040 33.795 120.545 ;
        RECT 33.965 119.975 34.205 120.350 ;
        RECT 34.485 120.215 34.655 120.360 ;
        RECT 34.485 120.020 34.885 120.215 ;
        RECT 35.245 120.050 35.645 120.545 ;
        RECT 32.905 119.805 33.285 119.890 ;
        RECT 32.195 119.635 32.395 119.805 ;
        RECT 33.060 119.765 33.285 119.805 ;
        RECT 31.150 119.305 32.025 119.635 ;
        RECT 32.195 119.305 32.945 119.635 ;
        RECT 29.960 118.165 30.210 118.495 ;
        RECT 31.150 118.465 31.320 119.305 ;
        RECT 32.195 119.100 32.385 119.305 ;
        RECT 33.115 119.185 33.285 119.765 ;
        RECT 33.515 119.695 33.820 119.865 ;
        RECT 33.070 119.135 33.285 119.185 ;
        RECT 31.490 118.725 32.385 119.100 ;
        RECT 32.895 119.055 33.285 119.135 ;
        RECT 30.435 118.295 31.320 118.465 ;
        RECT 31.500 117.995 31.815 118.495 ;
        RECT 32.045 118.165 32.385 118.725 ;
        RECT 32.555 117.995 32.725 119.005 ;
        RECT 32.895 118.210 33.225 119.055 ;
        RECT 33.520 119.015 33.820 119.695 ;
        RECT 33.990 119.825 34.205 119.975 ;
        RECT 33.990 119.495 34.545 119.825 ;
        RECT 34.715 119.685 34.885 120.020 ;
        RECT 35.815 119.855 36.050 120.375 ;
        RECT 36.235 119.910 36.505 120.545 ;
        RECT 36.675 120.000 42.020 120.545 ;
        RECT 33.990 118.845 34.225 119.495 ;
        RECT 34.715 119.325 35.705 119.685 ;
        RECT 33.545 118.615 34.225 118.845 ;
        RECT 34.415 119.305 35.705 119.325 ;
        RECT 34.415 119.155 35.275 119.305 ;
        RECT 33.545 118.185 33.715 118.615 ;
        RECT 33.885 117.995 34.215 118.445 ;
        RECT 34.415 118.210 34.700 119.155 ;
        RECT 35.875 119.050 36.050 119.855 ;
        RECT 38.260 119.170 38.600 120.000 ;
        RECT 43.115 119.820 43.405 120.545 ;
        RECT 43.575 120.000 48.920 120.545 ;
        RECT 49.095 120.000 54.440 120.545 ;
        RECT 54.615 120.000 59.960 120.545 ;
        RECT 60.135 120.000 65.480 120.545 ;
        RECT 34.875 118.675 35.570 118.985 ;
        RECT 34.880 117.995 35.565 118.465 ;
        RECT 35.745 118.265 36.050 119.050 ;
        RECT 36.235 117.995 36.505 118.950 ;
        RECT 40.080 118.430 40.430 119.680 ;
        RECT 45.160 119.170 45.500 120.000 ;
        RECT 36.675 117.995 42.020 118.430 ;
        RECT 43.115 117.995 43.405 119.160 ;
        RECT 46.980 118.430 47.330 119.680 ;
        RECT 50.680 119.170 51.020 120.000 ;
        RECT 52.500 118.430 52.850 119.680 ;
        RECT 56.200 119.170 56.540 120.000 ;
        RECT 58.020 118.430 58.370 119.680 ;
        RECT 61.720 119.170 62.060 120.000 ;
        RECT 65.655 119.775 68.245 120.545 ;
        RECT 68.875 119.820 69.165 120.545 ;
        RECT 69.335 119.775 72.845 120.545 ;
        RECT 73.940 120.040 74.275 120.545 ;
        RECT 74.445 119.975 74.685 120.350 ;
        RECT 74.965 120.215 75.135 120.360 ;
        RECT 74.965 120.020 75.340 120.215 ;
        RECT 75.700 120.050 76.095 120.545 ;
        RECT 63.540 118.430 63.890 119.680 ;
        RECT 65.655 119.255 66.865 119.775 ;
        RECT 67.035 119.085 68.245 119.605 ;
        RECT 69.335 119.255 70.985 119.775 ;
        RECT 43.575 117.995 48.920 118.430 ;
        RECT 49.095 117.995 54.440 118.430 ;
        RECT 54.615 117.995 59.960 118.430 ;
        RECT 60.135 117.995 65.480 118.430 ;
        RECT 65.655 117.995 68.245 119.085 ;
        RECT 68.875 117.995 69.165 119.160 ;
        RECT 71.155 119.085 72.845 119.605 ;
        RECT 69.335 117.995 72.845 119.085 ;
        RECT 73.995 119.015 74.295 119.865 ;
        RECT 74.465 119.825 74.685 119.975 ;
        RECT 74.465 119.495 75.000 119.825 ;
        RECT 75.170 119.685 75.340 120.020 ;
        RECT 76.265 119.855 76.505 120.375 ;
        RECT 74.465 118.845 74.700 119.495 ;
        RECT 75.170 119.325 76.155 119.685 ;
        RECT 74.025 118.615 74.700 118.845 ;
        RECT 74.870 119.305 76.155 119.325 ;
        RECT 74.870 119.155 75.730 119.305 ;
        RECT 74.025 118.185 74.195 118.615 ;
        RECT 74.365 117.995 74.695 118.445 ;
        RECT 74.870 118.210 75.155 119.155 ;
        RECT 76.330 119.050 76.505 119.855 ;
        RECT 76.695 119.795 77.905 120.545 ;
        RECT 78.080 119.805 78.335 120.375 ;
        RECT 78.505 120.145 78.835 120.545 ;
        RECT 79.260 120.010 79.790 120.375 ;
        RECT 79.980 120.205 80.255 120.375 ;
        RECT 79.975 120.035 80.255 120.205 ;
        RECT 79.260 119.975 79.435 120.010 ;
        RECT 78.505 119.805 79.435 119.975 ;
        RECT 76.695 119.255 77.215 119.795 ;
        RECT 77.385 119.085 77.905 119.625 ;
        RECT 75.330 118.675 76.025 118.985 ;
        RECT 75.335 117.995 76.020 118.465 ;
        RECT 76.200 118.265 76.505 119.050 ;
        RECT 76.695 117.995 77.905 119.085 ;
        RECT 78.080 119.135 78.250 119.805 ;
        RECT 78.505 119.635 78.675 119.805 ;
        RECT 78.420 119.305 78.675 119.635 ;
        RECT 78.900 119.305 79.095 119.635 ;
        RECT 78.080 118.165 78.415 119.135 ;
        RECT 78.585 117.995 78.755 119.135 ;
        RECT 78.925 118.335 79.095 119.305 ;
        RECT 79.265 118.675 79.435 119.805 ;
        RECT 79.605 119.015 79.775 119.815 ;
        RECT 79.980 119.215 80.255 120.035 ;
        RECT 80.425 119.015 80.615 120.375 ;
        RECT 80.795 120.010 81.305 120.545 ;
        RECT 81.525 119.735 81.770 120.340 ;
        RECT 82.215 119.775 83.885 120.545 ;
        RECT 84.520 119.805 84.775 120.375 ;
        RECT 84.945 120.145 85.275 120.545 ;
        RECT 85.700 120.010 86.230 120.375 ;
        RECT 86.420 120.205 86.695 120.375 ;
        RECT 86.415 120.035 86.695 120.205 ;
        RECT 85.700 119.975 85.875 120.010 ;
        RECT 84.945 119.805 85.875 119.975 ;
        RECT 80.815 119.565 82.045 119.735 ;
        RECT 79.605 118.845 80.615 119.015 ;
        RECT 80.785 119.000 81.535 119.190 ;
        RECT 79.265 118.505 80.390 118.675 ;
        RECT 80.785 118.335 80.955 119.000 ;
        RECT 81.705 118.755 82.045 119.565 ;
        RECT 82.215 119.255 82.965 119.775 ;
        RECT 83.135 119.085 83.885 119.605 ;
        RECT 78.925 118.165 80.955 118.335 ;
        RECT 81.125 117.995 81.295 118.755 ;
        RECT 81.530 118.345 82.045 118.755 ;
        RECT 82.215 117.995 83.885 119.085 ;
        RECT 84.520 119.135 84.690 119.805 ;
        RECT 84.945 119.635 85.115 119.805 ;
        RECT 84.860 119.305 85.115 119.635 ;
        RECT 85.340 119.305 85.535 119.635 ;
        RECT 84.520 118.165 84.855 119.135 ;
        RECT 85.025 117.995 85.195 119.135 ;
        RECT 85.365 118.335 85.535 119.305 ;
        RECT 85.705 118.675 85.875 119.805 ;
        RECT 86.045 119.015 86.215 119.815 ;
        RECT 86.420 119.215 86.695 120.035 ;
        RECT 86.865 119.015 87.055 120.375 ;
        RECT 87.235 120.010 87.745 120.545 ;
        RECT 87.965 119.735 88.210 120.340 ;
        RECT 88.655 119.775 90.325 120.545 ;
        RECT 90.500 119.915 90.835 120.375 ;
        RECT 91.005 120.085 91.175 120.545 ;
        RECT 91.345 119.915 91.675 120.375 ;
        RECT 91.845 120.085 92.015 120.545 ;
        RECT 92.185 120.165 94.195 120.375 ;
        RECT 92.185 119.915 92.435 120.165 ;
        RECT 87.255 119.565 88.485 119.735 ;
        RECT 86.045 118.845 87.055 119.015 ;
        RECT 87.225 119.000 87.975 119.190 ;
        RECT 85.705 118.505 86.830 118.675 ;
        RECT 87.225 118.335 87.395 119.000 ;
        RECT 88.145 118.755 88.485 119.565 ;
        RECT 88.655 119.255 89.405 119.775 ;
        RECT 90.500 119.725 92.435 119.915 ;
        RECT 92.605 119.825 93.775 119.995 ;
        RECT 89.575 119.085 90.325 119.605 ;
        RECT 92.605 119.555 92.855 119.825 ;
        RECT 93.945 119.745 94.195 120.165 ;
        RECT 94.635 119.820 94.925 120.545 ;
        RECT 96.020 119.705 96.280 120.545 ;
        RECT 96.455 119.800 96.710 120.375 ;
        RECT 96.880 120.165 97.210 120.545 ;
        RECT 97.425 119.995 97.595 120.375 ;
        RECT 96.880 119.825 97.595 119.995 ;
        RECT 90.520 119.305 92.140 119.555 ;
        RECT 92.320 119.135 92.855 119.555 ;
        RECT 93.025 119.305 94.465 119.555 ;
        RECT 85.365 118.165 87.395 118.335 ;
        RECT 87.565 117.995 87.735 118.755 ;
        RECT 87.970 118.345 88.485 118.755 ;
        RECT 88.655 117.995 90.325 119.085 ;
        RECT 90.500 117.995 90.755 119.135 ;
        RECT 90.925 118.965 93.775 119.135 ;
        RECT 90.925 118.165 91.255 118.965 ;
        RECT 91.425 117.995 91.595 118.795 ;
        RECT 91.765 118.165 92.095 118.965 ;
        RECT 92.265 117.995 92.435 118.795 ;
        RECT 92.605 118.165 92.935 118.965 ;
        RECT 93.105 117.995 93.275 118.795 ;
        RECT 93.445 118.165 93.775 118.965 ;
        RECT 93.945 117.995 94.195 118.795 ;
        RECT 94.635 117.995 94.925 119.160 ;
        RECT 96.020 117.995 96.280 119.145 ;
        RECT 96.455 119.070 96.625 119.800 ;
        RECT 96.880 119.635 97.050 119.825 ;
        RECT 97.860 119.725 98.135 120.545 ;
        RECT 98.305 119.905 98.635 120.375 ;
        RECT 98.805 120.075 98.975 120.545 ;
        RECT 99.145 119.905 99.475 120.375 ;
        RECT 99.645 120.075 100.375 120.545 ;
        RECT 100.545 119.905 100.875 120.375 ;
        RECT 98.305 119.725 100.875 119.905 ;
        RECT 101.045 119.735 101.250 120.545 ;
        RECT 101.460 119.725 101.815 120.250 ;
        RECT 101.985 119.805 102.275 120.545 ;
        RECT 102.520 120.275 103.005 120.375 ;
        RECT 102.520 120.085 103.970 120.275 ;
        RECT 104.150 120.185 104.480 120.545 ;
        RECT 105.015 120.185 105.345 120.545 ;
        RECT 102.520 119.825 103.005 120.085 ;
        RECT 103.790 120.015 103.970 120.085 ;
        RECT 104.655 120.015 104.845 120.115 ;
        RECT 105.515 120.015 105.705 120.375 ;
        RECT 105.875 120.185 106.205 120.545 ;
        RECT 100.585 119.695 100.845 119.725 ;
        RECT 96.795 119.305 97.050 119.635 ;
        RECT 96.880 119.095 97.050 119.305 ;
        RECT 97.330 119.275 97.685 119.645 ;
        RECT 97.880 119.345 98.735 119.555 ;
        RECT 98.905 119.345 100.410 119.555 ;
        RECT 96.455 118.165 96.710 119.070 ;
        RECT 96.880 118.925 97.595 119.095 ;
        RECT 96.880 117.995 97.210 118.755 ;
        RECT 97.425 118.165 97.595 118.925 ;
        RECT 97.860 119.005 99.855 119.175 ;
        RECT 97.860 118.165 98.175 119.005 ;
        RECT 98.345 117.995 98.595 118.835 ;
        RECT 98.765 118.165 99.015 119.005 ;
        RECT 99.185 118.335 99.435 118.835 ;
        RECT 99.605 118.505 99.855 119.005 ;
        RECT 100.145 118.335 100.415 119.175 ;
        RECT 100.585 118.505 100.835 119.695 ;
        RECT 101.460 119.555 101.630 119.725 ;
        RECT 101.005 119.345 101.630 119.555 ;
        RECT 101.800 119.345 102.285 119.555 ;
        RECT 101.460 119.175 101.630 119.345 ;
        RECT 101.005 118.335 101.250 119.175 ;
        RECT 101.460 118.760 101.815 119.175 ;
        RECT 102.520 119.135 102.740 119.825 ;
        RECT 102.910 119.305 103.220 119.635 ;
        RECT 99.185 118.165 101.250 118.335 ;
        RECT 101.985 117.995 102.235 119.090 ;
        RECT 102.520 118.465 102.880 119.135 ;
        RECT 103.050 118.755 103.220 119.305 ;
        RECT 103.390 119.290 103.605 119.905 ;
        RECT 103.790 119.825 104.485 120.015 ;
        RECT 103.895 119.290 104.085 119.635 ;
        RECT 104.255 119.610 104.485 119.825 ;
        RECT 104.655 119.785 105.905 120.015 ;
        RECT 104.255 119.275 105.470 119.610 ;
        RECT 104.255 119.105 104.425 119.275 ;
        RECT 103.650 118.935 104.425 119.105 ;
        RECT 105.640 119.095 105.905 119.785 ;
        RECT 104.595 118.925 105.905 119.095 ;
        RECT 106.085 118.925 106.365 120.015 ;
        RECT 106.535 118.755 106.815 120.205 ;
        RECT 107.790 119.735 108.035 120.340 ;
        RECT 108.255 120.010 108.765 120.545 ;
        RECT 103.050 118.525 106.815 118.755 ;
        RECT 107.515 119.565 108.745 119.735 ;
        RECT 107.515 118.755 107.855 119.565 ;
        RECT 108.025 119.000 108.775 119.190 ;
        RECT 103.100 117.995 103.550 118.355 ;
        RECT 104.115 117.995 104.445 118.355 ;
        RECT 105.015 117.995 105.350 118.355 ;
        RECT 105.875 117.995 106.205 118.355 ;
        RECT 107.515 118.345 108.030 118.755 ;
        RECT 108.265 117.995 108.435 118.755 ;
        RECT 108.605 118.335 108.775 119.000 ;
        RECT 108.945 119.015 109.135 120.375 ;
        RECT 109.305 120.205 109.580 120.375 ;
        RECT 109.305 120.035 109.585 120.205 ;
        RECT 109.305 119.215 109.580 120.035 ;
        RECT 109.770 120.010 110.300 120.375 ;
        RECT 110.725 120.145 111.055 120.545 ;
        RECT 110.125 119.975 110.300 120.010 ;
        RECT 109.785 119.015 109.955 119.815 ;
        RECT 108.945 118.845 109.955 119.015 ;
        RECT 110.125 119.805 111.055 119.975 ;
        RECT 111.225 119.805 111.480 120.375 ;
        RECT 112.580 120.040 112.915 120.545 ;
        RECT 113.085 119.975 113.325 120.350 ;
        RECT 113.605 120.215 113.775 120.360 ;
        RECT 113.605 120.020 113.980 120.215 ;
        RECT 114.340 120.050 114.735 120.545 ;
        RECT 110.125 118.675 110.295 119.805 ;
        RECT 110.885 119.635 111.055 119.805 ;
        RECT 109.170 118.505 110.295 118.675 ;
        RECT 110.465 119.305 110.660 119.635 ;
        RECT 110.885 119.305 111.140 119.635 ;
        RECT 110.465 118.335 110.635 119.305 ;
        RECT 111.310 119.135 111.480 119.805 ;
        RECT 108.605 118.165 110.635 118.335 ;
        RECT 110.805 117.995 110.975 119.135 ;
        RECT 111.145 118.165 111.480 119.135 ;
        RECT 112.635 119.015 112.935 119.865 ;
        RECT 113.105 119.825 113.325 119.975 ;
        RECT 113.105 119.495 113.640 119.825 ;
        RECT 113.810 119.685 113.980 120.020 ;
        RECT 114.905 119.855 115.145 120.375 ;
        RECT 113.105 118.845 113.340 119.495 ;
        RECT 113.810 119.325 114.795 119.685 ;
        RECT 112.665 118.615 113.340 118.845 ;
        RECT 113.510 119.305 114.795 119.325 ;
        RECT 113.510 119.155 114.370 119.305 ;
        RECT 112.665 118.185 112.835 118.615 ;
        RECT 113.005 117.995 113.335 118.445 ;
        RECT 113.510 118.210 113.795 119.155 ;
        RECT 114.970 119.050 115.145 119.855 ;
        RECT 115.335 119.775 118.845 120.545 ;
        RECT 119.015 119.795 120.225 120.545 ;
        RECT 120.395 119.820 120.685 120.545 ;
        RECT 121.405 119.995 121.575 120.285 ;
        RECT 121.745 120.165 122.075 120.545 ;
        RECT 121.405 119.825 122.070 119.995 ;
        RECT 115.335 119.255 116.985 119.775 ;
        RECT 117.155 119.085 118.845 119.605 ;
        RECT 119.015 119.255 119.535 119.795 ;
        RECT 119.705 119.085 120.225 119.625 ;
        RECT 113.970 118.675 114.665 118.985 ;
        RECT 113.975 117.995 114.660 118.465 ;
        RECT 114.840 118.265 115.145 119.050 ;
        RECT 115.335 117.995 118.845 119.085 ;
        RECT 119.015 117.995 120.225 119.085 ;
        RECT 120.395 117.995 120.685 119.160 ;
        RECT 121.320 119.005 121.670 119.655 ;
        RECT 121.840 118.835 122.070 119.825 ;
        RECT 121.405 118.665 122.070 118.835 ;
        RECT 121.405 118.165 121.575 118.665 ;
        RECT 121.745 117.995 122.075 118.495 ;
        RECT 122.245 118.165 122.430 120.285 ;
        RECT 122.685 120.085 122.935 120.545 ;
        RECT 123.105 120.095 123.440 120.265 ;
        RECT 123.635 120.095 124.310 120.265 ;
        RECT 123.105 119.955 123.275 120.095 ;
        RECT 122.600 118.965 122.880 119.915 ;
        RECT 123.050 119.825 123.275 119.955 ;
        RECT 123.050 118.720 123.220 119.825 ;
        RECT 123.445 119.675 123.970 119.895 ;
        RECT 123.390 118.910 123.630 119.505 ;
        RECT 123.800 118.975 123.970 119.675 ;
        RECT 124.140 119.315 124.310 120.095 ;
        RECT 124.630 120.045 125.000 120.545 ;
        RECT 125.180 120.095 125.585 120.265 ;
        RECT 125.755 120.095 126.540 120.265 ;
        RECT 125.180 119.865 125.350 120.095 ;
        RECT 124.520 119.565 125.350 119.865 ;
        RECT 125.735 119.595 126.200 119.925 ;
        RECT 124.520 119.535 124.720 119.565 ;
        RECT 124.840 119.315 125.010 119.385 ;
        RECT 124.140 119.145 125.010 119.315 ;
        RECT 124.500 119.055 125.010 119.145 ;
        RECT 123.050 118.590 123.355 118.720 ;
        RECT 123.800 118.610 124.330 118.975 ;
        RECT 122.670 117.995 122.935 118.455 ;
        RECT 123.105 118.165 123.355 118.590 ;
        RECT 124.500 118.440 124.670 119.055 ;
        RECT 123.565 118.270 124.670 118.440 ;
        RECT 124.840 117.995 125.010 118.795 ;
        RECT 125.180 118.495 125.350 119.565 ;
        RECT 125.520 118.665 125.710 119.385 ;
        RECT 125.880 118.635 126.200 119.595 ;
        RECT 126.370 119.635 126.540 120.095 ;
        RECT 126.815 120.015 127.025 120.545 ;
        RECT 127.285 119.805 127.615 120.330 ;
        RECT 127.785 119.935 127.955 120.545 ;
        RECT 128.125 119.890 128.455 120.325 ;
        RECT 128.125 119.805 128.505 119.890 ;
        RECT 127.415 119.635 127.615 119.805 ;
        RECT 128.280 119.765 128.505 119.805 ;
        RECT 126.370 119.305 127.245 119.635 ;
        RECT 127.415 119.305 128.165 119.635 ;
        RECT 125.180 118.165 125.430 118.495 ;
        RECT 126.370 118.465 126.540 119.305 ;
        RECT 127.415 119.100 127.605 119.305 ;
        RECT 128.335 119.185 128.505 119.765 ;
        RECT 128.290 119.135 128.505 119.185 ;
        RECT 126.710 118.725 127.605 119.100 ;
        RECT 128.115 119.055 128.505 119.135 ;
        RECT 128.680 119.805 128.935 120.375 ;
        RECT 129.105 120.145 129.435 120.545 ;
        RECT 129.860 120.010 130.390 120.375 ;
        RECT 129.860 119.975 130.035 120.010 ;
        RECT 129.105 119.805 130.035 119.975 ;
        RECT 128.680 119.135 128.850 119.805 ;
        RECT 129.105 119.635 129.275 119.805 ;
        RECT 129.020 119.305 129.275 119.635 ;
        RECT 129.500 119.305 129.695 119.635 ;
        RECT 125.655 118.295 126.540 118.465 ;
        RECT 126.720 117.995 127.035 118.495 ;
        RECT 127.265 118.165 127.605 118.725 ;
        RECT 127.775 117.995 127.945 119.005 ;
        RECT 128.115 118.210 128.445 119.055 ;
        RECT 128.680 118.165 129.015 119.135 ;
        RECT 129.185 117.995 129.355 119.135 ;
        RECT 129.525 118.335 129.695 119.305 ;
        RECT 129.865 118.675 130.035 119.805 ;
        RECT 130.205 119.015 130.375 119.815 ;
        RECT 130.580 119.525 130.855 120.375 ;
        RECT 130.575 119.355 130.855 119.525 ;
        RECT 130.580 119.215 130.855 119.355 ;
        RECT 131.025 119.015 131.215 120.375 ;
        RECT 131.395 120.010 131.905 120.545 ;
        RECT 132.125 119.735 132.370 120.340 ;
        RECT 132.815 119.775 134.485 120.545 ;
        RECT 134.660 120.040 134.995 120.545 ;
        RECT 135.165 119.975 135.405 120.350 ;
        RECT 135.685 120.215 135.855 120.360 ;
        RECT 135.685 120.020 136.060 120.215 ;
        RECT 136.420 120.050 136.815 120.545 ;
        RECT 131.415 119.565 132.645 119.735 ;
        RECT 130.205 118.845 131.215 119.015 ;
        RECT 131.385 119.000 132.135 119.190 ;
        RECT 129.865 118.505 130.990 118.675 ;
        RECT 131.385 118.335 131.555 119.000 ;
        RECT 132.305 118.755 132.645 119.565 ;
        RECT 132.815 119.255 133.565 119.775 ;
        RECT 133.735 119.085 134.485 119.605 ;
        RECT 129.525 118.165 131.555 118.335 ;
        RECT 131.725 117.995 131.895 118.755 ;
        RECT 132.130 118.345 132.645 118.755 ;
        RECT 132.815 117.995 134.485 119.085 ;
        RECT 134.715 119.015 135.015 119.865 ;
        RECT 135.185 119.825 135.405 119.975 ;
        RECT 135.185 119.495 135.720 119.825 ;
        RECT 135.890 119.685 136.060 120.020 ;
        RECT 136.985 119.855 137.225 120.375 ;
        RECT 135.185 118.845 135.420 119.495 ;
        RECT 135.890 119.325 136.875 119.685 ;
        RECT 134.745 118.615 135.420 118.845 ;
        RECT 135.590 119.305 136.875 119.325 ;
        RECT 135.590 119.155 136.450 119.305 ;
        RECT 134.745 118.185 134.915 118.615 ;
        RECT 135.085 117.995 135.415 118.445 ;
        RECT 135.590 118.210 135.875 119.155 ;
        RECT 137.050 119.050 137.225 119.855 ;
        RECT 137.505 119.995 137.675 120.285 ;
        RECT 137.845 120.165 138.175 120.545 ;
        RECT 137.505 119.825 138.170 119.995 ;
        RECT 136.050 118.675 136.745 118.985 ;
        RECT 136.055 117.995 136.740 118.465 ;
        RECT 136.920 118.265 137.225 119.050 ;
        RECT 137.420 119.005 137.770 119.655 ;
        RECT 137.940 118.835 138.170 119.825 ;
        RECT 137.505 118.665 138.170 118.835 ;
        RECT 137.505 118.165 137.675 118.665 ;
        RECT 137.845 117.995 138.175 118.495 ;
        RECT 138.345 118.165 138.530 120.285 ;
        RECT 138.785 120.085 139.035 120.545 ;
        RECT 139.205 120.095 139.540 120.265 ;
        RECT 139.735 120.095 140.410 120.265 ;
        RECT 139.205 119.955 139.375 120.095 ;
        RECT 138.700 118.965 138.980 119.915 ;
        RECT 139.150 119.825 139.375 119.955 ;
        RECT 139.150 118.720 139.320 119.825 ;
        RECT 139.545 119.675 140.070 119.895 ;
        RECT 139.490 118.910 139.730 119.505 ;
        RECT 139.900 118.975 140.070 119.675 ;
        RECT 140.240 119.315 140.410 120.095 ;
        RECT 140.730 120.045 141.100 120.545 ;
        RECT 141.280 120.095 141.685 120.265 ;
        RECT 141.855 120.095 142.640 120.265 ;
        RECT 141.280 119.865 141.450 120.095 ;
        RECT 140.620 119.565 141.450 119.865 ;
        RECT 141.835 119.595 142.300 119.925 ;
        RECT 140.620 119.535 140.820 119.565 ;
        RECT 140.940 119.315 141.110 119.385 ;
        RECT 140.240 119.145 141.110 119.315 ;
        RECT 140.600 119.055 141.110 119.145 ;
        RECT 139.150 118.590 139.455 118.720 ;
        RECT 139.900 118.610 140.430 118.975 ;
        RECT 138.770 117.995 139.035 118.455 ;
        RECT 139.205 118.165 139.455 118.590 ;
        RECT 140.600 118.440 140.770 119.055 ;
        RECT 139.665 118.270 140.770 118.440 ;
        RECT 140.940 117.995 141.110 118.795 ;
        RECT 141.280 118.495 141.450 119.565 ;
        RECT 141.620 118.665 141.810 119.385 ;
        RECT 141.980 118.635 142.300 119.595 ;
        RECT 142.470 119.635 142.640 120.095 ;
        RECT 142.915 120.015 143.125 120.545 ;
        RECT 143.385 119.805 143.715 120.330 ;
        RECT 143.885 119.935 144.055 120.545 ;
        RECT 144.225 119.890 144.555 120.325 ;
        RECT 144.225 119.805 144.605 119.890 ;
        RECT 143.515 119.635 143.715 119.805 ;
        RECT 144.380 119.765 144.605 119.805 ;
        RECT 145.695 119.795 146.905 120.545 ;
        RECT 142.470 119.305 143.345 119.635 ;
        RECT 143.515 119.305 144.265 119.635 ;
        RECT 141.280 118.165 141.530 118.495 ;
        RECT 142.470 118.465 142.640 119.305 ;
        RECT 143.515 119.100 143.705 119.305 ;
        RECT 144.435 119.185 144.605 119.765 ;
        RECT 144.390 119.135 144.605 119.185 ;
        RECT 142.810 118.725 143.705 119.100 ;
        RECT 144.215 119.055 144.605 119.135 ;
        RECT 145.695 119.085 146.215 119.625 ;
        RECT 146.385 119.255 146.905 119.795 ;
        RECT 141.755 118.295 142.640 118.465 ;
        RECT 142.820 117.995 143.135 118.495 ;
        RECT 143.365 118.165 143.705 118.725 ;
        RECT 143.875 117.995 144.045 119.005 ;
        RECT 144.215 118.210 144.545 119.055 ;
        RECT 145.695 117.995 146.905 119.085 ;
        RECT 17.270 117.825 146.990 117.995 ;
        RECT 17.355 116.735 18.565 117.825 ;
        RECT 18.735 117.390 24.080 117.825 ;
        RECT 17.355 116.025 17.875 116.565 ;
        RECT 18.045 116.195 18.565 116.735 ;
        RECT 17.355 115.275 18.565 116.025 ;
        RECT 20.320 115.820 20.660 116.650 ;
        RECT 22.140 116.140 22.490 117.390 ;
        RECT 24.255 116.735 27.765 117.825 ;
        RECT 24.255 116.045 25.905 116.565 ;
        RECT 26.075 116.215 27.765 116.735 ;
        RECT 28.865 116.685 29.195 117.825 ;
        RECT 29.725 116.855 30.055 117.640 ;
        RECT 29.375 116.685 30.055 116.855 ;
        RECT 28.855 116.265 29.205 116.515 ;
        RECT 29.375 116.085 29.545 116.685 ;
        RECT 30.235 116.660 30.525 117.825 ;
        RECT 30.695 117.390 36.040 117.825 ;
        RECT 36.215 117.390 41.560 117.825 ;
        RECT 41.735 117.390 47.080 117.825 ;
        RECT 47.255 117.390 52.600 117.825 ;
        RECT 29.715 116.265 30.065 116.515 ;
        RECT 18.735 115.275 24.080 115.820 ;
        RECT 24.255 115.275 27.765 116.045 ;
        RECT 28.865 115.275 29.135 116.085 ;
        RECT 29.305 115.445 29.635 116.085 ;
        RECT 29.805 115.275 30.045 116.085 ;
        RECT 30.235 115.275 30.525 116.000 ;
        RECT 32.280 115.820 32.620 116.650 ;
        RECT 34.100 116.140 34.450 117.390 ;
        RECT 37.800 115.820 38.140 116.650 ;
        RECT 39.620 116.140 39.970 117.390 ;
        RECT 43.320 115.820 43.660 116.650 ;
        RECT 45.140 116.140 45.490 117.390 ;
        RECT 48.840 115.820 49.180 116.650 ;
        RECT 50.660 116.140 51.010 117.390 ;
        RECT 52.775 116.735 55.365 117.825 ;
        RECT 52.775 116.045 53.985 116.565 ;
        RECT 54.155 116.215 55.365 116.735 ;
        RECT 55.995 116.660 56.285 117.825 ;
        RECT 56.455 117.390 61.800 117.825 ;
        RECT 61.975 117.390 67.320 117.825 ;
        RECT 30.695 115.275 36.040 115.820 ;
        RECT 36.215 115.275 41.560 115.820 ;
        RECT 41.735 115.275 47.080 115.820 ;
        RECT 47.255 115.275 52.600 115.820 ;
        RECT 52.775 115.275 55.365 116.045 ;
        RECT 55.995 115.275 56.285 116.000 ;
        RECT 58.040 115.820 58.380 116.650 ;
        RECT 59.860 116.140 60.210 117.390 ;
        RECT 63.560 115.820 63.900 116.650 ;
        RECT 65.380 116.140 65.730 117.390 ;
        RECT 67.495 116.735 71.005 117.825 ;
        RECT 71.265 117.205 71.435 117.635 ;
        RECT 71.605 117.375 71.935 117.825 ;
        RECT 71.265 116.975 71.940 117.205 ;
        RECT 67.495 116.045 69.145 116.565 ;
        RECT 69.315 116.215 71.005 116.735 ;
        RECT 56.455 115.275 61.800 115.820 ;
        RECT 61.975 115.275 67.320 115.820 ;
        RECT 67.495 115.275 71.005 116.045 ;
        RECT 71.235 115.955 71.535 116.805 ;
        RECT 71.705 116.325 71.940 116.975 ;
        RECT 72.110 116.665 72.395 117.610 ;
        RECT 72.575 117.355 73.260 117.825 ;
        RECT 72.570 116.835 73.265 117.145 ;
        RECT 73.440 116.770 73.745 117.555 ;
        RECT 74.025 117.155 74.195 117.655 ;
        RECT 74.365 117.325 74.695 117.825 ;
        RECT 74.025 116.985 74.690 117.155 ;
        RECT 72.110 116.515 72.970 116.665 ;
        RECT 72.110 116.495 73.395 116.515 ;
        RECT 71.705 115.995 72.240 116.325 ;
        RECT 72.410 116.135 73.395 116.495 ;
        RECT 71.705 115.845 71.925 115.995 ;
        RECT 71.180 115.275 71.515 115.780 ;
        RECT 71.685 115.470 71.925 115.845 ;
        RECT 72.410 115.800 72.580 116.135 ;
        RECT 73.570 115.965 73.745 116.770 ;
        RECT 73.940 116.165 74.290 116.815 ;
        RECT 74.460 115.995 74.690 116.985 ;
        RECT 72.205 115.605 72.580 115.800 ;
        RECT 72.205 115.460 72.375 115.605 ;
        RECT 72.940 115.275 73.335 115.770 ;
        RECT 73.505 115.445 73.745 115.965 ;
        RECT 74.025 115.825 74.690 115.995 ;
        RECT 74.025 115.535 74.195 115.825 ;
        RECT 74.365 115.275 74.695 115.655 ;
        RECT 74.865 115.535 75.050 117.655 ;
        RECT 75.290 117.365 75.555 117.825 ;
        RECT 75.725 117.230 75.975 117.655 ;
        RECT 76.185 117.380 77.290 117.550 ;
        RECT 75.670 117.100 75.975 117.230 ;
        RECT 75.220 115.905 75.500 116.855 ;
        RECT 75.670 115.995 75.840 117.100 ;
        RECT 76.010 116.315 76.250 116.910 ;
        RECT 76.420 116.845 76.950 117.210 ;
        RECT 76.420 116.145 76.590 116.845 ;
        RECT 77.120 116.765 77.290 117.380 ;
        RECT 77.460 117.025 77.630 117.825 ;
        RECT 77.800 117.325 78.050 117.655 ;
        RECT 78.275 117.355 79.160 117.525 ;
        RECT 77.120 116.675 77.630 116.765 ;
        RECT 75.670 115.865 75.895 115.995 ;
        RECT 76.065 115.925 76.590 116.145 ;
        RECT 76.760 116.505 77.630 116.675 ;
        RECT 75.305 115.275 75.555 115.735 ;
        RECT 75.725 115.725 75.895 115.865 ;
        RECT 76.760 115.725 76.930 116.505 ;
        RECT 77.460 116.435 77.630 116.505 ;
        RECT 77.140 116.255 77.340 116.285 ;
        RECT 77.800 116.255 77.970 117.325 ;
        RECT 78.140 116.435 78.330 117.155 ;
        RECT 77.140 115.955 77.970 116.255 ;
        RECT 78.500 116.225 78.820 117.185 ;
        RECT 75.725 115.555 76.060 115.725 ;
        RECT 76.255 115.555 76.930 115.725 ;
        RECT 77.250 115.275 77.620 115.775 ;
        RECT 77.800 115.725 77.970 115.955 ;
        RECT 78.355 115.895 78.820 116.225 ;
        RECT 78.990 116.515 79.160 117.355 ;
        RECT 79.340 117.325 79.655 117.825 ;
        RECT 79.885 117.095 80.225 117.655 ;
        RECT 79.330 116.720 80.225 117.095 ;
        RECT 80.395 116.815 80.565 117.825 ;
        RECT 80.035 116.515 80.225 116.720 ;
        RECT 80.735 116.765 81.065 117.610 ;
        RECT 80.735 116.685 81.125 116.765 ;
        RECT 80.910 116.635 81.125 116.685 ;
        RECT 81.755 116.660 82.045 117.825 ;
        RECT 82.305 117.155 82.475 117.655 ;
        RECT 82.645 117.325 82.975 117.825 ;
        RECT 82.305 116.985 82.970 117.155 ;
        RECT 78.990 116.185 79.865 116.515 ;
        RECT 80.035 116.185 80.785 116.515 ;
        RECT 78.990 115.725 79.160 116.185 ;
        RECT 80.035 116.015 80.235 116.185 ;
        RECT 80.955 116.055 81.125 116.635 ;
        RECT 82.220 116.165 82.570 116.815 ;
        RECT 80.900 116.015 81.125 116.055 ;
        RECT 77.800 115.555 78.205 115.725 ;
        RECT 78.375 115.555 79.160 115.725 ;
        RECT 79.435 115.275 79.645 115.805 ;
        RECT 79.905 115.490 80.235 116.015 ;
        RECT 80.745 115.930 81.125 116.015 ;
        RECT 80.405 115.275 80.575 115.885 ;
        RECT 80.745 115.495 81.075 115.930 ;
        RECT 81.755 115.275 82.045 116.000 ;
        RECT 82.740 115.995 82.970 116.985 ;
        RECT 82.305 115.825 82.970 115.995 ;
        RECT 82.305 115.535 82.475 115.825 ;
        RECT 82.645 115.275 82.975 115.655 ;
        RECT 83.145 115.535 83.330 117.655 ;
        RECT 83.570 117.365 83.835 117.825 ;
        RECT 84.005 117.230 84.255 117.655 ;
        RECT 84.465 117.380 85.570 117.550 ;
        RECT 83.950 117.100 84.255 117.230 ;
        RECT 83.500 115.905 83.780 116.855 ;
        RECT 83.950 115.995 84.120 117.100 ;
        RECT 84.290 116.315 84.530 116.910 ;
        RECT 84.700 116.845 85.230 117.210 ;
        RECT 84.700 116.145 84.870 116.845 ;
        RECT 85.400 116.765 85.570 117.380 ;
        RECT 85.740 117.025 85.910 117.825 ;
        RECT 86.080 117.325 86.330 117.655 ;
        RECT 86.555 117.355 87.440 117.525 ;
        RECT 85.400 116.675 85.910 116.765 ;
        RECT 83.950 115.865 84.175 115.995 ;
        RECT 84.345 115.925 84.870 116.145 ;
        RECT 85.040 116.505 85.910 116.675 ;
        RECT 83.585 115.275 83.835 115.735 ;
        RECT 84.005 115.725 84.175 115.865 ;
        RECT 85.040 115.725 85.210 116.505 ;
        RECT 85.740 116.435 85.910 116.505 ;
        RECT 85.420 116.255 85.620 116.285 ;
        RECT 86.080 116.255 86.250 117.325 ;
        RECT 86.420 116.435 86.610 117.155 ;
        RECT 85.420 115.955 86.250 116.255 ;
        RECT 86.780 116.225 87.100 117.185 ;
        RECT 84.005 115.555 84.340 115.725 ;
        RECT 84.535 115.555 85.210 115.725 ;
        RECT 85.530 115.275 85.900 115.775 ;
        RECT 86.080 115.725 86.250 115.955 ;
        RECT 86.635 115.895 87.100 116.225 ;
        RECT 87.270 116.515 87.440 117.355 ;
        RECT 87.620 117.325 87.935 117.825 ;
        RECT 88.165 117.095 88.505 117.655 ;
        RECT 87.610 116.720 88.505 117.095 ;
        RECT 88.675 116.815 88.845 117.825 ;
        RECT 88.315 116.515 88.505 116.720 ;
        RECT 89.015 116.765 89.345 117.610 ;
        RECT 89.015 116.685 89.405 116.765 ;
        RECT 89.190 116.635 89.405 116.685 ;
        RECT 87.270 116.185 88.145 116.515 ;
        RECT 88.315 116.185 89.065 116.515 ;
        RECT 87.270 115.725 87.440 116.185 ;
        RECT 88.315 116.015 88.515 116.185 ;
        RECT 89.235 116.055 89.405 116.635 ;
        RECT 89.180 116.015 89.405 116.055 ;
        RECT 86.080 115.555 86.485 115.725 ;
        RECT 86.655 115.555 87.440 115.725 ;
        RECT 87.715 115.275 87.925 115.805 ;
        RECT 88.185 115.490 88.515 116.015 ;
        RECT 89.025 115.930 89.405 116.015 ;
        RECT 90.500 116.685 90.835 117.655 ;
        RECT 91.005 116.685 91.175 117.825 ;
        RECT 91.345 117.485 93.375 117.655 ;
        RECT 90.500 116.015 90.670 116.685 ;
        RECT 91.345 116.515 91.515 117.485 ;
        RECT 90.840 116.185 91.095 116.515 ;
        RECT 91.320 116.185 91.515 116.515 ;
        RECT 91.685 117.145 92.810 117.315 ;
        RECT 90.925 116.015 91.095 116.185 ;
        RECT 91.685 116.015 91.855 117.145 ;
        RECT 88.685 115.275 88.855 115.885 ;
        RECT 89.025 115.495 89.355 115.930 ;
        RECT 90.500 115.445 90.755 116.015 ;
        RECT 90.925 115.845 91.855 116.015 ;
        RECT 92.025 116.805 93.035 116.975 ;
        RECT 92.025 116.005 92.195 116.805 ;
        RECT 91.680 115.810 91.855 115.845 ;
        RECT 90.925 115.275 91.255 115.675 ;
        RECT 91.680 115.445 92.210 115.810 ;
        RECT 92.400 115.785 92.675 116.605 ;
        RECT 92.395 115.615 92.675 115.785 ;
        RECT 92.400 115.445 92.675 115.615 ;
        RECT 92.845 115.445 93.035 116.805 ;
        RECT 93.205 116.820 93.375 117.485 ;
        RECT 93.545 117.065 93.715 117.825 ;
        RECT 93.950 117.065 94.465 117.475 ;
        RECT 93.205 116.630 93.955 116.820 ;
        RECT 94.125 116.255 94.465 117.065 ;
        RECT 94.640 116.685 94.895 117.825 ;
        RECT 95.065 116.855 95.395 117.655 ;
        RECT 95.565 117.025 95.735 117.825 ;
        RECT 95.905 116.855 96.235 117.655 ;
        RECT 96.405 117.025 96.575 117.825 ;
        RECT 96.745 116.855 97.075 117.655 ;
        RECT 97.245 117.025 97.415 117.825 ;
        RECT 97.585 116.855 97.915 117.655 ;
        RECT 98.085 117.025 98.335 117.825 ;
        RECT 99.045 117.025 99.295 117.825 ;
        RECT 95.065 116.685 97.915 116.855 ;
        RECT 99.465 116.855 99.795 117.655 ;
        RECT 99.965 117.025 100.135 117.825 ;
        RECT 100.305 116.855 100.635 117.655 ;
        RECT 100.805 117.025 100.975 117.825 ;
        RECT 101.145 116.855 101.475 117.655 ;
        RECT 101.645 117.025 101.815 117.825 ;
        RECT 101.985 116.855 102.315 117.655 ;
        RECT 99.465 116.685 102.315 116.855 ;
        RECT 102.485 116.685 102.740 117.825 ;
        RECT 103.380 116.685 103.715 117.655 ;
        RECT 103.885 116.685 104.055 117.825 ;
        RECT 104.225 117.485 106.255 117.655 ;
        RECT 94.660 116.265 96.280 116.515 ;
        RECT 96.460 116.265 96.995 116.685 ;
        RECT 97.165 116.265 98.605 116.515 ;
        RECT 98.775 116.265 100.215 116.515 ;
        RECT 100.385 116.265 100.920 116.685 ;
        RECT 101.100 116.265 102.720 116.515 ;
        RECT 93.235 116.085 94.465 116.255 ;
        RECT 93.215 115.275 93.725 115.810 ;
        RECT 93.945 115.480 94.190 116.085 ;
        RECT 94.640 115.905 96.575 116.095 ;
        RECT 94.640 115.445 94.975 115.905 ;
        RECT 95.145 115.275 95.315 115.735 ;
        RECT 95.485 115.445 95.815 115.905 ;
        RECT 95.985 115.275 96.155 115.735 ;
        RECT 96.325 115.655 96.575 115.905 ;
        RECT 96.745 115.995 96.995 116.265 ;
        RECT 96.745 115.825 97.915 115.995 ;
        RECT 98.085 115.655 98.335 116.075 ;
        RECT 96.325 115.445 98.335 115.655 ;
        RECT 99.045 115.655 99.295 116.075 ;
        RECT 100.385 115.995 100.635 116.265 ;
        RECT 99.465 115.825 100.635 115.995 ;
        RECT 100.805 115.905 102.740 116.095 ;
        RECT 100.805 115.655 101.055 115.905 ;
        RECT 99.045 115.445 101.055 115.655 ;
        RECT 101.225 115.275 101.395 115.735 ;
        RECT 101.565 115.445 101.895 115.905 ;
        RECT 102.065 115.275 102.235 115.735 ;
        RECT 102.405 115.445 102.740 115.905 ;
        RECT 103.380 116.015 103.550 116.685 ;
        RECT 104.225 116.515 104.395 117.485 ;
        RECT 103.720 116.185 103.975 116.515 ;
        RECT 104.200 116.185 104.395 116.515 ;
        RECT 104.565 117.145 105.690 117.315 ;
        RECT 103.805 116.015 103.975 116.185 ;
        RECT 104.565 116.015 104.735 117.145 ;
        RECT 103.380 115.445 103.635 116.015 ;
        RECT 103.805 115.845 104.735 116.015 ;
        RECT 104.905 116.805 105.915 116.975 ;
        RECT 104.905 116.005 105.075 116.805 ;
        RECT 105.280 116.465 105.555 116.605 ;
        RECT 105.275 116.295 105.555 116.465 ;
        RECT 104.560 115.810 104.735 115.845 ;
        RECT 103.805 115.275 104.135 115.675 ;
        RECT 104.560 115.445 105.090 115.810 ;
        RECT 105.280 115.445 105.555 116.295 ;
        RECT 105.725 115.445 105.915 116.805 ;
        RECT 106.085 116.820 106.255 117.485 ;
        RECT 106.425 117.065 106.595 117.825 ;
        RECT 106.830 117.065 107.345 117.475 ;
        RECT 106.085 116.630 106.835 116.820 ;
        RECT 107.005 116.255 107.345 117.065 ;
        RECT 107.515 116.660 107.805 117.825 ;
        RECT 108.035 116.765 108.365 117.610 ;
        RECT 108.535 116.815 108.705 117.825 ;
        RECT 108.875 117.095 109.215 117.655 ;
        RECT 109.445 117.325 109.760 117.825 ;
        RECT 109.940 117.355 110.825 117.525 ;
        RECT 107.975 116.685 108.365 116.765 ;
        RECT 108.875 116.720 109.770 117.095 ;
        RECT 106.115 116.085 107.345 116.255 ;
        RECT 107.975 116.635 108.190 116.685 ;
        RECT 106.095 115.275 106.605 115.810 ;
        RECT 106.825 115.480 107.070 116.085 ;
        RECT 107.975 116.055 108.145 116.635 ;
        RECT 108.875 116.515 109.065 116.720 ;
        RECT 109.940 116.515 110.110 117.355 ;
        RECT 111.050 117.325 111.300 117.655 ;
        RECT 108.315 116.185 109.065 116.515 ;
        RECT 109.235 116.185 110.110 116.515 ;
        RECT 107.975 116.015 108.200 116.055 ;
        RECT 108.865 116.015 109.065 116.185 ;
        RECT 107.515 115.275 107.805 116.000 ;
        RECT 107.975 115.930 108.355 116.015 ;
        RECT 108.025 115.495 108.355 115.930 ;
        RECT 108.525 115.275 108.695 115.885 ;
        RECT 108.865 115.490 109.195 116.015 ;
        RECT 109.455 115.275 109.665 115.805 ;
        RECT 109.940 115.725 110.110 116.185 ;
        RECT 110.280 116.225 110.600 117.185 ;
        RECT 110.770 116.435 110.960 117.155 ;
        RECT 111.130 116.255 111.300 117.325 ;
        RECT 111.470 117.025 111.640 117.825 ;
        RECT 111.810 117.380 112.915 117.550 ;
        RECT 111.810 116.765 111.980 117.380 ;
        RECT 113.125 117.230 113.375 117.655 ;
        RECT 113.545 117.365 113.810 117.825 ;
        RECT 112.150 116.845 112.680 117.210 ;
        RECT 113.125 117.100 113.430 117.230 ;
        RECT 111.470 116.675 111.980 116.765 ;
        RECT 111.470 116.505 112.340 116.675 ;
        RECT 111.470 116.435 111.640 116.505 ;
        RECT 111.760 116.255 111.960 116.285 ;
        RECT 110.280 115.895 110.745 116.225 ;
        RECT 111.130 115.955 111.960 116.255 ;
        RECT 111.130 115.725 111.300 115.955 ;
        RECT 109.940 115.555 110.725 115.725 ;
        RECT 110.895 115.555 111.300 115.725 ;
        RECT 111.480 115.275 111.850 115.775 ;
        RECT 112.170 115.725 112.340 116.505 ;
        RECT 112.510 116.145 112.680 116.845 ;
        RECT 112.850 116.315 113.090 116.910 ;
        RECT 112.510 115.925 113.035 116.145 ;
        RECT 113.260 115.995 113.430 117.100 ;
        RECT 113.205 115.865 113.430 115.995 ;
        RECT 113.600 115.905 113.880 116.855 ;
        RECT 113.205 115.725 113.375 115.865 ;
        RECT 112.170 115.555 112.845 115.725 ;
        RECT 113.040 115.555 113.375 115.725 ;
        RECT 113.545 115.275 113.795 115.735 ;
        RECT 114.050 115.535 114.235 117.655 ;
        RECT 114.405 117.325 114.735 117.825 ;
        RECT 114.905 117.155 115.075 117.655 ;
        RECT 115.335 117.390 120.680 117.825 ;
        RECT 114.410 116.985 115.075 117.155 ;
        RECT 114.410 115.995 114.640 116.985 ;
        RECT 114.810 116.165 115.160 116.815 ;
        RECT 114.410 115.825 115.075 115.995 ;
        RECT 114.405 115.275 114.735 115.655 ;
        RECT 114.905 115.535 115.075 115.825 ;
        RECT 116.920 115.820 117.260 116.650 ;
        RECT 118.740 116.140 119.090 117.390 ;
        RECT 121.405 117.205 121.575 117.635 ;
        RECT 121.745 117.375 122.075 117.825 ;
        RECT 121.405 116.975 122.080 117.205 ;
        RECT 121.375 115.955 121.675 116.805 ;
        RECT 121.845 116.325 122.080 116.975 ;
        RECT 122.250 116.665 122.535 117.610 ;
        RECT 122.715 117.355 123.400 117.825 ;
        RECT 122.710 116.835 123.405 117.145 ;
        RECT 123.580 116.770 123.885 117.555 ;
        RECT 122.250 116.515 123.110 116.665 ;
        RECT 122.250 116.495 123.535 116.515 ;
        RECT 121.845 115.995 122.380 116.325 ;
        RECT 122.550 116.135 123.535 116.495 ;
        RECT 121.845 115.845 122.065 115.995 ;
        RECT 115.335 115.275 120.680 115.820 ;
        RECT 121.320 115.275 121.655 115.780 ;
        RECT 121.825 115.470 122.065 115.845 ;
        RECT 122.550 115.800 122.720 116.135 ;
        RECT 123.710 115.965 123.885 116.770 ;
        RECT 122.345 115.605 122.720 115.800 ;
        RECT 122.345 115.460 122.515 115.605 ;
        RECT 123.080 115.275 123.475 115.770 ;
        RECT 123.645 115.445 123.885 115.965 ;
        RECT 124.095 116.770 124.400 117.555 ;
        RECT 124.580 117.355 125.265 117.825 ;
        RECT 124.575 116.835 125.270 117.145 ;
        RECT 124.095 115.965 124.270 116.770 ;
        RECT 125.445 116.665 125.730 117.610 ;
        RECT 125.905 117.375 126.235 117.825 ;
        RECT 126.405 117.205 126.575 117.635 ;
        RECT 126.835 117.390 132.180 117.825 ;
        RECT 124.870 116.515 125.730 116.665 ;
        RECT 124.445 116.495 125.730 116.515 ;
        RECT 125.900 116.975 126.575 117.205 ;
        RECT 124.445 116.135 125.430 116.495 ;
        RECT 125.900 116.325 126.135 116.975 ;
        RECT 124.095 115.445 124.335 115.965 ;
        RECT 125.260 115.800 125.430 116.135 ;
        RECT 125.600 115.995 126.135 116.325 ;
        RECT 125.915 115.845 126.135 115.995 ;
        RECT 126.305 115.955 126.605 116.805 ;
        RECT 124.505 115.275 124.900 115.770 ;
        RECT 125.260 115.605 125.635 115.800 ;
        RECT 125.465 115.460 125.635 115.605 ;
        RECT 125.915 115.470 126.155 115.845 ;
        RECT 128.420 115.820 128.760 116.650 ;
        RECT 130.240 116.140 130.590 117.390 ;
        RECT 133.275 116.660 133.565 117.825 ;
        RECT 133.735 116.735 136.325 117.825 ;
        RECT 133.735 116.045 134.945 116.565 ;
        RECT 135.115 116.215 136.325 116.735 ;
        RECT 136.500 116.685 136.835 117.655 ;
        RECT 137.005 116.685 137.175 117.825 ;
        RECT 137.345 117.485 139.375 117.655 ;
        RECT 126.325 115.275 126.660 115.780 ;
        RECT 126.835 115.275 132.180 115.820 ;
        RECT 133.275 115.275 133.565 116.000 ;
        RECT 133.735 115.275 136.325 116.045 ;
        RECT 136.500 116.015 136.670 116.685 ;
        RECT 137.345 116.515 137.515 117.485 ;
        RECT 136.840 116.185 137.095 116.515 ;
        RECT 137.320 116.185 137.515 116.515 ;
        RECT 137.685 117.145 138.810 117.315 ;
        RECT 136.925 116.015 137.095 116.185 ;
        RECT 137.685 116.015 137.855 117.145 ;
        RECT 136.500 115.445 136.755 116.015 ;
        RECT 136.925 115.845 137.855 116.015 ;
        RECT 138.025 116.805 139.035 116.975 ;
        RECT 138.025 116.005 138.195 116.805 ;
        RECT 138.400 116.465 138.675 116.605 ;
        RECT 138.395 116.295 138.675 116.465 ;
        RECT 137.680 115.810 137.855 115.845 ;
        RECT 136.925 115.275 137.255 115.675 ;
        RECT 137.680 115.445 138.210 115.810 ;
        RECT 138.400 115.445 138.675 116.295 ;
        RECT 138.845 115.445 139.035 116.805 ;
        RECT 139.205 116.820 139.375 117.485 ;
        RECT 139.545 117.065 139.715 117.825 ;
        RECT 139.950 117.065 140.465 117.475 ;
        RECT 139.205 116.630 139.955 116.820 ;
        RECT 140.125 116.255 140.465 117.065 ;
        RECT 139.235 116.085 140.465 116.255 ;
        RECT 140.655 116.985 140.910 117.655 ;
        RECT 141.080 117.065 141.410 117.825 ;
        RECT 141.580 117.225 141.830 117.655 ;
        RECT 142.000 117.405 142.355 117.825 ;
        RECT 142.545 117.485 143.715 117.655 ;
        RECT 142.545 117.445 142.875 117.485 ;
        RECT 142.985 117.225 143.215 117.315 ;
        RECT 141.580 116.985 143.215 117.225 ;
        RECT 143.385 116.985 143.715 117.485 ;
        RECT 139.215 115.275 139.725 115.810 ;
        RECT 139.945 115.480 140.190 116.085 ;
        RECT 140.655 115.855 140.825 116.985 ;
        RECT 143.885 116.815 144.055 117.655 ;
        RECT 140.995 116.645 144.055 116.815 ;
        RECT 144.315 116.735 145.525 117.825 ;
        RECT 140.995 116.095 141.165 116.645 ;
        RECT 141.395 116.265 141.760 116.465 ;
        RECT 141.930 116.265 142.260 116.465 ;
        RECT 140.995 115.925 141.795 116.095 ;
        RECT 140.655 115.785 140.840 115.855 ;
        RECT 140.655 115.775 140.865 115.785 ;
        RECT 140.655 115.445 140.910 115.775 ;
        RECT 141.125 115.275 141.455 115.755 ;
        RECT 141.625 115.695 141.795 115.925 ;
        RECT 141.975 115.865 142.260 116.265 ;
        RECT 142.530 116.265 143.005 116.465 ;
        RECT 143.175 116.265 143.620 116.465 ;
        RECT 143.790 116.265 144.140 116.475 ;
        RECT 142.530 115.865 142.810 116.265 ;
        RECT 142.990 115.925 144.055 116.095 ;
        RECT 142.990 115.695 143.160 115.925 ;
        RECT 141.625 115.445 143.160 115.695 ;
        RECT 143.385 115.275 143.715 115.755 ;
        RECT 143.885 115.445 144.055 115.925 ;
        RECT 144.315 116.025 144.835 116.565 ;
        RECT 145.005 116.195 145.525 116.735 ;
        RECT 145.695 116.735 146.905 117.825 ;
        RECT 145.695 116.195 146.215 116.735 ;
        RECT 146.385 116.025 146.905 116.565 ;
        RECT 144.315 115.275 145.525 116.025 ;
        RECT 145.695 115.275 146.905 116.025 ;
        RECT 17.270 115.105 146.990 115.275 ;
        RECT 17.355 114.355 18.565 115.105 ;
        RECT 17.355 113.815 17.875 114.355 ;
        RECT 18.740 114.265 19.000 115.105 ;
        RECT 19.175 114.360 19.430 114.935 ;
        RECT 19.600 114.725 19.930 115.105 ;
        RECT 20.145 114.555 20.315 114.935 ;
        RECT 19.600 114.385 20.315 114.555 ;
        RECT 18.045 113.645 18.565 114.185 ;
        RECT 17.355 112.555 18.565 113.645 ;
        RECT 18.740 112.555 19.000 113.705 ;
        RECT 19.175 113.630 19.345 114.360 ;
        RECT 19.600 114.195 19.770 114.385 ;
        RECT 20.575 114.335 22.245 115.105 ;
        RECT 19.515 113.865 19.770 114.195 ;
        RECT 19.600 113.655 19.770 113.865 ;
        RECT 20.050 113.835 20.405 114.205 ;
        RECT 20.575 113.815 21.325 114.335 ;
        RECT 22.690 114.295 22.935 114.900 ;
        RECT 23.155 114.570 23.665 115.105 ;
        RECT 19.175 112.725 19.430 113.630 ;
        RECT 19.600 113.485 20.315 113.655 ;
        RECT 21.495 113.645 22.245 114.165 ;
        RECT 19.600 112.555 19.930 113.315 ;
        RECT 20.145 112.725 20.315 113.485 ;
        RECT 20.575 112.555 22.245 113.645 ;
        RECT 22.415 114.125 23.645 114.295 ;
        RECT 22.415 113.315 22.755 114.125 ;
        RECT 22.925 113.560 23.675 113.750 ;
        RECT 22.415 112.905 22.930 113.315 ;
        RECT 23.165 112.555 23.335 113.315 ;
        RECT 23.505 112.895 23.675 113.560 ;
        RECT 23.845 113.575 24.035 114.935 ;
        RECT 24.205 114.085 24.480 114.935 ;
        RECT 24.670 114.570 25.200 114.935 ;
        RECT 25.625 114.705 25.955 115.105 ;
        RECT 25.025 114.535 25.200 114.570 ;
        RECT 24.205 113.915 24.485 114.085 ;
        RECT 24.205 113.775 24.480 113.915 ;
        RECT 24.685 113.575 24.855 114.375 ;
        RECT 23.845 113.405 24.855 113.575 ;
        RECT 25.025 114.365 25.955 114.535 ;
        RECT 26.125 114.365 26.380 114.935 ;
        RECT 27.105 114.555 27.275 114.845 ;
        RECT 27.445 114.725 27.775 115.105 ;
        RECT 27.105 114.385 27.770 114.555 ;
        RECT 25.025 113.235 25.195 114.365 ;
        RECT 25.785 114.195 25.955 114.365 ;
        RECT 24.070 113.065 25.195 113.235 ;
        RECT 25.365 113.865 25.560 114.195 ;
        RECT 25.785 113.865 26.040 114.195 ;
        RECT 25.365 112.895 25.535 113.865 ;
        RECT 26.210 113.695 26.380 114.365 ;
        RECT 23.505 112.725 25.535 112.895 ;
        RECT 25.705 112.555 25.875 113.695 ;
        RECT 26.045 112.725 26.380 113.695 ;
        RECT 27.020 113.565 27.370 114.215 ;
        RECT 27.540 113.395 27.770 114.385 ;
        RECT 27.105 113.225 27.770 113.395 ;
        RECT 27.105 112.725 27.275 113.225 ;
        RECT 27.445 112.555 27.775 113.055 ;
        RECT 27.945 112.725 28.130 114.845 ;
        RECT 28.385 114.645 28.635 115.105 ;
        RECT 28.805 114.655 29.140 114.825 ;
        RECT 29.335 114.655 30.010 114.825 ;
        RECT 28.805 114.515 28.975 114.655 ;
        RECT 28.300 113.525 28.580 114.475 ;
        RECT 28.750 114.385 28.975 114.515 ;
        RECT 28.750 113.280 28.920 114.385 ;
        RECT 29.145 114.235 29.670 114.455 ;
        RECT 29.090 113.470 29.330 114.065 ;
        RECT 29.500 113.535 29.670 114.235 ;
        RECT 29.840 113.875 30.010 114.655 ;
        RECT 30.330 114.605 30.700 115.105 ;
        RECT 30.880 114.655 31.285 114.825 ;
        RECT 31.455 114.655 32.240 114.825 ;
        RECT 30.880 114.425 31.050 114.655 ;
        RECT 30.220 114.125 31.050 114.425 ;
        RECT 31.435 114.155 31.900 114.485 ;
        RECT 30.220 114.095 30.420 114.125 ;
        RECT 30.540 113.875 30.710 113.945 ;
        RECT 29.840 113.705 30.710 113.875 ;
        RECT 30.200 113.615 30.710 113.705 ;
        RECT 28.750 113.150 29.055 113.280 ;
        RECT 29.500 113.170 30.030 113.535 ;
        RECT 28.370 112.555 28.635 113.015 ;
        RECT 28.805 112.725 29.055 113.150 ;
        RECT 30.200 113.000 30.370 113.615 ;
        RECT 29.265 112.830 30.370 113.000 ;
        RECT 30.540 112.555 30.710 113.355 ;
        RECT 30.880 113.055 31.050 114.125 ;
        RECT 31.220 113.225 31.410 113.945 ;
        RECT 31.580 113.195 31.900 114.155 ;
        RECT 32.070 114.195 32.240 114.655 ;
        RECT 32.515 114.575 32.725 115.105 ;
        RECT 32.985 114.365 33.315 114.890 ;
        RECT 33.485 114.495 33.655 115.105 ;
        RECT 33.825 114.450 34.155 114.885 ;
        RECT 34.375 114.560 39.720 115.105 ;
        RECT 33.825 114.365 34.205 114.450 ;
        RECT 33.115 114.195 33.315 114.365 ;
        RECT 33.980 114.325 34.205 114.365 ;
        RECT 32.070 113.865 32.945 114.195 ;
        RECT 33.115 113.865 33.865 114.195 ;
        RECT 30.880 112.725 31.130 113.055 ;
        RECT 32.070 113.025 32.240 113.865 ;
        RECT 33.115 113.660 33.305 113.865 ;
        RECT 34.035 113.745 34.205 114.325 ;
        RECT 33.990 113.695 34.205 113.745 ;
        RECT 35.960 113.730 36.300 114.560 ;
        RECT 39.895 114.335 42.485 115.105 ;
        RECT 43.115 114.380 43.405 115.105 ;
        RECT 43.575 114.560 48.920 115.105 ;
        RECT 49.095 114.560 54.440 115.105 ;
        RECT 54.615 114.560 59.960 115.105 ;
        RECT 60.135 114.560 65.480 115.105 ;
        RECT 32.410 113.285 33.305 113.660 ;
        RECT 33.815 113.615 34.205 113.695 ;
        RECT 31.355 112.855 32.240 113.025 ;
        RECT 32.420 112.555 32.735 113.055 ;
        RECT 32.965 112.725 33.305 113.285 ;
        RECT 33.475 112.555 33.645 113.565 ;
        RECT 33.815 112.770 34.145 113.615 ;
        RECT 37.780 112.990 38.130 114.240 ;
        RECT 39.895 113.815 41.105 114.335 ;
        RECT 41.275 113.645 42.485 114.165 ;
        RECT 45.160 113.730 45.500 114.560 ;
        RECT 34.375 112.555 39.720 112.990 ;
        RECT 39.895 112.555 42.485 113.645 ;
        RECT 43.115 112.555 43.405 113.720 ;
        RECT 46.980 112.990 47.330 114.240 ;
        RECT 50.680 113.730 51.020 114.560 ;
        RECT 52.500 112.990 52.850 114.240 ;
        RECT 56.200 113.730 56.540 114.560 ;
        RECT 58.020 112.990 58.370 114.240 ;
        RECT 61.720 113.730 62.060 114.560 ;
        RECT 65.655 114.335 68.245 115.105 ;
        RECT 68.875 114.380 69.165 115.105 ;
        RECT 69.335 114.335 71.005 115.105 ;
        RECT 71.265 114.555 71.435 114.845 ;
        RECT 71.605 114.725 71.935 115.105 ;
        RECT 71.265 114.385 71.930 114.555 ;
        RECT 63.540 112.990 63.890 114.240 ;
        RECT 65.655 113.815 66.865 114.335 ;
        RECT 67.035 113.645 68.245 114.165 ;
        RECT 69.335 113.815 70.085 114.335 ;
        RECT 43.575 112.555 48.920 112.990 ;
        RECT 49.095 112.555 54.440 112.990 ;
        RECT 54.615 112.555 59.960 112.990 ;
        RECT 60.135 112.555 65.480 112.990 ;
        RECT 65.655 112.555 68.245 113.645 ;
        RECT 68.875 112.555 69.165 113.720 ;
        RECT 70.255 113.645 71.005 114.165 ;
        RECT 69.335 112.555 71.005 113.645 ;
        RECT 71.180 113.565 71.530 114.215 ;
        RECT 71.700 113.395 71.930 114.385 ;
        RECT 71.265 113.225 71.930 113.395 ;
        RECT 71.265 112.725 71.435 113.225 ;
        RECT 71.605 112.555 71.935 113.055 ;
        RECT 72.105 112.725 72.290 114.845 ;
        RECT 72.545 114.645 72.795 115.105 ;
        RECT 72.965 114.655 73.300 114.825 ;
        RECT 73.495 114.655 74.170 114.825 ;
        RECT 72.965 114.515 73.135 114.655 ;
        RECT 72.460 113.525 72.740 114.475 ;
        RECT 72.910 114.385 73.135 114.515 ;
        RECT 72.910 113.280 73.080 114.385 ;
        RECT 73.305 114.235 73.830 114.455 ;
        RECT 73.250 113.470 73.490 114.065 ;
        RECT 73.660 113.535 73.830 114.235 ;
        RECT 74.000 113.875 74.170 114.655 ;
        RECT 74.490 114.605 74.860 115.105 ;
        RECT 75.040 114.655 75.445 114.825 ;
        RECT 75.615 114.655 76.400 114.825 ;
        RECT 75.040 114.425 75.210 114.655 ;
        RECT 74.380 114.125 75.210 114.425 ;
        RECT 75.595 114.155 76.060 114.485 ;
        RECT 74.380 114.095 74.580 114.125 ;
        RECT 74.700 113.875 74.870 113.945 ;
        RECT 74.000 113.705 74.870 113.875 ;
        RECT 74.360 113.615 74.870 113.705 ;
        RECT 72.910 113.150 73.215 113.280 ;
        RECT 73.660 113.170 74.190 113.535 ;
        RECT 72.530 112.555 72.795 113.015 ;
        RECT 72.965 112.725 73.215 113.150 ;
        RECT 74.360 113.000 74.530 113.615 ;
        RECT 73.425 112.830 74.530 113.000 ;
        RECT 74.700 112.555 74.870 113.355 ;
        RECT 75.040 113.055 75.210 114.125 ;
        RECT 75.380 113.225 75.570 113.945 ;
        RECT 75.740 113.195 76.060 114.155 ;
        RECT 76.230 114.195 76.400 114.655 ;
        RECT 76.675 114.575 76.885 115.105 ;
        RECT 77.145 114.365 77.475 114.890 ;
        RECT 77.645 114.495 77.815 115.105 ;
        RECT 77.985 114.450 78.315 114.885 ;
        RECT 77.985 114.365 78.365 114.450 ;
        RECT 77.275 114.195 77.475 114.365 ;
        RECT 78.140 114.325 78.365 114.365 ;
        RECT 76.230 113.865 77.105 114.195 ;
        RECT 77.275 113.865 78.025 114.195 ;
        RECT 75.040 112.725 75.290 113.055 ;
        RECT 76.230 113.025 76.400 113.865 ;
        RECT 77.275 113.660 77.465 113.865 ;
        RECT 78.195 113.745 78.365 114.325 ;
        RECT 78.150 113.695 78.365 113.745 ;
        RECT 76.570 113.285 77.465 113.660 ;
        RECT 77.975 113.615 78.365 113.695 ;
        RECT 78.540 114.365 78.795 114.935 ;
        RECT 78.965 114.705 79.295 115.105 ;
        RECT 79.720 114.570 80.250 114.935 ;
        RECT 79.720 114.535 79.895 114.570 ;
        RECT 78.965 114.365 79.895 114.535 ;
        RECT 80.440 114.425 80.715 114.935 ;
        RECT 78.540 113.695 78.710 114.365 ;
        RECT 78.965 114.195 79.135 114.365 ;
        RECT 78.880 113.865 79.135 114.195 ;
        RECT 79.360 113.865 79.555 114.195 ;
        RECT 75.515 112.855 76.400 113.025 ;
        RECT 76.580 112.555 76.895 113.055 ;
        RECT 77.125 112.725 77.465 113.285 ;
        RECT 77.635 112.555 77.805 113.565 ;
        RECT 77.975 112.770 78.305 113.615 ;
        RECT 78.540 112.725 78.875 113.695 ;
        RECT 79.045 112.555 79.215 113.695 ;
        RECT 79.385 112.895 79.555 113.865 ;
        RECT 79.725 113.235 79.895 114.365 ;
        RECT 80.065 113.575 80.235 114.375 ;
        RECT 80.435 114.255 80.715 114.425 ;
        RECT 80.440 113.775 80.715 114.255 ;
        RECT 80.885 113.575 81.075 114.935 ;
        RECT 81.255 114.570 81.765 115.105 ;
        RECT 81.985 114.295 82.230 114.900 ;
        RECT 82.765 114.455 82.935 114.935 ;
        RECT 83.105 114.625 83.435 115.105 ;
        RECT 83.660 114.685 85.195 114.935 ;
        RECT 83.660 114.455 83.830 114.685 ;
        RECT 81.275 114.125 82.505 114.295 ;
        RECT 82.765 114.285 83.830 114.455 ;
        RECT 80.065 113.405 81.075 113.575 ;
        RECT 81.245 113.560 81.995 113.750 ;
        RECT 79.725 113.065 80.850 113.235 ;
        RECT 81.245 112.895 81.415 113.560 ;
        RECT 82.165 113.315 82.505 114.125 ;
        RECT 84.010 114.115 84.290 114.515 ;
        RECT 82.680 113.905 83.030 114.115 ;
        RECT 83.200 113.915 83.645 114.115 ;
        RECT 83.815 113.915 84.290 114.115 ;
        RECT 84.560 114.115 84.845 114.515 ;
        RECT 85.025 114.455 85.195 114.685 ;
        RECT 85.365 114.625 85.695 115.105 ;
        RECT 85.910 114.605 86.165 114.935 ;
        RECT 85.955 114.595 86.165 114.605 ;
        RECT 85.980 114.525 86.165 114.595 ;
        RECT 85.025 114.285 85.825 114.455 ;
        RECT 84.560 113.915 84.890 114.115 ;
        RECT 85.060 113.915 85.425 114.115 ;
        RECT 85.655 113.735 85.825 114.285 ;
        RECT 79.385 112.725 81.415 112.895 ;
        RECT 81.585 112.555 81.755 113.315 ;
        RECT 81.990 112.905 82.505 113.315 ;
        RECT 82.765 113.565 85.825 113.735 ;
        RECT 82.765 112.725 82.935 113.565 ;
        RECT 85.995 113.395 86.165 114.525 ;
        RECT 86.905 114.555 87.075 114.845 ;
        RECT 87.245 114.725 87.575 115.105 ;
        RECT 86.905 114.385 87.570 114.555 ;
        RECT 86.820 113.565 87.170 114.215 ;
        RECT 87.340 113.395 87.570 114.385 ;
        RECT 83.105 112.895 83.435 113.395 ;
        RECT 83.605 113.155 85.240 113.395 ;
        RECT 83.605 113.065 83.835 113.155 ;
        RECT 83.945 112.895 84.275 112.935 ;
        RECT 83.105 112.725 84.275 112.895 ;
        RECT 84.465 112.555 84.820 112.975 ;
        RECT 84.990 112.725 85.240 113.155 ;
        RECT 85.410 112.555 85.740 113.315 ;
        RECT 85.910 112.725 86.165 113.395 ;
        RECT 86.905 113.225 87.570 113.395 ;
        RECT 86.905 112.725 87.075 113.225 ;
        RECT 87.245 112.555 87.575 113.055 ;
        RECT 87.745 112.725 87.930 114.845 ;
        RECT 88.185 114.645 88.435 115.105 ;
        RECT 88.605 114.655 88.940 114.825 ;
        RECT 89.135 114.655 89.810 114.825 ;
        RECT 88.605 114.515 88.775 114.655 ;
        RECT 88.100 113.525 88.380 114.475 ;
        RECT 88.550 114.385 88.775 114.515 ;
        RECT 88.550 113.280 88.720 114.385 ;
        RECT 88.945 114.235 89.470 114.455 ;
        RECT 88.890 113.470 89.130 114.065 ;
        RECT 89.300 113.535 89.470 114.235 ;
        RECT 89.640 113.875 89.810 114.655 ;
        RECT 90.130 114.605 90.500 115.105 ;
        RECT 90.680 114.655 91.085 114.825 ;
        RECT 91.255 114.655 92.040 114.825 ;
        RECT 90.680 114.425 90.850 114.655 ;
        RECT 90.020 114.125 90.850 114.425 ;
        RECT 91.235 114.155 91.700 114.485 ;
        RECT 90.020 114.095 90.220 114.125 ;
        RECT 90.340 113.875 90.510 113.945 ;
        RECT 89.640 113.705 90.510 113.875 ;
        RECT 90.000 113.615 90.510 113.705 ;
        RECT 88.550 113.150 88.855 113.280 ;
        RECT 89.300 113.170 89.830 113.535 ;
        RECT 88.170 112.555 88.435 113.015 ;
        RECT 88.605 112.725 88.855 113.150 ;
        RECT 90.000 113.000 90.170 113.615 ;
        RECT 89.065 112.830 90.170 113.000 ;
        RECT 90.340 112.555 90.510 113.355 ;
        RECT 90.680 113.055 90.850 114.125 ;
        RECT 91.020 113.225 91.210 113.945 ;
        RECT 91.380 113.195 91.700 114.155 ;
        RECT 91.870 114.195 92.040 114.655 ;
        RECT 92.315 114.575 92.525 115.105 ;
        RECT 92.785 114.365 93.115 114.890 ;
        RECT 93.285 114.495 93.455 115.105 ;
        RECT 93.625 114.450 93.955 114.885 ;
        RECT 93.625 114.365 94.005 114.450 ;
        RECT 94.635 114.380 94.925 115.105 ;
        RECT 95.365 114.725 97.375 114.935 ;
        RECT 92.915 114.195 93.115 114.365 ;
        RECT 93.780 114.325 94.005 114.365 ;
        RECT 91.870 113.865 92.745 114.195 ;
        RECT 92.915 113.865 93.665 114.195 ;
        RECT 90.680 112.725 90.930 113.055 ;
        RECT 91.870 113.025 92.040 113.865 ;
        RECT 92.915 113.660 93.105 113.865 ;
        RECT 93.835 113.745 94.005 114.325 ;
        RECT 95.365 114.305 95.615 114.725 ;
        RECT 95.785 114.385 96.955 114.555 ;
        RECT 96.705 114.115 96.955 114.385 ;
        RECT 97.125 114.475 97.375 114.725 ;
        RECT 97.545 114.645 97.715 115.105 ;
        RECT 97.885 114.475 98.215 114.935 ;
        RECT 98.385 114.645 98.555 115.105 ;
        RECT 98.725 114.475 99.060 114.935 ;
        RECT 97.125 114.285 99.060 114.475 ;
        RECT 99.235 114.355 100.445 115.105 ;
        RECT 100.620 114.705 100.955 115.105 ;
        RECT 101.125 114.535 101.330 114.935 ;
        RECT 101.540 114.625 101.815 115.105 ;
        RECT 102.025 114.605 102.285 114.935 ;
        RECT 100.645 114.365 101.330 114.535 ;
        RECT 95.095 113.865 96.535 114.115 ;
        RECT 93.790 113.695 94.005 113.745 ;
        RECT 92.210 113.285 93.105 113.660 ;
        RECT 93.615 113.615 94.005 113.695 ;
        RECT 91.155 112.855 92.040 113.025 ;
        RECT 92.220 112.555 92.535 113.055 ;
        RECT 92.765 112.725 93.105 113.285 ;
        RECT 93.275 112.555 93.445 113.565 ;
        RECT 93.615 112.770 93.945 113.615 ;
        RECT 94.635 112.555 94.925 113.720 ;
        RECT 96.705 113.695 97.240 114.115 ;
        RECT 97.420 113.865 99.040 114.115 ;
        RECT 99.235 113.815 99.755 114.355 ;
        RECT 95.785 113.525 98.635 113.695 ;
        RECT 95.365 112.555 95.615 113.355 ;
        RECT 95.785 112.725 96.115 113.525 ;
        RECT 96.285 112.555 96.455 113.355 ;
        RECT 96.625 112.725 96.955 113.525 ;
        RECT 97.125 112.555 97.295 113.355 ;
        RECT 97.465 112.725 97.795 113.525 ;
        RECT 97.965 112.555 98.135 113.355 ;
        RECT 98.305 112.725 98.635 113.525 ;
        RECT 98.805 112.555 99.060 113.695 ;
        RECT 99.925 113.645 100.445 114.185 ;
        RECT 99.235 112.555 100.445 113.645 ;
        RECT 100.645 113.335 100.985 114.365 ;
        RECT 101.155 113.695 101.405 114.195 ;
        RECT 101.585 113.865 101.945 114.445 ;
        RECT 102.115 113.695 102.285 114.605 ;
        RECT 102.545 114.555 102.715 114.845 ;
        RECT 102.885 114.725 103.215 115.105 ;
        RECT 102.545 114.385 103.210 114.555 ;
        RECT 101.155 113.525 102.285 113.695 ;
        RECT 102.460 113.565 102.810 114.215 ;
        RECT 100.645 113.160 101.310 113.335 ;
        RECT 100.620 112.555 100.955 112.980 ;
        RECT 101.125 112.755 101.310 113.160 ;
        RECT 101.515 112.555 101.845 113.335 ;
        RECT 102.015 112.755 102.285 113.525 ;
        RECT 102.980 113.395 103.210 114.385 ;
        RECT 102.545 113.225 103.210 113.395 ;
        RECT 102.545 112.725 102.715 113.225 ;
        RECT 102.885 112.555 103.215 113.055 ;
        RECT 103.385 112.725 103.570 114.845 ;
        RECT 103.825 114.645 104.075 115.105 ;
        RECT 104.245 114.655 104.580 114.825 ;
        RECT 104.775 114.655 105.450 114.825 ;
        RECT 104.245 114.515 104.415 114.655 ;
        RECT 103.740 113.525 104.020 114.475 ;
        RECT 104.190 114.385 104.415 114.515 ;
        RECT 104.190 113.280 104.360 114.385 ;
        RECT 104.585 114.235 105.110 114.455 ;
        RECT 104.530 113.470 104.770 114.065 ;
        RECT 104.940 113.535 105.110 114.235 ;
        RECT 105.280 113.875 105.450 114.655 ;
        RECT 105.770 114.605 106.140 115.105 ;
        RECT 106.320 114.655 106.725 114.825 ;
        RECT 106.895 114.655 107.680 114.825 ;
        RECT 106.320 114.425 106.490 114.655 ;
        RECT 105.660 114.125 106.490 114.425 ;
        RECT 106.875 114.155 107.340 114.485 ;
        RECT 105.660 114.095 105.860 114.125 ;
        RECT 105.980 113.875 106.150 113.945 ;
        RECT 105.280 113.705 106.150 113.875 ;
        RECT 105.640 113.615 106.150 113.705 ;
        RECT 104.190 113.150 104.495 113.280 ;
        RECT 104.940 113.170 105.470 113.535 ;
        RECT 103.810 112.555 104.075 113.015 ;
        RECT 104.245 112.725 104.495 113.150 ;
        RECT 105.640 113.000 105.810 113.615 ;
        RECT 104.705 112.830 105.810 113.000 ;
        RECT 105.980 112.555 106.150 113.355 ;
        RECT 106.320 113.055 106.490 114.125 ;
        RECT 106.660 113.225 106.850 113.945 ;
        RECT 107.020 113.195 107.340 114.155 ;
        RECT 107.510 114.195 107.680 114.655 ;
        RECT 107.955 114.575 108.165 115.105 ;
        RECT 108.425 114.365 108.755 114.890 ;
        RECT 108.925 114.495 109.095 115.105 ;
        RECT 109.265 114.450 109.595 114.885 ;
        RECT 109.265 114.365 109.645 114.450 ;
        RECT 108.555 114.195 108.755 114.365 ;
        RECT 109.420 114.325 109.645 114.365 ;
        RECT 109.820 114.340 110.275 115.105 ;
        RECT 110.550 114.725 111.850 114.935 ;
        RECT 112.105 114.745 112.435 115.105 ;
        RECT 111.680 114.575 111.850 114.725 ;
        RECT 112.605 114.605 112.865 114.935 ;
        RECT 112.635 114.595 112.865 114.605 ;
        RECT 107.510 113.865 108.385 114.195 ;
        RECT 108.555 113.865 109.305 114.195 ;
        RECT 106.320 112.725 106.570 113.055 ;
        RECT 107.510 113.025 107.680 113.865 ;
        RECT 108.555 113.660 108.745 113.865 ;
        RECT 109.475 113.745 109.645 114.325 ;
        RECT 110.750 114.115 110.970 114.515 ;
        RECT 109.815 113.915 110.305 114.115 ;
        RECT 110.495 113.905 110.970 114.115 ;
        RECT 111.215 114.115 111.425 114.515 ;
        RECT 111.680 114.450 112.435 114.575 ;
        RECT 111.680 114.405 112.525 114.450 ;
        RECT 112.255 114.285 112.525 114.405 ;
        RECT 111.215 113.905 111.545 114.115 ;
        RECT 111.715 113.845 112.125 114.150 ;
        RECT 109.430 113.695 109.645 113.745 ;
        RECT 107.850 113.285 108.745 113.660 ;
        RECT 109.255 113.615 109.645 113.695 ;
        RECT 109.820 113.675 110.995 113.735 ;
        RECT 112.355 113.710 112.525 114.285 ;
        RECT 112.325 113.675 112.525 113.710 ;
        RECT 106.795 112.855 107.680 113.025 ;
        RECT 107.860 112.555 108.175 113.055 ;
        RECT 108.405 112.725 108.745 113.285 ;
        RECT 108.915 112.555 109.085 113.565 ;
        RECT 109.255 112.770 109.585 113.615 ;
        RECT 109.820 113.565 112.525 113.675 ;
        RECT 109.820 112.945 110.075 113.565 ;
        RECT 110.665 113.505 112.465 113.565 ;
        RECT 110.665 113.475 110.995 113.505 ;
        RECT 112.695 113.405 112.865 114.595 ;
        RECT 113.035 114.560 118.380 115.105 ;
        RECT 114.620 113.730 114.960 114.560 ;
        RECT 118.555 114.335 120.225 115.105 ;
        RECT 120.395 114.380 120.685 115.105 ;
        RECT 120.855 114.355 122.065 115.105 ;
        RECT 122.325 114.555 122.495 114.845 ;
        RECT 122.665 114.725 122.995 115.105 ;
        RECT 122.325 114.385 122.990 114.555 ;
        RECT 110.325 113.305 110.510 113.395 ;
        RECT 111.100 113.305 111.935 113.315 ;
        RECT 110.325 113.105 111.935 113.305 ;
        RECT 110.325 113.065 110.555 113.105 ;
        RECT 109.820 112.725 110.155 112.945 ;
        RECT 111.160 112.555 111.515 112.935 ;
        RECT 111.685 112.725 111.935 113.105 ;
        RECT 112.185 112.555 112.435 113.335 ;
        RECT 112.605 112.725 112.865 113.405 ;
        RECT 116.440 112.990 116.790 114.240 ;
        RECT 118.555 113.815 119.305 114.335 ;
        RECT 119.475 113.645 120.225 114.165 ;
        RECT 120.855 113.815 121.375 114.355 ;
        RECT 113.035 112.555 118.380 112.990 ;
        RECT 118.555 112.555 120.225 113.645 ;
        RECT 120.395 112.555 120.685 113.720 ;
        RECT 121.545 113.645 122.065 114.185 ;
        RECT 120.855 112.555 122.065 113.645 ;
        RECT 122.240 113.565 122.590 114.215 ;
        RECT 122.760 113.395 122.990 114.385 ;
        RECT 122.325 113.225 122.990 113.395 ;
        RECT 122.325 112.725 122.495 113.225 ;
        RECT 122.665 112.555 122.995 113.055 ;
        RECT 123.165 112.725 123.350 114.845 ;
        RECT 123.605 114.645 123.855 115.105 ;
        RECT 124.025 114.655 124.360 114.825 ;
        RECT 124.555 114.655 125.230 114.825 ;
        RECT 124.025 114.515 124.195 114.655 ;
        RECT 123.520 113.525 123.800 114.475 ;
        RECT 123.970 114.385 124.195 114.515 ;
        RECT 123.970 113.280 124.140 114.385 ;
        RECT 124.365 114.235 124.890 114.455 ;
        RECT 124.310 113.470 124.550 114.065 ;
        RECT 124.720 113.535 124.890 114.235 ;
        RECT 125.060 113.875 125.230 114.655 ;
        RECT 125.550 114.605 125.920 115.105 ;
        RECT 126.100 114.655 126.505 114.825 ;
        RECT 126.675 114.655 127.460 114.825 ;
        RECT 126.100 114.425 126.270 114.655 ;
        RECT 125.440 114.125 126.270 114.425 ;
        RECT 126.655 114.155 127.120 114.485 ;
        RECT 125.440 114.095 125.640 114.125 ;
        RECT 125.760 113.875 125.930 113.945 ;
        RECT 125.060 113.705 125.930 113.875 ;
        RECT 125.420 113.615 125.930 113.705 ;
        RECT 123.970 113.150 124.275 113.280 ;
        RECT 124.720 113.170 125.250 113.535 ;
        RECT 123.590 112.555 123.855 113.015 ;
        RECT 124.025 112.725 124.275 113.150 ;
        RECT 125.420 113.000 125.590 113.615 ;
        RECT 124.485 112.830 125.590 113.000 ;
        RECT 125.760 112.555 125.930 113.355 ;
        RECT 126.100 113.055 126.270 114.125 ;
        RECT 126.440 113.225 126.630 113.945 ;
        RECT 126.800 113.195 127.120 114.155 ;
        RECT 127.290 114.195 127.460 114.655 ;
        RECT 127.735 114.575 127.945 115.105 ;
        RECT 128.205 114.365 128.535 114.890 ;
        RECT 128.705 114.495 128.875 115.105 ;
        RECT 129.045 114.450 129.375 114.885 ;
        RECT 129.045 114.365 129.425 114.450 ;
        RECT 128.335 114.195 128.535 114.365 ;
        RECT 129.200 114.325 129.425 114.365 ;
        RECT 127.290 113.865 128.165 114.195 ;
        RECT 128.335 113.865 129.085 114.195 ;
        RECT 126.100 112.725 126.350 113.055 ;
        RECT 127.290 113.025 127.460 113.865 ;
        RECT 128.335 113.660 128.525 113.865 ;
        RECT 129.255 113.745 129.425 114.325 ;
        RECT 129.210 113.695 129.425 113.745 ;
        RECT 127.630 113.285 128.525 113.660 ;
        RECT 129.035 113.615 129.425 113.695 ;
        RECT 129.600 114.365 129.855 114.935 ;
        RECT 130.025 114.705 130.355 115.105 ;
        RECT 130.780 114.570 131.310 114.935 ;
        RECT 131.500 114.765 131.775 114.935 ;
        RECT 131.495 114.595 131.775 114.765 ;
        RECT 130.780 114.535 130.955 114.570 ;
        RECT 130.025 114.365 130.955 114.535 ;
        RECT 129.600 113.695 129.770 114.365 ;
        RECT 130.025 114.195 130.195 114.365 ;
        RECT 129.940 113.865 130.195 114.195 ;
        RECT 130.420 113.865 130.615 114.195 ;
        RECT 126.575 112.855 127.460 113.025 ;
        RECT 127.640 112.555 127.955 113.055 ;
        RECT 128.185 112.725 128.525 113.285 ;
        RECT 128.695 112.555 128.865 113.565 ;
        RECT 129.035 112.770 129.365 113.615 ;
        RECT 129.600 112.725 129.935 113.695 ;
        RECT 130.105 112.555 130.275 113.695 ;
        RECT 130.445 112.895 130.615 113.865 ;
        RECT 130.785 113.235 130.955 114.365 ;
        RECT 131.125 113.575 131.295 114.375 ;
        RECT 131.500 113.775 131.775 114.595 ;
        RECT 131.945 113.575 132.135 114.935 ;
        RECT 132.315 114.570 132.825 115.105 ;
        RECT 133.045 114.295 133.290 114.900 ;
        RECT 133.735 114.335 135.405 115.105 ;
        RECT 135.580 114.365 135.835 114.935 ;
        RECT 136.005 114.705 136.335 115.105 ;
        RECT 136.760 114.570 137.290 114.935 ;
        RECT 137.480 114.765 137.755 114.935 ;
        RECT 137.475 114.595 137.755 114.765 ;
        RECT 136.760 114.535 136.935 114.570 ;
        RECT 136.005 114.365 136.935 114.535 ;
        RECT 132.335 114.125 133.565 114.295 ;
        RECT 131.125 113.405 132.135 113.575 ;
        RECT 132.305 113.560 133.055 113.750 ;
        RECT 130.785 113.065 131.910 113.235 ;
        RECT 132.305 112.895 132.475 113.560 ;
        RECT 133.225 113.315 133.565 114.125 ;
        RECT 133.735 113.815 134.485 114.335 ;
        RECT 134.655 113.645 135.405 114.165 ;
        RECT 130.445 112.725 132.475 112.895 ;
        RECT 132.645 112.555 132.815 113.315 ;
        RECT 133.050 112.905 133.565 113.315 ;
        RECT 133.735 112.555 135.405 113.645 ;
        RECT 135.580 113.695 135.750 114.365 ;
        RECT 136.005 114.195 136.175 114.365 ;
        RECT 135.920 113.865 136.175 114.195 ;
        RECT 136.400 113.865 136.595 114.195 ;
        RECT 135.580 112.725 135.915 113.695 ;
        RECT 136.085 112.555 136.255 113.695 ;
        RECT 136.425 112.895 136.595 113.865 ;
        RECT 136.765 113.235 136.935 114.365 ;
        RECT 137.105 113.575 137.275 114.375 ;
        RECT 137.480 113.775 137.755 114.595 ;
        RECT 137.925 113.575 138.115 114.935 ;
        RECT 138.295 114.570 138.805 115.105 ;
        RECT 139.025 114.295 139.270 114.900 ;
        RECT 139.720 114.365 139.975 114.935 ;
        RECT 140.145 114.705 140.475 115.105 ;
        RECT 140.900 114.570 141.430 114.935 ;
        RECT 140.900 114.535 141.075 114.570 ;
        RECT 140.145 114.365 141.075 114.535 ;
        RECT 138.315 114.125 139.545 114.295 ;
        RECT 137.105 113.405 138.115 113.575 ;
        RECT 138.285 113.560 139.035 113.750 ;
        RECT 136.765 113.065 137.890 113.235 ;
        RECT 138.285 112.895 138.455 113.560 ;
        RECT 139.205 113.315 139.545 114.125 ;
        RECT 136.425 112.725 138.455 112.895 ;
        RECT 138.625 112.555 138.795 113.315 ;
        RECT 139.030 112.905 139.545 113.315 ;
        RECT 139.720 113.695 139.890 114.365 ;
        RECT 140.145 114.195 140.315 114.365 ;
        RECT 140.060 113.865 140.315 114.195 ;
        RECT 140.540 113.865 140.735 114.195 ;
        RECT 139.720 112.725 140.055 113.695 ;
        RECT 140.225 112.555 140.395 113.695 ;
        RECT 140.565 112.895 140.735 113.865 ;
        RECT 140.905 113.235 141.075 114.365 ;
        RECT 141.245 113.575 141.415 114.375 ;
        RECT 141.620 114.085 141.895 114.935 ;
        RECT 141.615 113.915 141.895 114.085 ;
        RECT 141.620 113.775 141.895 113.915 ;
        RECT 142.065 113.575 142.255 114.935 ;
        RECT 142.435 114.570 142.945 115.105 ;
        RECT 143.165 114.295 143.410 114.900 ;
        RECT 143.945 114.555 144.115 114.935 ;
        RECT 144.330 114.725 144.660 115.105 ;
        RECT 143.945 114.385 144.660 114.555 ;
        RECT 142.455 114.125 143.685 114.295 ;
        RECT 141.245 113.405 142.255 113.575 ;
        RECT 142.425 113.560 143.175 113.750 ;
        RECT 140.905 113.065 142.030 113.235 ;
        RECT 142.425 112.895 142.595 113.560 ;
        RECT 143.345 113.315 143.685 114.125 ;
        RECT 143.855 113.835 144.210 114.205 ;
        RECT 144.490 114.195 144.660 114.385 ;
        RECT 144.830 114.360 145.085 114.935 ;
        RECT 144.490 113.865 144.745 114.195 ;
        RECT 144.490 113.655 144.660 113.865 ;
        RECT 140.565 112.725 142.595 112.895 ;
        RECT 142.765 112.555 142.935 113.315 ;
        RECT 143.170 112.905 143.685 113.315 ;
        RECT 143.945 113.485 144.660 113.655 ;
        RECT 144.915 113.630 145.085 114.360 ;
        RECT 145.260 114.265 145.520 115.105 ;
        RECT 145.695 114.355 146.905 115.105 ;
        RECT 143.945 112.725 144.115 113.485 ;
        RECT 144.330 112.555 144.660 113.315 ;
        RECT 144.830 112.725 145.085 113.630 ;
        RECT 145.260 112.555 145.520 113.705 ;
        RECT 145.695 113.645 146.215 114.185 ;
        RECT 146.385 113.815 146.905 114.355 ;
        RECT 145.695 112.555 146.905 113.645 ;
        RECT 17.270 112.385 146.990 112.555 ;
        RECT 17.355 111.295 18.565 112.385 ;
        RECT 19.255 111.325 19.585 112.170 ;
        RECT 19.755 111.375 19.925 112.385 ;
        RECT 20.095 111.655 20.435 112.215 ;
        RECT 20.665 111.885 20.980 112.385 ;
        RECT 21.160 111.915 22.045 112.085 ;
        RECT 17.355 110.585 17.875 111.125 ;
        RECT 18.045 110.755 18.565 111.295 ;
        RECT 19.195 111.245 19.585 111.325 ;
        RECT 20.095 111.280 20.990 111.655 ;
        RECT 19.195 111.195 19.410 111.245 ;
        RECT 19.195 110.615 19.365 111.195 ;
        RECT 20.095 111.075 20.285 111.280 ;
        RECT 21.160 111.075 21.330 111.915 ;
        RECT 22.270 111.885 22.520 112.215 ;
        RECT 19.535 110.745 20.285 111.075 ;
        RECT 20.455 110.745 21.330 111.075 ;
        RECT 17.355 109.835 18.565 110.585 ;
        RECT 19.195 110.575 19.420 110.615 ;
        RECT 20.085 110.575 20.285 110.745 ;
        RECT 19.195 110.490 19.575 110.575 ;
        RECT 19.245 110.055 19.575 110.490 ;
        RECT 19.745 109.835 19.915 110.445 ;
        RECT 20.085 110.050 20.415 110.575 ;
        RECT 20.675 109.835 20.885 110.365 ;
        RECT 21.160 110.285 21.330 110.745 ;
        RECT 21.500 110.785 21.820 111.745 ;
        RECT 21.990 110.995 22.180 111.715 ;
        RECT 22.350 110.815 22.520 111.885 ;
        RECT 22.690 111.585 22.860 112.385 ;
        RECT 23.030 111.940 24.135 112.110 ;
        RECT 23.030 111.325 23.200 111.940 ;
        RECT 24.345 111.790 24.595 112.215 ;
        RECT 24.765 111.925 25.030 112.385 ;
        RECT 23.370 111.405 23.900 111.770 ;
        RECT 24.345 111.660 24.650 111.790 ;
        RECT 22.690 111.235 23.200 111.325 ;
        RECT 22.690 111.065 23.560 111.235 ;
        RECT 22.690 110.995 22.860 111.065 ;
        RECT 22.980 110.815 23.180 110.845 ;
        RECT 21.500 110.455 21.965 110.785 ;
        RECT 22.350 110.515 23.180 110.815 ;
        RECT 22.350 110.285 22.520 110.515 ;
        RECT 21.160 110.115 21.945 110.285 ;
        RECT 22.115 110.115 22.520 110.285 ;
        RECT 22.700 109.835 23.070 110.335 ;
        RECT 23.390 110.285 23.560 111.065 ;
        RECT 23.730 110.705 23.900 111.405 ;
        RECT 24.070 110.875 24.310 111.470 ;
        RECT 23.730 110.485 24.255 110.705 ;
        RECT 24.480 110.555 24.650 111.660 ;
        RECT 24.425 110.425 24.650 110.555 ;
        RECT 24.820 110.465 25.100 111.415 ;
        RECT 24.425 110.285 24.595 110.425 ;
        RECT 23.390 110.115 24.065 110.285 ;
        RECT 24.260 110.115 24.595 110.285 ;
        RECT 24.765 109.835 25.015 110.295 ;
        RECT 25.270 110.095 25.455 112.215 ;
        RECT 25.625 111.885 25.955 112.385 ;
        RECT 26.125 111.715 26.295 112.215 ;
        RECT 25.630 111.545 26.295 111.715 ;
        RECT 25.630 110.555 25.860 111.545 ;
        RECT 26.030 110.725 26.380 111.375 ;
        RECT 26.555 111.295 30.065 112.385 ;
        RECT 26.555 110.605 28.205 111.125 ;
        RECT 28.375 110.775 30.065 111.295 ;
        RECT 30.235 111.220 30.525 112.385 ;
        RECT 30.700 111.245 31.035 112.215 ;
        RECT 31.205 111.245 31.375 112.385 ;
        RECT 31.545 112.045 33.575 112.215 ;
        RECT 25.630 110.385 26.295 110.555 ;
        RECT 25.625 109.835 25.955 110.215 ;
        RECT 26.125 110.095 26.295 110.385 ;
        RECT 26.555 109.835 30.065 110.605 ;
        RECT 30.700 110.575 30.870 111.245 ;
        RECT 31.545 111.075 31.715 112.045 ;
        RECT 31.040 110.745 31.295 111.075 ;
        RECT 31.520 110.745 31.715 111.075 ;
        RECT 31.885 111.705 33.010 111.875 ;
        RECT 31.125 110.575 31.295 110.745 ;
        RECT 31.885 110.575 32.055 111.705 ;
        RECT 30.235 109.835 30.525 110.560 ;
        RECT 30.700 110.005 30.955 110.575 ;
        RECT 31.125 110.405 32.055 110.575 ;
        RECT 32.225 111.365 33.235 111.535 ;
        RECT 32.225 110.565 32.395 111.365 ;
        RECT 32.600 111.025 32.875 111.165 ;
        RECT 32.595 110.855 32.875 111.025 ;
        RECT 31.880 110.370 32.055 110.405 ;
        RECT 31.125 109.835 31.455 110.235 ;
        RECT 31.880 110.005 32.410 110.370 ;
        RECT 32.600 110.005 32.875 110.855 ;
        RECT 33.045 110.005 33.235 111.365 ;
        RECT 33.405 111.380 33.575 112.045 ;
        RECT 33.745 111.625 33.915 112.385 ;
        RECT 34.150 111.625 34.665 112.035 ;
        RECT 34.835 111.950 40.180 112.385 ;
        RECT 40.355 111.950 45.700 112.385 ;
        RECT 45.875 111.950 51.220 112.385 ;
        RECT 33.405 111.190 34.155 111.380 ;
        RECT 34.325 110.815 34.665 111.625 ;
        RECT 33.435 110.645 34.665 110.815 ;
        RECT 33.415 109.835 33.925 110.370 ;
        RECT 34.145 110.040 34.390 110.645 ;
        RECT 36.420 110.380 36.760 111.210 ;
        RECT 38.240 110.700 38.590 111.950 ;
        RECT 41.940 110.380 42.280 111.210 ;
        RECT 43.760 110.700 44.110 111.950 ;
        RECT 47.460 110.380 47.800 111.210 ;
        RECT 49.280 110.700 49.630 111.950 ;
        RECT 51.395 111.295 54.905 112.385 ;
        RECT 51.395 110.605 53.045 111.125 ;
        RECT 53.215 110.775 54.905 111.295 ;
        RECT 55.995 111.220 56.285 112.385 ;
        RECT 56.455 111.950 61.800 112.385 ;
        RECT 34.835 109.835 40.180 110.380 ;
        RECT 40.355 109.835 45.700 110.380 ;
        RECT 45.875 109.835 51.220 110.380 ;
        RECT 51.395 109.835 54.905 110.605 ;
        RECT 55.995 109.835 56.285 110.560 ;
        RECT 58.040 110.380 58.380 111.210 ;
        RECT 59.860 110.700 60.210 111.950 ;
        RECT 61.975 111.295 63.185 112.385 ;
        RECT 63.445 111.715 63.615 112.215 ;
        RECT 63.785 111.885 64.115 112.385 ;
        RECT 63.445 111.545 64.110 111.715 ;
        RECT 61.975 110.585 62.495 111.125 ;
        RECT 62.665 110.755 63.185 111.295 ;
        RECT 63.360 110.725 63.710 111.375 ;
        RECT 56.455 109.835 61.800 110.380 ;
        RECT 61.975 109.835 63.185 110.585 ;
        RECT 63.880 110.555 64.110 111.545 ;
        RECT 63.445 110.385 64.110 110.555 ;
        RECT 63.445 110.095 63.615 110.385 ;
        RECT 63.785 109.835 64.115 110.215 ;
        RECT 64.285 110.095 64.470 112.215 ;
        RECT 64.710 111.925 64.975 112.385 ;
        RECT 65.145 111.790 65.395 112.215 ;
        RECT 65.605 111.940 66.710 112.110 ;
        RECT 65.090 111.660 65.395 111.790 ;
        RECT 64.640 110.465 64.920 111.415 ;
        RECT 65.090 110.555 65.260 111.660 ;
        RECT 65.430 110.875 65.670 111.470 ;
        RECT 65.840 111.405 66.370 111.770 ;
        RECT 65.840 110.705 66.010 111.405 ;
        RECT 66.540 111.325 66.710 111.940 ;
        RECT 66.880 111.585 67.050 112.385 ;
        RECT 67.220 111.885 67.470 112.215 ;
        RECT 67.695 111.915 68.580 112.085 ;
        RECT 66.540 111.235 67.050 111.325 ;
        RECT 65.090 110.425 65.315 110.555 ;
        RECT 65.485 110.485 66.010 110.705 ;
        RECT 66.180 111.065 67.050 111.235 ;
        RECT 64.725 109.835 64.975 110.295 ;
        RECT 65.145 110.285 65.315 110.425 ;
        RECT 66.180 110.285 66.350 111.065 ;
        RECT 66.880 110.995 67.050 111.065 ;
        RECT 66.560 110.815 66.760 110.845 ;
        RECT 67.220 110.815 67.390 111.885 ;
        RECT 67.560 110.995 67.750 111.715 ;
        RECT 66.560 110.515 67.390 110.815 ;
        RECT 67.920 110.785 68.240 111.745 ;
        RECT 65.145 110.115 65.480 110.285 ;
        RECT 65.675 110.115 66.350 110.285 ;
        RECT 66.670 109.835 67.040 110.335 ;
        RECT 67.220 110.285 67.390 110.515 ;
        RECT 67.775 110.455 68.240 110.785 ;
        RECT 68.410 111.075 68.580 111.915 ;
        RECT 68.760 111.885 69.075 112.385 ;
        RECT 69.305 111.655 69.645 112.215 ;
        RECT 68.750 111.280 69.645 111.655 ;
        RECT 69.815 111.375 69.985 112.385 ;
        RECT 69.455 111.075 69.645 111.280 ;
        RECT 70.155 111.325 70.485 112.170 ;
        RECT 70.155 111.245 70.545 111.325 ;
        RECT 70.330 111.195 70.545 111.245 ;
        RECT 68.410 110.745 69.285 111.075 ;
        RECT 69.455 110.745 70.205 111.075 ;
        RECT 68.410 110.285 68.580 110.745 ;
        RECT 69.455 110.575 69.655 110.745 ;
        RECT 70.375 110.615 70.545 111.195 ;
        RECT 70.320 110.575 70.545 110.615 ;
        RECT 67.220 110.115 67.625 110.285 ;
        RECT 67.795 110.115 68.580 110.285 ;
        RECT 68.855 109.835 69.065 110.365 ;
        RECT 69.325 110.050 69.655 110.575 ;
        RECT 70.165 110.490 70.545 110.575 ;
        RECT 70.720 111.245 71.055 112.215 ;
        RECT 71.225 111.245 71.395 112.385 ;
        RECT 71.565 112.045 73.595 112.215 ;
        RECT 70.720 110.575 70.890 111.245 ;
        RECT 71.565 111.075 71.735 112.045 ;
        RECT 71.060 110.745 71.315 111.075 ;
        RECT 71.540 110.745 71.735 111.075 ;
        RECT 71.905 111.705 73.030 111.875 ;
        RECT 71.145 110.575 71.315 110.745 ;
        RECT 71.905 110.575 72.075 111.705 ;
        RECT 69.825 109.835 69.995 110.445 ;
        RECT 70.165 110.055 70.495 110.490 ;
        RECT 70.720 110.005 70.975 110.575 ;
        RECT 71.145 110.405 72.075 110.575 ;
        RECT 72.245 111.365 73.255 111.535 ;
        RECT 72.245 110.565 72.415 111.365 ;
        RECT 72.620 111.025 72.895 111.165 ;
        RECT 72.615 110.855 72.895 111.025 ;
        RECT 71.900 110.370 72.075 110.405 ;
        RECT 71.145 109.835 71.475 110.235 ;
        RECT 71.900 110.005 72.430 110.370 ;
        RECT 72.620 110.005 72.895 110.855 ;
        RECT 73.065 110.005 73.255 111.365 ;
        RECT 73.425 111.380 73.595 112.045 ;
        RECT 73.765 111.625 73.935 112.385 ;
        RECT 74.170 111.625 74.685 112.035 ;
        RECT 74.855 111.950 80.200 112.385 ;
        RECT 73.425 111.190 74.175 111.380 ;
        RECT 74.345 110.815 74.685 111.625 ;
        RECT 73.455 110.645 74.685 110.815 ;
        RECT 73.435 109.835 73.945 110.370 ;
        RECT 74.165 110.040 74.410 110.645 ;
        RECT 76.440 110.380 76.780 111.210 ;
        RECT 78.260 110.700 78.610 111.950 ;
        RECT 80.375 111.295 81.585 112.385 ;
        RECT 80.375 110.585 80.895 111.125 ;
        RECT 81.065 110.755 81.585 111.295 ;
        RECT 81.755 111.220 82.045 112.385 ;
        RECT 82.305 111.765 82.475 112.195 ;
        RECT 82.645 111.935 82.975 112.385 ;
        RECT 82.305 111.535 82.980 111.765 ;
        RECT 74.855 109.835 80.200 110.380 ;
        RECT 80.375 109.835 81.585 110.585 ;
        RECT 81.755 109.835 82.045 110.560 ;
        RECT 82.275 110.515 82.575 111.365 ;
        RECT 82.745 110.885 82.980 111.535 ;
        RECT 83.150 111.225 83.435 112.170 ;
        RECT 83.615 111.915 84.300 112.385 ;
        RECT 83.610 111.395 84.305 111.705 ;
        RECT 84.480 111.330 84.785 112.115 ;
        RECT 83.150 111.075 84.010 111.225 ;
        RECT 83.150 111.055 84.435 111.075 ;
        RECT 82.745 110.555 83.280 110.885 ;
        RECT 83.450 110.695 84.435 111.055 ;
        RECT 82.745 110.405 82.965 110.555 ;
        RECT 82.220 109.835 82.555 110.340 ;
        RECT 82.725 110.030 82.965 110.405 ;
        RECT 83.450 110.360 83.620 110.695 ;
        RECT 84.610 110.525 84.785 111.330 ;
        RECT 84.975 111.295 88.485 112.385 ;
        RECT 83.245 110.165 83.620 110.360 ;
        RECT 83.245 110.020 83.415 110.165 ;
        RECT 83.980 109.835 84.375 110.330 ;
        RECT 84.545 110.005 84.785 110.525 ;
        RECT 84.975 110.605 86.625 111.125 ;
        RECT 86.795 110.775 88.485 111.295 ;
        RECT 88.655 111.535 88.915 112.215 ;
        RECT 89.085 111.605 89.335 112.385 ;
        RECT 89.585 111.835 89.835 112.215 ;
        RECT 90.005 112.005 90.360 112.385 ;
        RECT 91.365 111.995 91.700 112.215 ;
        RECT 90.965 111.835 91.195 111.875 ;
        RECT 89.585 111.635 91.195 111.835 ;
        RECT 89.585 111.625 90.420 111.635 ;
        RECT 91.010 111.545 91.195 111.635 ;
        RECT 84.975 109.835 88.485 110.605 ;
        RECT 88.655 110.335 88.825 111.535 ;
        RECT 90.525 111.435 90.855 111.465 ;
        RECT 89.055 111.375 90.855 111.435 ;
        RECT 91.445 111.375 91.700 111.995 ;
        RECT 91.875 111.950 97.220 112.385 ;
        RECT 97.395 111.950 102.740 112.385 ;
        RECT 88.995 111.265 91.700 111.375 ;
        RECT 88.995 111.230 89.195 111.265 ;
        RECT 88.995 110.655 89.165 111.230 ;
        RECT 90.525 111.205 91.700 111.265 ;
        RECT 89.395 110.790 89.805 111.095 ;
        RECT 89.975 110.825 90.305 111.035 ;
        RECT 88.995 110.535 89.265 110.655 ;
        RECT 88.995 110.490 89.840 110.535 ;
        RECT 89.085 110.365 89.840 110.490 ;
        RECT 90.095 110.425 90.305 110.825 ;
        RECT 90.550 110.825 91.025 111.035 ;
        RECT 91.215 110.825 91.705 111.025 ;
        RECT 90.550 110.425 90.770 110.825 ;
        RECT 88.655 110.005 88.915 110.335 ;
        RECT 89.670 110.215 89.840 110.365 ;
        RECT 89.085 109.835 89.415 110.195 ;
        RECT 89.670 110.005 90.970 110.215 ;
        RECT 91.245 109.835 91.700 110.600 ;
        RECT 93.460 110.380 93.800 111.210 ;
        RECT 95.280 110.700 95.630 111.950 ;
        RECT 98.980 110.380 99.320 111.210 ;
        RECT 100.800 110.700 101.150 111.950 ;
        RECT 102.935 111.330 103.240 112.115 ;
        RECT 103.420 111.915 104.105 112.385 ;
        RECT 103.415 111.395 104.110 111.705 ;
        RECT 102.935 110.525 103.110 111.330 ;
        RECT 104.285 111.225 104.570 112.170 ;
        RECT 104.745 111.935 105.075 112.385 ;
        RECT 105.245 111.765 105.415 112.195 ;
        RECT 103.710 111.075 104.570 111.225 ;
        RECT 103.285 111.055 104.570 111.075 ;
        RECT 104.740 111.535 105.415 111.765 ;
        RECT 103.285 110.695 104.270 111.055 ;
        RECT 104.740 110.885 104.975 111.535 ;
        RECT 91.875 109.835 97.220 110.380 ;
        RECT 97.395 109.835 102.740 110.380 ;
        RECT 102.935 110.005 103.175 110.525 ;
        RECT 104.100 110.360 104.270 110.695 ;
        RECT 104.440 110.555 104.975 110.885 ;
        RECT 104.755 110.405 104.975 110.555 ;
        RECT 105.145 110.515 105.445 111.365 ;
        RECT 105.675 111.295 107.345 112.385 ;
        RECT 105.675 110.605 106.425 111.125 ;
        RECT 106.595 110.775 107.345 111.295 ;
        RECT 107.515 111.220 107.805 112.385 ;
        RECT 108.065 111.765 108.235 112.195 ;
        RECT 108.405 111.935 108.735 112.385 ;
        RECT 108.065 111.535 108.740 111.765 ;
        RECT 103.345 109.835 103.740 110.330 ;
        RECT 104.100 110.165 104.475 110.360 ;
        RECT 104.305 110.020 104.475 110.165 ;
        RECT 104.755 110.030 104.995 110.405 ;
        RECT 105.165 109.835 105.500 110.340 ;
        RECT 105.675 109.835 107.345 110.605 ;
        RECT 107.515 109.835 107.805 110.560 ;
        RECT 108.035 110.515 108.335 111.365 ;
        RECT 108.505 110.885 108.740 111.535 ;
        RECT 108.910 111.225 109.195 112.170 ;
        RECT 109.375 111.915 110.060 112.385 ;
        RECT 109.370 111.395 110.065 111.705 ;
        RECT 110.240 111.330 110.545 112.115 ;
        RECT 108.910 111.075 109.770 111.225 ;
        RECT 108.910 111.055 110.195 111.075 ;
        RECT 108.505 110.555 109.040 110.885 ;
        RECT 109.210 110.695 110.195 111.055 ;
        RECT 108.505 110.405 108.725 110.555 ;
        RECT 107.980 109.835 108.315 110.340 ;
        RECT 108.485 110.030 108.725 110.405 ;
        RECT 109.210 110.360 109.380 110.695 ;
        RECT 110.370 110.525 110.545 111.330 ;
        RECT 110.735 111.295 112.405 112.385 ;
        RECT 109.005 110.165 109.380 110.360 ;
        RECT 109.005 110.020 109.175 110.165 ;
        RECT 109.740 109.835 110.135 110.330 ;
        RECT 110.305 110.005 110.545 110.525 ;
        RECT 110.735 110.605 111.485 111.125 ;
        RECT 111.655 110.775 112.405 111.295 ;
        RECT 113.035 111.625 113.550 112.035 ;
        RECT 113.785 111.625 113.955 112.385 ;
        RECT 114.125 112.045 116.155 112.215 ;
        RECT 113.035 110.815 113.375 111.625 ;
        RECT 114.125 111.380 114.295 112.045 ;
        RECT 114.690 111.705 115.815 111.875 ;
        RECT 113.545 111.190 114.295 111.380 ;
        RECT 114.465 111.365 115.475 111.535 ;
        RECT 113.035 110.645 114.265 110.815 ;
        RECT 110.735 109.835 112.405 110.605 ;
        RECT 113.310 110.040 113.555 110.645 ;
        RECT 113.775 109.835 114.285 110.370 ;
        RECT 114.465 110.005 114.655 111.365 ;
        RECT 114.825 111.025 115.100 111.165 ;
        RECT 114.825 110.855 115.105 111.025 ;
        RECT 114.825 110.005 115.100 110.855 ;
        RECT 115.305 110.565 115.475 111.365 ;
        RECT 115.645 110.575 115.815 111.705 ;
        RECT 115.985 111.075 116.155 112.045 ;
        RECT 116.325 111.245 116.495 112.385 ;
        RECT 116.665 111.245 117.000 112.215 ;
        RECT 117.265 111.715 117.435 112.215 ;
        RECT 117.605 111.885 117.935 112.385 ;
        RECT 117.265 111.545 117.930 111.715 ;
        RECT 115.985 110.745 116.180 111.075 ;
        RECT 116.405 110.745 116.660 111.075 ;
        RECT 116.405 110.575 116.575 110.745 ;
        RECT 116.830 110.575 117.000 111.245 ;
        RECT 117.180 110.725 117.530 111.375 ;
        RECT 115.645 110.405 116.575 110.575 ;
        RECT 115.645 110.370 115.820 110.405 ;
        RECT 115.290 110.005 115.820 110.370 ;
        RECT 116.245 109.835 116.575 110.235 ;
        RECT 116.745 110.005 117.000 110.575 ;
        RECT 117.700 110.555 117.930 111.545 ;
        RECT 117.265 110.385 117.930 110.555 ;
        RECT 117.265 110.095 117.435 110.385 ;
        RECT 117.605 109.835 117.935 110.215 ;
        RECT 118.105 110.095 118.290 112.215 ;
        RECT 118.530 111.925 118.795 112.385 ;
        RECT 118.965 111.790 119.215 112.215 ;
        RECT 119.425 111.940 120.530 112.110 ;
        RECT 118.910 111.660 119.215 111.790 ;
        RECT 118.460 110.465 118.740 111.415 ;
        RECT 118.910 110.555 119.080 111.660 ;
        RECT 119.250 110.875 119.490 111.470 ;
        RECT 119.660 111.405 120.190 111.770 ;
        RECT 119.660 110.705 119.830 111.405 ;
        RECT 120.360 111.325 120.530 111.940 ;
        RECT 120.700 111.585 120.870 112.385 ;
        RECT 121.040 111.885 121.290 112.215 ;
        RECT 121.515 111.915 122.400 112.085 ;
        RECT 120.360 111.235 120.870 111.325 ;
        RECT 118.910 110.425 119.135 110.555 ;
        RECT 119.305 110.485 119.830 110.705 ;
        RECT 120.000 111.065 120.870 111.235 ;
        RECT 118.545 109.835 118.795 110.295 ;
        RECT 118.965 110.285 119.135 110.425 ;
        RECT 120.000 110.285 120.170 111.065 ;
        RECT 120.700 110.995 120.870 111.065 ;
        RECT 120.380 110.815 120.580 110.845 ;
        RECT 121.040 110.815 121.210 111.885 ;
        RECT 121.380 110.995 121.570 111.715 ;
        RECT 120.380 110.515 121.210 110.815 ;
        RECT 121.740 110.785 122.060 111.745 ;
        RECT 118.965 110.115 119.300 110.285 ;
        RECT 119.495 110.115 120.170 110.285 ;
        RECT 120.490 109.835 120.860 110.335 ;
        RECT 121.040 110.285 121.210 110.515 ;
        RECT 121.595 110.455 122.060 110.785 ;
        RECT 122.230 111.075 122.400 111.915 ;
        RECT 122.580 111.885 122.895 112.385 ;
        RECT 123.125 111.655 123.465 112.215 ;
        RECT 122.570 111.280 123.465 111.655 ;
        RECT 123.635 111.375 123.805 112.385 ;
        RECT 123.275 111.075 123.465 111.280 ;
        RECT 123.975 111.325 124.305 112.170 ;
        RECT 124.535 111.950 129.880 112.385 ;
        RECT 123.975 111.245 124.365 111.325 ;
        RECT 124.150 111.195 124.365 111.245 ;
        RECT 122.230 110.745 123.105 111.075 ;
        RECT 123.275 110.745 124.025 111.075 ;
        RECT 122.230 110.285 122.400 110.745 ;
        RECT 123.275 110.575 123.475 110.745 ;
        RECT 124.195 110.615 124.365 111.195 ;
        RECT 124.140 110.575 124.365 110.615 ;
        RECT 121.040 110.115 121.445 110.285 ;
        RECT 121.615 110.115 122.400 110.285 ;
        RECT 122.675 109.835 122.885 110.365 ;
        RECT 123.145 110.050 123.475 110.575 ;
        RECT 123.985 110.490 124.365 110.575 ;
        RECT 123.645 109.835 123.815 110.445 ;
        RECT 123.985 110.055 124.315 110.490 ;
        RECT 126.120 110.380 126.460 111.210 ;
        RECT 127.940 110.700 128.290 111.950 ;
        RECT 130.605 111.765 130.775 112.195 ;
        RECT 130.945 111.935 131.275 112.385 ;
        RECT 130.605 111.535 131.280 111.765 ;
        RECT 130.575 110.515 130.875 111.365 ;
        RECT 131.045 110.885 131.280 111.535 ;
        RECT 131.450 111.225 131.735 112.170 ;
        RECT 131.915 111.915 132.600 112.385 ;
        RECT 131.910 111.395 132.605 111.705 ;
        RECT 132.780 111.330 133.085 112.115 ;
        RECT 131.450 111.075 132.310 111.225 ;
        RECT 131.450 111.055 132.735 111.075 ;
        RECT 131.045 110.555 131.580 110.885 ;
        RECT 131.750 110.695 132.735 111.055 ;
        RECT 131.045 110.405 131.265 110.555 ;
        RECT 124.535 109.835 129.880 110.380 ;
        RECT 130.520 109.835 130.855 110.340 ;
        RECT 131.025 110.030 131.265 110.405 ;
        RECT 131.750 110.360 131.920 110.695 ;
        RECT 132.910 110.525 133.085 111.330 ;
        RECT 133.275 111.220 133.565 112.385 ;
        RECT 133.735 111.295 135.405 112.385 ;
        RECT 136.125 111.715 136.295 112.215 ;
        RECT 136.465 111.885 136.795 112.385 ;
        RECT 136.125 111.545 136.790 111.715 ;
        RECT 133.735 110.605 134.485 111.125 ;
        RECT 134.655 110.775 135.405 111.295 ;
        RECT 136.040 110.725 136.390 111.375 ;
        RECT 131.545 110.165 131.920 110.360 ;
        RECT 131.545 110.020 131.715 110.165 ;
        RECT 132.280 109.835 132.675 110.330 ;
        RECT 132.845 110.005 133.085 110.525 ;
        RECT 133.275 109.835 133.565 110.560 ;
        RECT 133.735 109.835 135.405 110.605 ;
        RECT 136.560 110.555 136.790 111.545 ;
        RECT 136.125 110.385 136.790 110.555 ;
        RECT 136.125 110.095 136.295 110.385 ;
        RECT 136.465 109.835 136.795 110.215 ;
        RECT 136.965 110.095 137.150 112.215 ;
        RECT 137.390 111.925 137.655 112.385 ;
        RECT 137.825 111.790 138.075 112.215 ;
        RECT 138.285 111.940 139.390 112.110 ;
        RECT 137.770 111.660 138.075 111.790 ;
        RECT 137.320 110.465 137.600 111.415 ;
        RECT 137.770 110.555 137.940 111.660 ;
        RECT 138.110 110.875 138.350 111.470 ;
        RECT 138.520 111.405 139.050 111.770 ;
        RECT 138.520 110.705 138.690 111.405 ;
        RECT 139.220 111.325 139.390 111.940 ;
        RECT 139.560 111.585 139.730 112.385 ;
        RECT 139.900 111.885 140.150 112.215 ;
        RECT 140.375 111.915 141.260 112.085 ;
        RECT 139.220 111.235 139.730 111.325 ;
        RECT 137.770 110.425 137.995 110.555 ;
        RECT 138.165 110.485 138.690 110.705 ;
        RECT 138.860 111.065 139.730 111.235 ;
        RECT 137.405 109.835 137.655 110.295 ;
        RECT 137.825 110.285 137.995 110.425 ;
        RECT 138.860 110.285 139.030 111.065 ;
        RECT 139.560 110.995 139.730 111.065 ;
        RECT 139.240 110.815 139.440 110.845 ;
        RECT 139.900 110.815 140.070 111.885 ;
        RECT 140.240 110.995 140.430 111.715 ;
        RECT 139.240 110.515 140.070 110.815 ;
        RECT 140.600 110.785 140.920 111.745 ;
        RECT 137.825 110.115 138.160 110.285 ;
        RECT 138.355 110.115 139.030 110.285 ;
        RECT 139.350 109.835 139.720 110.335 ;
        RECT 139.900 110.285 140.070 110.515 ;
        RECT 140.455 110.455 140.920 110.785 ;
        RECT 141.090 111.075 141.260 111.915 ;
        RECT 141.440 111.885 141.755 112.385 ;
        RECT 141.985 111.655 142.325 112.215 ;
        RECT 141.430 111.280 142.325 111.655 ;
        RECT 142.495 111.375 142.665 112.385 ;
        RECT 142.135 111.075 142.325 111.280 ;
        RECT 142.835 111.325 143.165 112.170 ;
        RECT 143.945 111.455 144.115 112.215 ;
        RECT 144.330 111.625 144.660 112.385 ;
        RECT 142.835 111.245 143.225 111.325 ;
        RECT 143.945 111.285 144.660 111.455 ;
        RECT 144.830 111.310 145.085 112.215 ;
        RECT 143.010 111.195 143.225 111.245 ;
        RECT 141.090 110.745 141.965 111.075 ;
        RECT 142.135 110.745 142.885 111.075 ;
        RECT 141.090 110.285 141.260 110.745 ;
        RECT 142.135 110.575 142.335 110.745 ;
        RECT 143.055 110.615 143.225 111.195 ;
        RECT 143.855 110.735 144.210 111.105 ;
        RECT 144.490 111.075 144.660 111.285 ;
        RECT 144.490 110.745 144.745 111.075 ;
        RECT 143.000 110.575 143.225 110.615 ;
        RECT 139.900 110.115 140.305 110.285 ;
        RECT 140.475 110.115 141.260 110.285 ;
        RECT 141.535 109.835 141.745 110.365 ;
        RECT 142.005 110.050 142.335 110.575 ;
        RECT 142.845 110.490 143.225 110.575 ;
        RECT 144.490 110.555 144.660 110.745 ;
        RECT 144.915 110.580 145.085 111.310 ;
        RECT 145.260 111.235 145.520 112.385 ;
        RECT 145.695 111.295 146.905 112.385 ;
        RECT 145.695 110.755 146.215 111.295 ;
        RECT 142.505 109.835 142.675 110.445 ;
        RECT 142.845 110.055 143.175 110.490 ;
        RECT 143.945 110.385 144.660 110.555 ;
        RECT 143.945 110.005 144.115 110.385 ;
        RECT 144.330 109.835 144.660 110.215 ;
        RECT 144.830 110.005 145.085 110.580 ;
        RECT 145.260 109.835 145.520 110.675 ;
        RECT 146.385 110.585 146.905 111.125 ;
        RECT 145.695 109.835 146.905 110.585 ;
        RECT 17.270 109.665 146.990 109.835 ;
        RECT 17.355 108.915 18.565 109.665 ;
        RECT 17.355 108.375 17.875 108.915 ;
        RECT 18.740 108.825 19.000 109.665 ;
        RECT 19.175 108.920 19.430 109.495 ;
        RECT 19.600 109.285 19.930 109.665 ;
        RECT 20.145 109.115 20.315 109.495 ;
        RECT 19.600 108.945 20.315 109.115 ;
        RECT 21.085 109.010 21.415 109.445 ;
        RECT 21.585 109.055 21.755 109.665 ;
        RECT 18.045 108.205 18.565 108.745 ;
        RECT 17.355 107.115 18.565 108.205 ;
        RECT 18.740 107.115 19.000 108.265 ;
        RECT 19.175 108.190 19.345 108.920 ;
        RECT 19.600 108.755 19.770 108.945 ;
        RECT 21.035 108.925 21.415 109.010 ;
        RECT 21.925 108.925 22.255 109.450 ;
        RECT 22.515 109.135 22.725 109.665 ;
        RECT 23.000 109.215 23.785 109.385 ;
        RECT 23.955 109.215 24.360 109.385 ;
        RECT 21.035 108.885 21.260 108.925 ;
        RECT 19.515 108.425 19.770 108.755 ;
        RECT 19.600 108.215 19.770 108.425 ;
        RECT 20.050 108.395 20.405 108.765 ;
        RECT 21.035 108.305 21.205 108.885 ;
        RECT 21.925 108.755 22.125 108.925 ;
        RECT 23.000 108.755 23.170 109.215 ;
        RECT 21.375 108.425 22.125 108.755 ;
        RECT 22.295 108.425 23.170 108.755 ;
        RECT 21.035 108.255 21.250 108.305 ;
        RECT 19.175 107.285 19.430 108.190 ;
        RECT 19.600 108.045 20.315 108.215 ;
        RECT 21.035 108.175 21.425 108.255 ;
        RECT 19.600 107.115 19.930 107.875 ;
        RECT 20.145 107.285 20.315 108.045 ;
        RECT 21.095 107.330 21.425 108.175 ;
        RECT 21.935 108.220 22.125 108.425 ;
        RECT 21.595 107.115 21.765 108.125 ;
        RECT 21.935 107.845 22.830 108.220 ;
        RECT 21.935 107.285 22.275 107.845 ;
        RECT 22.505 107.115 22.820 107.615 ;
        RECT 23.000 107.585 23.170 108.425 ;
        RECT 23.340 108.715 23.805 109.045 ;
        RECT 24.190 108.985 24.360 109.215 ;
        RECT 24.540 109.165 24.910 109.665 ;
        RECT 25.230 109.215 25.905 109.385 ;
        RECT 26.100 109.215 26.435 109.385 ;
        RECT 23.340 107.755 23.660 108.715 ;
        RECT 24.190 108.685 25.020 108.985 ;
        RECT 23.830 107.785 24.020 108.505 ;
        RECT 24.190 107.615 24.360 108.685 ;
        RECT 24.820 108.655 25.020 108.685 ;
        RECT 24.530 108.435 24.700 108.505 ;
        RECT 25.230 108.435 25.400 109.215 ;
        RECT 26.265 109.075 26.435 109.215 ;
        RECT 26.605 109.205 26.855 109.665 ;
        RECT 24.530 108.265 25.400 108.435 ;
        RECT 25.570 108.795 26.095 109.015 ;
        RECT 26.265 108.945 26.490 109.075 ;
        RECT 24.530 108.175 25.040 108.265 ;
        RECT 23.000 107.415 23.885 107.585 ;
        RECT 24.110 107.285 24.360 107.615 ;
        RECT 24.530 107.115 24.700 107.915 ;
        RECT 24.870 107.560 25.040 108.175 ;
        RECT 25.570 108.095 25.740 108.795 ;
        RECT 25.210 107.730 25.740 108.095 ;
        RECT 25.910 108.030 26.150 108.625 ;
        RECT 26.320 107.840 26.490 108.945 ;
        RECT 26.660 108.085 26.940 109.035 ;
        RECT 26.185 107.710 26.490 107.840 ;
        RECT 24.870 107.390 25.975 107.560 ;
        RECT 26.185 107.285 26.435 107.710 ;
        RECT 26.605 107.115 26.870 107.575 ;
        RECT 27.110 107.285 27.295 109.405 ;
        RECT 27.465 109.285 27.795 109.665 ;
        RECT 27.965 109.115 28.135 109.405 ;
        RECT 27.470 108.945 28.135 109.115 ;
        RECT 27.470 107.955 27.700 108.945 ;
        RECT 28.400 108.925 28.655 109.495 ;
        RECT 28.825 109.265 29.155 109.665 ;
        RECT 29.580 109.130 30.110 109.495 ;
        RECT 29.580 109.095 29.755 109.130 ;
        RECT 28.825 108.925 29.755 109.095 ;
        RECT 30.300 108.985 30.575 109.495 ;
        RECT 27.870 108.125 28.220 108.775 ;
        RECT 28.400 108.255 28.570 108.925 ;
        RECT 28.825 108.755 28.995 108.925 ;
        RECT 28.740 108.425 28.995 108.755 ;
        RECT 29.220 108.425 29.415 108.755 ;
        RECT 27.470 107.785 28.135 107.955 ;
        RECT 27.465 107.115 27.795 107.615 ;
        RECT 27.965 107.285 28.135 107.785 ;
        RECT 28.400 107.285 28.735 108.255 ;
        RECT 28.905 107.115 29.075 108.255 ;
        RECT 29.245 107.455 29.415 108.425 ;
        RECT 29.585 107.795 29.755 108.925 ;
        RECT 29.925 108.135 30.095 108.935 ;
        RECT 30.295 108.815 30.575 108.985 ;
        RECT 30.300 108.335 30.575 108.815 ;
        RECT 30.745 108.135 30.935 109.495 ;
        RECT 31.115 109.130 31.625 109.665 ;
        RECT 31.845 108.855 32.090 109.460 ;
        RECT 32.535 109.120 37.880 109.665 ;
        RECT 31.135 108.685 32.365 108.855 ;
        RECT 29.925 107.965 30.935 108.135 ;
        RECT 31.105 108.120 31.855 108.310 ;
        RECT 29.585 107.625 30.710 107.795 ;
        RECT 31.105 107.455 31.275 108.120 ;
        RECT 32.025 107.875 32.365 108.685 ;
        RECT 34.120 108.290 34.460 109.120 ;
        RECT 38.055 108.895 41.565 109.665 ;
        RECT 41.735 108.915 42.945 109.665 ;
        RECT 43.115 108.940 43.405 109.665 ;
        RECT 43.575 109.120 48.920 109.665 ;
        RECT 49.095 109.120 54.440 109.665 ;
        RECT 54.615 109.120 59.960 109.665 ;
        RECT 29.245 107.285 31.275 107.455 ;
        RECT 31.445 107.115 31.615 107.875 ;
        RECT 31.850 107.465 32.365 107.875 ;
        RECT 35.940 107.550 36.290 108.800 ;
        RECT 38.055 108.375 39.705 108.895 ;
        RECT 39.875 108.205 41.565 108.725 ;
        RECT 41.735 108.375 42.255 108.915 ;
        RECT 42.425 108.205 42.945 108.745 ;
        RECT 45.160 108.290 45.500 109.120 ;
        RECT 32.535 107.115 37.880 107.550 ;
        RECT 38.055 107.115 41.565 108.205 ;
        RECT 41.735 107.115 42.945 108.205 ;
        RECT 43.115 107.115 43.405 108.280 ;
        RECT 46.980 107.550 47.330 108.800 ;
        RECT 50.680 108.290 51.020 109.120 ;
        RECT 52.500 107.550 52.850 108.800 ;
        RECT 56.200 108.290 56.540 109.120 ;
        RECT 60.135 108.895 63.645 109.665 ;
        RECT 64.295 108.975 64.535 109.495 ;
        RECT 64.705 109.170 65.100 109.665 ;
        RECT 65.665 109.335 65.835 109.480 ;
        RECT 65.460 109.140 65.835 109.335 ;
        RECT 58.020 107.550 58.370 108.800 ;
        RECT 60.135 108.375 61.785 108.895 ;
        RECT 61.955 108.205 63.645 108.725 ;
        RECT 43.575 107.115 48.920 107.550 ;
        RECT 49.095 107.115 54.440 107.550 ;
        RECT 54.615 107.115 59.960 107.550 ;
        RECT 60.135 107.115 63.645 108.205 ;
        RECT 64.295 108.170 64.470 108.975 ;
        RECT 65.460 108.805 65.630 109.140 ;
        RECT 66.115 109.095 66.355 109.470 ;
        RECT 66.525 109.160 66.860 109.665 ;
        RECT 66.115 108.945 66.335 109.095 ;
        RECT 64.645 108.445 65.630 108.805 ;
        RECT 65.800 108.615 66.335 108.945 ;
        RECT 64.645 108.425 65.930 108.445 ;
        RECT 65.070 108.275 65.930 108.425 ;
        RECT 64.295 107.385 64.600 108.170 ;
        RECT 64.775 107.795 65.470 108.105 ;
        RECT 64.780 107.115 65.465 107.585 ;
        RECT 65.645 107.330 65.930 108.275 ;
        RECT 66.100 107.965 66.335 108.615 ;
        RECT 66.505 108.135 66.805 108.985 ;
        RECT 67.035 108.895 68.705 109.665 ;
        RECT 68.875 108.940 69.165 109.665 ;
        RECT 69.335 109.120 74.680 109.665 ;
        RECT 74.855 109.120 80.200 109.665 ;
        RECT 80.375 109.120 85.720 109.665 ;
        RECT 85.895 109.120 91.240 109.665 ;
        RECT 67.035 108.375 67.785 108.895 ;
        RECT 67.955 108.205 68.705 108.725 ;
        RECT 70.920 108.290 71.260 109.120 ;
        RECT 66.100 107.735 66.775 107.965 ;
        RECT 66.105 107.115 66.435 107.565 ;
        RECT 66.605 107.305 66.775 107.735 ;
        RECT 67.035 107.115 68.705 108.205 ;
        RECT 68.875 107.115 69.165 108.280 ;
        RECT 72.740 107.550 73.090 108.800 ;
        RECT 76.440 108.290 76.780 109.120 ;
        RECT 78.260 107.550 78.610 108.800 ;
        RECT 81.960 108.290 82.300 109.120 ;
        RECT 83.780 107.550 84.130 108.800 ;
        RECT 87.480 108.290 87.820 109.120 ;
        RECT 91.415 108.895 94.005 109.665 ;
        RECT 94.635 108.940 94.925 109.665 ;
        RECT 95.095 109.120 100.440 109.665 ;
        RECT 100.615 109.120 105.960 109.665 ;
        RECT 107.060 109.160 107.395 109.665 ;
        RECT 89.300 107.550 89.650 108.800 ;
        RECT 91.415 108.375 92.625 108.895 ;
        RECT 92.795 108.205 94.005 108.725 ;
        RECT 96.680 108.290 97.020 109.120 ;
        RECT 69.335 107.115 74.680 107.550 ;
        RECT 74.855 107.115 80.200 107.550 ;
        RECT 80.375 107.115 85.720 107.550 ;
        RECT 85.895 107.115 91.240 107.550 ;
        RECT 91.415 107.115 94.005 108.205 ;
        RECT 94.635 107.115 94.925 108.280 ;
        RECT 98.500 107.550 98.850 108.800 ;
        RECT 102.200 108.290 102.540 109.120 ;
        RECT 107.565 109.095 107.805 109.470 ;
        RECT 108.085 109.335 108.255 109.480 ;
        RECT 108.085 109.140 108.460 109.335 ;
        RECT 108.820 109.170 109.215 109.665 ;
        RECT 104.020 107.550 104.370 108.800 ;
        RECT 107.115 108.135 107.415 108.985 ;
        RECT 107.585 108.945 107.805 109.095 ;
        RECT 107.585 108.615 108.120 108.945 ;
        RECT 108.290 108.805 108.460 109.140 ;
        RECT 109.385 108.975 109.625 109.495 ;
        RECT 109.815 109.120 115.160 109.665 ;
        RECT 116.260 109.160 116.595 109.665 ;
        RECT 107.585 107.965 107.820 108.615 ;
        RECT 108.290 108.445 109.275 108.805 ;
        RECT 107.145 107.735 107.820 107.965 ;
        RECT 107.990 108.425 109.275 108.445 ;
        RECT 107.990 108.275 108.850 108.425 ;
        RECT 95.095 107.115 100.440 107.550 ;
        RECT 100.615 107.115 105.960 107.550 ;
        RECT 107.145 107.305 107.315 107.735 ;
        RECT 107.485 107.115 107.815 107.565 ;
        RECT 107.990 107.330 108.275 108.275 ;
        RECT 109.450 108.170 109.625 108.975 ;
        RECT 111.400 108.290 111.740 109.120 ;
        RECT 116.765 109.095 117.005 109.470 ;
        RECT 117.285 109.335 117.455 109.480 ;
        RECT 117.285 109.140 117.660 109.335 ;
        RECT 118.020 109.170 118.415 109.665 ;
        RECT 108.450 107.795 109.145 108.105 ;
        RECT 108.455 107.115 109.140 107.585 ;
        RECT 109.320 107.385 109.625 108.170 ;
        RECT 113.220 107.550 113.570 108.800 ;
        RECT 116.315 108.135 116.615 108.985 ;
        RECT 116.785 108.945 117.005 109.095 ;
        RECT 116.785 108.615 117.320 108.945 ;
        RECT 117.490 108.805 117.660 109.140 ;
        RECT 118.585 108.975 118.825 109.495 ;
        RECT 116.785 107.965 117.020 108.615 ;
        RECT 117.490 108.445 118.475 108.805 ;
        RECT 116.345 107.735 117.020 107.965 ;
        RECT 117.190 108.425 118.475 108.445 ;
        RECT 117.190 108.275 118.050 108.425 ;
        RECT 109.815 107.115 115.160 107.550 ;
        RECT 116.345 107.305 116.515 107.735 ;
        RECT 116.685 107.115 117.015 107.565 ;
        RECT 117.190 107.330 117.475 108.275 ;
        RECT 118.650 108.170 118.825 108.975 ;
        RECT 119.015 108.915 120.225 109.665 ;
        RECT 120.395 108.940 120.685 109.665 ;
        RECT 120.855 109.120 126.200 109.665 ;
        RECT 126.375 109.120 131.720 109.665 ;
        RECT 119.015 108.375 119.535 108.915 ;
        RECT 119.705 108.205 120.225 108.745 ;
        RECT 122.440 108.290 122.780 109.120 ;
        RECT 117.650 107.795 118.345 108.105 ;
        RECT 117.655 107.115 118.340 107.585 ;
        RECT 118.520 107.385 118.825 108.170 ;
        RECT 119.015 107.115 120.225 108.205 ;
        RECT 120.395 107.115 120.685 108.280 ;
        RECT 124.260 107.550 124.610 108.800 ;
        RECT 127.960 108.290 128.300 109.120 ;
        RECT 131.895 108.895 133.565 109.665 ;
        RECT 133.740 109.160 134.075 109.665 ;
        RECT 134.245 109.095 134.485 109.470 ;
        RECT 134.765 109.335 134.935 109.480 ;
        RECT 134.765 109.140 135.140 109.335 ;
        RECT 135.500 109.170 135.895 109.665 ;
        RECT 129.780 107.550 130.130 108.800 ;
        RECT 131.895 108.375 132.645 108.895 ;
        RECT 132.815 108.205 133.565 108.725 ;
        RECT 120.855 107.115 126.200 107.550 ;
        RECT 126.375 107.115 131.720 107.550 ;
        RECT 131.895 107.115 133.565 108.205 ;
        RECT 133.795 108.135 134.095 108.985 ;
        RECT 134.265 108.945 134.485 109.095 ;
        RECT 134.265 108.615 134.800 108.945 ;
        RECT 134.970 108.805 135.140 109.140 ;
        RECT 136.065 108.975 136.305 109.495 ;
        RECT 134.265 107.965 134.500 108.615 ;
        RECT 134.970 108.445 135.955 108.805 ;
        RECT 133.825 107.735 134.500 107.965 ;
        RECT 134.670 108.425 135.955 108.445 ;
        RECT 134.670 108.275 135.530 108.425 ;
        RECT 133.825 107.305 133.995 107.735 ;
        RECT 134.165 107.115 134.495 107.565 ;
        RECT 134.670 107.330 134.955 108.275 ;
        RECT 136.130 108.170 136.305 108.975 ;
        RECT 136.585 109.115 136.755 109.405 ;
        RECT 136.925 109.285 137.255 109.665 ;
        RECT 136.585 108.945 137.250 109.115 ;
        RECT 135.130 107.795 135.825 108.105 ;
        RECT 135.135 107.115 135.820 107.585 ;
        RECT 136.000 107.385 136.305 108.170 ;
        RECT 136.500 108.125 136.850 108.775 ;
        RECT 137.020 107.955 137.250 108.945 ;
        RECT 136.585 107.785 137.250 107.955 ;
        RECT 136.585 107.285 136.755 107.785 ;
        RECT 136.925 107.115 137.255 107.615 ;
        RECT 137.425 107.285 137.610 109.405 ;
        RECT 137.865 109.205 138.115 109.665 ;
        RECT 138.285 109.215 138.620 109.385 ;
        RECT 138.815 109.215 139.490 109.385 ;
        RECT 138.285 109.075 138.455 109.215 ;
        RECT 137.780 108.085 138.060 109.035 ;
        RECT 138.230 108.945 138.455 109.075 ;
        RECT 138.230 107.840 138.400 108.945 ;
        RECT 138.625 108.795 139.150 109.015 ;
        RECT 138.570 108.030 138.810 108.625 ;
        RECT 138.980 108.095 139.150 108.795 ;
        RECT 139.320 108.435 139.490 109.215 ;
        RECT 139.810 109.165 140.180 109.665 ;
        RECT 140.360 109.215 140.765 109.385 ;
        RECT 140.935 109.215 141.720 109.385 ;
        RECT 140.360 108.985 140.530 109.215 ;
        RECT 139.700 108.685 140.530 108.985 ;
        RECT 140.915 108.715 141.380 109.045 ;
        RECT 139.700 108.655 139.900 108.685 ;
        RECT 140.020 108.435 140.190 108.505 ;
        RECT 139.320 108.265 140.190 108.435 ;
        RECT 139.680 108.175 140.190 108.265 ;
        RECT 138.230 107.710 138.535 107.840 ;
        RECT 138.980 107.730 139.510 108.095 ;
        RECT 137.850 107.115 138.115 107.575 ;
        RECT 138.285 107.285 138.535 107.710 ;
        RECT 139.680 107.560 139.850 108.175 ;
        RECT 138.745 107.390 139.850 107.560 ;
        RECT 140.020 107.115 140.190 107.915 ;
        RECT 140.360 107.615 140.530 108.685 ;
        RECT 140.700 107.785 140.890 108.505 ;
        RECT 141.060 107.755 141.380 108.715 ;
        RECT 141.550 108.755 141.720 109.215 ;
        RECT 141.995 109.135 142.205 109.665 ;
        RECT 142.465 108.925 142.795 109.450 ;
        RECT 142.965 109.055 143.135 109.665 ;
        RECT 143.305 109.010 143.635 109.445 ;
        RECT 143.945 109.115 144.115 109.495 ;
        RECT 144.330 109.285 144.660 109.665 ;
        RECT 143.305 108.925 143.685 109.010 ;
        RECT 143.945 108.945 144.660 109.115 ;
        RECT 142.595 108.755 142.795 108.925 ;
        RECT 143.460 108.885 143.685 108.925 ;
        RECT 141.550 108.425 142.425 108.755 ;
        RECT 142.595 108.425 143.345 108.755 ;
        RECT 140.360 107.285 140.610 107.615 ;
        RECT 141.550 107.585 141.720 108.425 ;
        RECT 142.595 108.220 142.785 108.425 ;
        RECT 143.515 108.305 143.685 108.885 ;
        RECT 143.855 108.395 144.210 108.765 ;
        RECT 144.490 108.755 144.660 108.945 ;
        RECT 144.830 108.920 145.085 109.495 ;
        RECT 144.490 108.425 144.745 108.755 ;
        RECT 143.470 108.255 143.685 108.305 ;
        RECT 141.890 107.845 142.785 108.220 ;
        RECT 143.295 108.175 143.685 108.255 ;
        RECT 144.490 108.215 144.660 108.425 ;
        RECT 140.835 107.415 141.720 107.585 ;
        RECT 141.900 107.115 142.215 107.615 ;
        RECT 142.445 107.285 142.785 107.845 ;
        RECT 142.955 107.115 143.125 108.125 ;
        RECT 143.295 107.330 143.625 108.175 ;
        RECT 143.945 108.045 144.660 108.215 ;
        RECT 144.915 108.190 145.085 108.920 ;
        RECT 145.260 108.825 145.520 109.665 ;
        RECT 145.695 108.915 146.905 109.665 ;
        RECT 143.945 107.285 144.115 108.045 ;
        RECT 144.330 107.115 144.660 107.875 ;
        RECT 144.830 107.285 145.085 108.190 ;
        RECT 145.260 107.115 145.520 108.265 ;
        RECT 145.695 108.205 146.215 108.745 ;
        RECT 146.385 108.375 146.905 108.915 ;
        RECT 145.695 107.115 146.905 108.205 ;
        RECT 17.270 106.945 146.990 107.115 ;
        RECT 17.355 105.855 18.565 106.945 ;
        RECT 19.255 105.885 19.585 106.730 ;
        RECT 19.755 105.935 19.925 106.945 ;
        RECT 20.095 106.215 20.435 106.775 ;
        RECT 20.665 106.445 20.980 106.945 ;
        RECT 21.160 106.475 22.045 106.645 ;
        RECT 17.355 105.145 17.875 105.685 ;
        RECT 18.045 105.315 18.565 105.855 ;
        RECT 19.195 105.805 19.585 105.885 ;
        RECT 20.095 105.840 20.990 106.215 ;
        RECT 19.195 105.755 19.410 105.805 ;
        RECT 19.195 105.175 19.365 105.755 ;
        RECT 20.095 105.635 20.285 105.840 ;
        RECT 21.160 105.635 21.330 106.475 ;
        RECT 22.270 106.445 22.520 106.775 ;
        RECT 19.535 105.305 20.285 105.635 ;
        RECT 20.455 105.305 21.330 105.635 ;
        RECT 17.355 104.395 18.565 105.145 ;
        RECT 19.195 105.135 19.420 105.175 ;
        RECT 20.085 105.135 20.285 105.305 ;
        RECT 19.195 105.050 19.575 105.135 ;
        RECT 19.245 104.615 19.575 105.050 ;
        RECT 19.745 104.395 19.915 105.005 ;
        RECT 20.085 104.610 20.415 105.135 ;
        RECT 20.675 104.395 20.885 104.925 ;
        RECT 21.160 104.845 21.330 105.305 ;
        RECT 21.500 105.345 21.820 106.305 ;
        RECT 21.990 105.555 22.180 106.275 ;
        RECT 22.350 105.375 22.520 106.445 ;
        RECT 22.690 106.145 22.860 106.945 ;
        RECT 23.030 106.500 24.135 106.670 ;
        RECT 23.030 105.885 23.200 106.500 ;
        RECT 24.345 106.350 24.595 106.775 ;
        RECT 24.765 106.485 25.030 106.945 ;
        RECT 23.370 105.965 23.900 106.330 ;
        RECT 24.345 106.220 24.650 106.350 ;
        RECT 22.690 105.795 23.200 105.885 ;
        RECT 22.690 105.625 23.560 105.795 ;
        RECT 22.690 105.555 22.860 105.625 ;
        RECT 22.980 105.375 23.180 105.405 ;
        RECT 21.500 105.015 21.965 105.345 ;
        RECT 22.350 105.075 23.180 105.375 ;
        RECT 22.350 104.845 22.520 105.075 ;
        RECT 21.160 104.675 21.945 104.845 ;
        RECT 22.115 104.675 22.520 104.845 ;
        RECT 22.700 104.395 23.070 104.895 ;
        RECT 23.390 104.845 23.560 105.625 ;
        RECT 23.730 105.265 23.900 105.965 ;
        RECT 24.070 105.435 24.310 106.030 ;
        RECT 23.730 105.045 24.255 105.265 ;
        RECT 24.480 105.115 24.650 106.220 ;
        RECT 24.425 104.985 24.650 105.115 ;
        RECT 24.820 105.025 25.100 105.975 ;
        RECT 24.425 104.845 24.595 104.985 ;
        RECT 23.390 104.675 24.065 104.845 ;
        RECT 24.260 104.675 24.595 104.845 ;
        RECT 24.765 104.395 25.015 104.855 ;
        RECT 25.270 104.655 25.455 106.775 ;
        RECT 25.625 106.445 25.955 106.945 ;
        RECT 26.125 106.275 26.295 106.775 ;
        RECT 25.630 106.105 26.295 106.275 ;
        RECT 25.630 105.115 25.860 106.105 ;
        RECT 26.030 105.285 26.380 105.935 ;
        RECT 26.555 105.855 27.765 106.945 ;
        RECT 26.555 105.145 27.075 105.685 ;
        RECT 27.245 105.315 27.765 105.855 ;
        RECT 27.940 105.805 28.215 106.775 ;
        RECT 28.425 106.145 28.705 106.945 ;
        RECT 28.875 106.435 30.065 106.725 ;
        RECT 28.875 106.095 30.045 106.265 ;
        RECT 28.875 105.975 29.045 106.095 ;
        RECT 28.385 105.805 29.045 105.975 ;
        RECT 25.630 104.945 26.295 105.115 ;
        RECT 25.625 104.395 25.955 104.775 ;
        RECT 26.125 104.655 26.295 104.945 ;
        RECT 26.555 104.395 27.765 105.145 ;
        RECT 27.940 105.070 28.110 105.805 ;
        RECT 28.385 105.635 28.555 105.805 ;
        RECT 29.355 105.635 29.550 105.925 ;
        RECT 29.720 105.805 30.045 106.095 ;
        RECT 30.235 105.780 30.525 106.945 ;
        RECT 30.695 105.790 31.035 106.775 ;
        RECT 31.205 106.515 31.615 106.945 ;
        RECT 32.360 106.525 32.690 106.945 ;
        RECT 32.860 106.345 33.185 106.775 ;
        RECT 31.205 106.175 33.185 106.345 ;
        RECT 28.280 105.305 28.555 105.635 ;
        RECT 28.725 105.305 29.550 105.635 ;
        RECT 29.720 105.305 30.065 105.635 ;
        RECT 28.385 105.135 28.555 105.305 ;
        RECT 30.695 105.135 30.950 105.790 ;
        RECT 31.205 105.635 31.470 106.175 ;
        RECT 31.685 105.835 32.310 106.005 ;
        RECT 31.120 105.305 31.470 105.635 ;
        RECT 31.640 105.305 31.970 105.635 ;
        RECT 32.140 105.135 32.310 105.835 ;
        RECT 27.940 104.725 28.215 105.070 ;
        RECT 28.385 104.965 30.050 105.135 ;
        RECT 28.405 104.395 28.785 104.795 ;
        RECT 28.955 104.615 29.125 104.965 ;
        RECT 29.295 104.395 29.625 104.795 ;
        RECT 29.795 104.615 30.050 104.965 ;
        RECT 30.235 104.395 30.525 105.120 ;
        RECT 30.695 104.760 31.055 105.135 ;
        RECT 31.320 104.395 31.490 105.135 ;
        RECT 31.770 104.965 32.310 105.135 ;
        RECT 32.480 105.765 33.185 106.175 ;
        RECT 33.660 105.845 33.990 106.945 ;
        RECT 34.380 106.435 36.035 106.725 ;
        RECT 34.380 106.095 35.970 106.265 ;
        RECT 36.205 106.145 36.485 106.945 ;
        RECT 34.380 105.805 34.700 106.095 ;
        RECT 35.800 105.975 35.970 106.095 ;
        RECT 31.770 104.760 31.940 104.965 ;
        RECT 32.480 104.565 32.650 105.765 ;
        RECT 34.895 105.755 35.610 105.925 ;
        RECT 35.800 105.805 36.525 105.975 ;
        RECT 36.695 105.805 36.965 106.775 ;
        RECT 37.135 106.510 42.480 106.945 ;
        RECT 42.655 106.510 48.000 106.945 ;
        RECT 48.175 106.510 53.520 106.945 ;
        RECT 32.820 105.385 33.390 105.595 ;
        RECT 33.560 105.385 34.205 105.595 ;
        RECT 32.880 105.045 34.050 105.215 ;
        RECT 34.380 105.065 34.730 105.635 ;
        RECT 34.900 105.305 35.610 105.755 ;
        RECT 36.355 105.635 36.525 105.805 ;
        RECT 35.780 105.305 36.185 105.635 ;
        RECT 36.355 105.305 36.625 105.635 ;
        RECT 36.355 105.135 36.525 105.305 ;
        RECT 32.880 104.565 33.210 105.045 ;
        RECT 33.380 104.395 33.550 104.865 ;
        RECT 33.720 104.580 34.050 105.045 ;
        RECT 34.915 104.965 36.525 105.135 ;
        RECT 36.795 105.070 36.965 105.805 ;
        RECT 34.385 104.395 34.715 104.895 ;
        RECT 34.915 104.615 35.085 104.965 ;
        RECT 35.285 104.395 35.615 104.795 ;
        RECT 35.785 104.615 35.955 104.965 ;
        RECT 36.125 104.395 36.505 104.795 ;
        RECT 36.695 104.725 36.965 105.070 ;
        RECT 38.720 104.940 39.060 105.770 ;
        RECT 40.540 105.260 40.890 106.510 ;
        RECT 44.240 104.940 44.580 105.770 ;
        RECT 46.060 105.260 46.410 106.510 ;
        RECT 49.760 104.940 50.100 105.770 ;
        RECT 51.580 105.260 51.930 106.510 ;
        RECT 53.695 105.855 55.365 106.945 ;
        RECT 53.695 105.165 54.445 105.685 ;
        RECT 54.615 105.335 55.365 105.855 ;
        RECT 55.995 105.780 56.285 106.945 ;
        RECT 56.455 106.510 61.800 106.945 ;
        RECT 37.135 104.395 42.480 104.940 ;
        RECT 42.655 104.395 48.000 104.940 ;
        RECT 48.175 104.395 53.520 104.940 ;
        RECT 53.695 104.395 55.365 105.165 ;
        RECT 55.995 104.395 56.285 105.120 ;
        RECT 58.040 104.940 58.380 105.770 ;
        RECT 59.860 105.260 60.210 106.510 ;
        RECT 62.065 106.325 62.235 106.755 ;
        RECT 62.405 106.495 62.735 106.945 ;
        RECT 62.065 106.095 62.740 106.325 ;
        RECT 62.035 105.075 62.335 105.925 ;
        RECT 62.505 105.445 62.740 106.095 ;
        RECT 62.910 105.785 63.195 106.730 ;
        RECT 63.375 106.475 64.060 106.945 ;
        RECT 63.370 105.955 64.065 106.265 ;
        RECT 64.240 105.890 64.545 106.675 ;
        RECT 62.910 105.635 63.770 105.785 ;
        RECT 62.910 105.615 64.195 105.635 ;
        RECT 62.505 105.115 63.040 105.445 ;
        RECT 63.210 105.255 64.195 105.615 ;
        RECT 62.505 104.965 62.725 105.115 ;
        RECT 56.455 104.395 61.800 104.940 ;
        RECT 61.980 104.395 62.315 104.900 ;
        RECT 62.485 104.590 62.725 104.965 ;
        RECT 63.210 104.920 63.380 105.255 ;
        RECT 64.370 105.085 64.545 105.890 ;
        RECT 64.735 105.855 67.325 106.945 ;
        RECT 63.005 104.725 63.380 104.920 ;
        RECT 63.005 104.580 63.175 104.725 ;
        RECT 63.740 104.395 64.135 104.890 ;
        RECT 64.305 104.565 64.545 105.085 ;
        RECT 64.735 105.165 65.945 105.685 ;
        RECT 66.115 105.335 67.325 105.855 ;
        RECT 67.500 105.805 67.835 106.775 ;
        RECT 68.005 105.805 68.175 106.945 ;
        RECT 68.345 106.605 70.375 106.775 ;
        RECT 64.735 104.395 67.325 105.165 ;
        RECT 67.500 105.135 67.670 105.805 ;
        RECT 68.345 105.635 68.515 106.605 ;
        RECT 67.840 105.305 68.095 105.635 ;
        RECT 68.320 105.305 68.515 105.635 ;
        RECT 68.685 106.265 69.810 106.435 ;
        RECT 67.925 105.135 68.095 105.305 ;
        RECT 68.685 105.135 68.855 106.265 ;
        RECT 67.500 104.565 67.755 105.135 ;
        RECT 67.925 104.965 68.855 105.135 ;
        RECT 69.025 105.925 70.035 106.095 ;
        RECT 69.025 105.125 69.195 105.925 ;
        RECT 69.400 105.245 69.675 105.725 ;
        RECT 69.395 105.075 69.675 105.245 ;
        RECT 68.680 104.930 68.855 104.965 ;
        RECT 67.925 104.395 68.255 104.795 ;
        RECT 68.680 104.565 69.210 104.930 ;
        RECT 69.400 104.565 69.675 105.075 ;
        RECT 69.845 104.565 70.035 105.925 ;
        RECT 70.205 105.940 70.375 106.605 ;
        RECT 70.545 106.185 70.715 106.945 ;
        RECT 70.950 106.185 71.465 106.595 ;
        RECT 70.205 105.750 70.955 105.940 ;
        RECT 71.125 105.375 71.465 106.185 ;
        RECT 71.640 106.555 71.975 106.775 ;
        RECT 72.980 106.565 73.335 106.945 ;
        RECT 71.640 105.935 71.895 106.555 ;
        RECT 72.145 106.395 72.375 106.435 ;
        RECT 73.505 106.395 73.755 106.775 ;
        RECT 72.145 106.195 73.755 106.395 ;
        RECT 72.145 106.105 72.330 106.195 ;
        RECT 72.920 106.185 73.755 106.195 ;
        RECT 74.005 106.165 74.255 106.945 ;
        RECT 74.425 106.095 74.685 106.775 ;
        RECT 72.485 105.995 72.815 106.025 ;
        RECT 72.485 105.935 74.285 105.995 ;
        RECT 71.640 105.825 74.345 105.935 ;
        RECT 71.640 105.765 72.815 105.825 ;
        RECT 74.145 105.790 74.345 105.825 ;
        RECT 71.635 105.385 72.125 105.585 ;
        RECT 72.315 105.385 72.790 105.595 ;
        RECT 70.235 105.205 71.465 105.375 ;
        RECT 70.215 104.395 70.725 104.930 ;
        RECT 70.945 104.600 71.190 105.205 ;
        RECT 71.640 104.395 72.095 105.160 ;
        RECT 72.570 104.985 72.790 105.385 ;
        RECT 73.035 105.385 73.365 105.595 ;
        RECT 73.035 104.985 73.245 105.385 ;
        RECT 73.535 105.350 73.945 105.655 ;
        RECT 74.175 105.215 74.345 105.790 ;
        RECT 74.075 105.095 74.345 105.215 ;
        RECT 73.500 105.050 74.345 105.095 ;
        RECT 73.500 104.925 74.255 105.050 ;
        RECT 73.500 104.775 73.670 104.925 ;
        RECT 74.515 104.895 74.685 106.095 ;
        RECT 74.855 105.855 78.365 106.945 ;
        RECT 79.085 106.325 79.255 106.755 ;
        RECT 79.425 106.495 79.755 106.945 ;
        RECT 79.085 106.095 79.760 106.325 ;
        RECT 72.370 104.565 73.670 104.775 ;
        RECT 73.925 104.395 74.255 104.755 ;
        RECT 74.425 104.565 74.685 104.895 ;
        RECT 74.855 105.165 76.505 105.685 ;
        RECT 76.675 105.335 78.365 105.855 ;
        RECT 74.855 104.395 78.365 105.165 ;
        RECT 79.055 105.075 79.355 105.925 ;
        RECT 79.525 105.445 79.760 106.095 ;
        RECT 79.930 105.785 80.215 106.730 ;
        RECT 80.395 106.475 81.080 106.945 ;
        RECT 80.390 105.955 81.085 106.265 ;
        RECT 81.260 105.890 81.565 106.675 ;
        RECT 79.930 105.635 80.790 105.785 ;
        RECT 79.930 105.615 81.215 105.635 ;
        RECT 79.525 105.115 80.060 105.445 ;
        RECT 80.230 105.255 81.215 105.615 ;
        RECT 79.525 104.965 79.745 105.115 ;
        RECT 79.000 104.395 79.335 104.900 ;
        RECT 79.505 104.590 79.745 104.965 ;
        RECT 80.230 104.920 80.400 105.255 ;
        RECT 81.390 105.085 81.565 105.890 ;
        RECT 81.755 105.780 82.045 106.945 ;
        RECT 82.215 105.855 83.885 106.945 ;
        RECT 82.215 105.165 82.965 105.685 ;
        RECT 83.135 105.335 83.885 105.855 ;
        RECT 84.060 105.805 84.395 106.775 ;
        RECT 84.565 105.805 84.735 106.945 ;
        RECT 84.905 106.605 86.935 106.775 ;
        RECT 80.025 104.725 80.400 104.920 ;
        RECT 80.025 104.580 80.195 104.725 ;
        RECT 80.760 104.395 81.155 104.890 ;
        RECT 81.325 104.565 81.565 105.085 ;
        RECT 81.755 104.395 82.045 105.120 ;
        RECT 82.215 104.395 83.885 105.165 ;
        RECT 84.060 105.135 84.230 105.805 ;
        RECT 84.905 105.635 85.075 106.605 ;
        RECT 84.400 105.305 84.655 105.635 ;
        RECT 84.880 105.305 85.075 105.635 ;
        RECT 85.245 106.265 86.370 106.435 ;
        RECT 84.485 105.135 84.655 105.305 ;
        RECT 85.245 105.135 85.415 106.265 ;
        RECT 84.060 104.565 84.315 105.135 ;
        RECT 84.485 104.965 85.415 105.135 ;
        RECT 85.585 105.925 86.595 106.095 ;
        RECT 85.585 105.125 85.755 105.925 ;
        RECT 85.240 104.930 85.415 104.965 ;
        RECT 84.485 104.395 84.815 104.795 ;
        RECT 85.240 104.565 85.770 104.930 ;
        RECT 85.960 104.905 86.235 105.725 ;
        RECT 85.955 104.735 86.235 104.905 ;
        RECT 85.960 104.565 86.235 104.735 ;
        RECT 86.405 104.565 86.595 105.925 ;
        RECT 86.765 105.940 86.935 106.605 ;
        RECT 87.105 106.185 87.275 106.945 ;
        RECT 87.510 106.185 88.025 106.595 ;
        RECT 86.765 105.750 87.515 105.940 ;
        RECT 87.685 105.375 88.025 106.185 ;
        RECT 88.195 105.855 89.865 106.945 ;
        RECT 86.795 105.205 88.025 105.375 ;
        RECT 86.775 104.395 87.285 104.930 ;
        RECT 87.505 104.600 87.750 105.205 ;
        RECT 88.195 105.165 88.945 105.685 ;
        RECT 89.115 105.335 89.865 105.855 ;
        RECT 90.585 105.935 90.755 106.775 ;
        RECT 90.925 106.605 92.095 106.775 ;
        RECT 90.925 106.105 91.255 106.605 ;
        RECT 91.765 106.565 92.095 106.605 ;
        RECT 92.285 106.525 92.640 106.945 ;
        RECT 91.425 106.345 91.655 106.435 ;
        RECT 92.810 106.345 93.060 106.775 ;
        RECT 91.425 106.105 93.060 106.345 ;
        RECT 93.230 106.185 93.560 106.945 ;
        RECT 93.730 106.105 93.985 106.775 ;
        RECT 90.585 105.765 93.645 105.935 ;
        RECT 90.500 105.385 90.850 105.595 ;
        RECT 91.020 105.385 91.465 105.585 ;
        RECT 91.635 105.385 92.110 105.585 ;
        RECT 88.195 104.395 89.865 105.165 ;
        RECT 90.585 105.045 91.650 105.215 ;
        RECT 90.585 104.565 90.755 105.045 ;
        RECT 90.925 104.395 91.255 104.875 ;
        RECT 91.480 104.815 91.650 105.045 ;
        RECT 91.830 104.985 92.110 105.385 ;
        RECT 92.380 105.385 92.710 105.585 ;
        RECT 92.880 105.385 93.245 105.585 ;
        RECT 92.380 104.985 92.665 105.385 ;
        RECT 93.475 105.215 93.645 105.765 ;
        RECT 92.845 105.045 93.645 105.215 ;
        RECT 92.845 104.815 93.015 105.045 ;
        RECT 93.815 104.975 93.985 106.105 ;
        RECT 94.175 105.855 95.385 106.945 ;
        RECT 93.800 104.905 93.985 104.975 ;
        RECT 93.775 104.895 93.985 104.905 ;
        RECT 91.480 104.565 93.015 104.815 ;
        RECT 93.185 104.395 93.515 104.875 ;
        RECT 93.730 104.565 93.985 104.895 ;
        RECT 94.175 105.145 94.695 105.685 ;
        RECT 94.865 105.315 95.385 105.855 ;
        RECT 95.555 105.975 95.825 106.745 ;
        RECT 95.995 106.165 96.325 106.945 ;
        RECT 96.530 106.340 96.715 106.745 ;
        RECT 96.885 106.520 97.220 106.945 ;
        RECT 96.530 106.165 97.195 106.340 ;
        RECT 95.555 105.805 96.685 105.975 ;
        RECT 94.175 104.395 95.385 105.145 ;
        RECT 95.555 104.895 95.725 105.805 ;
        RECT 95.895 105.055 96.255 105.635 ;
        RECT 96.435 105.305 96.685 105.805 ;
        RECT 96.855 105.135 97.195 106.165 ;
        RECT 96.510 104.965 97.195 105.135 ;
        RECT 97.395 105.805 97.655 106.775 ;
        RECT 97.825 106.520 98.210 106.945 ;
        RECT 98.380 106.350 98.635 106.775 ;
        RECT 97.825 106.155 98.635 106.350 ;
        RECT 97.395 105.135 97.580 105.805 ;
        RECT 97.825 105.635 98.175 106.155 ;
        RECT 98.825 105.985 99.070 106.775 ;
        RECT 99.240 106.520 99.625 106.945 ;
        RECT 99.795 106.350 100.070 106.775 ;
        RECT 97.750 105.305 98.175 105.635 ;
        RECT 98.345 105.805 99.070 105.985 ;
        RECT 99.240 106.155 100.070 106.350 ;
        RECT 98.345 105.305 98.995 105.805 ;
        RECT 99.240 105.635 99.590 106.155 ;
        RECT 100.240 105.985 100.665 106.775 ;
        RECT 100.835 106.520 101.220 106.945 ;
        RECT 101.390 106.350 101.825 106.775 ;
        RECT 99.165 105.305 99.590 105.635 ;
        RECT 99.760 105.805 100.665 105.985 ;
        RECT 100.835 106.180 101.825 106.350 ;
        RECT 99.760 105.305 100.590 105.805 ;
        RECT 100.835 105.635 101.170 106.180 ;
        RECT 100.760 105.305 101.170 105.635 ;
        RECT 101.340 105.305 101.825 106.010 ;
        RECT 102.000 105.805 102.335 106.775 ;
        RECT 102.505 105.805 102.675 106.945 ;
        RECT 102.845 106.605 104.875 106.775 ;
        RECT 97.825 105.135 98.175 105.305 ;
        RECT 98.825 105.135 98.995 105.305 ;
        RECT 99.240 105.135 99.590 105.305 ;
        RECT 100.240 105.135 100.590 105.305 ;
        RECT 100.835 105.135 101.170 105.305 ;
        RECT 102.000 105.135 102.170 105.805 ;
        RECT 102.845 105.635 103.015 106.605 ;
        RECT 102.340 105.305 102.595 105.635 ;
        RECT 102.820 105.305 103.015 105.635 ;
        RECT 103.185 106.265 104.310 106.435 ;
        RECT 102.425 105.135 102.595 105.305 ;
        RECT 103.185 105.135 103.355 106.265 ;
        RECT 95.555 104.565 95.815 104.895 ;
        RECT 96.025 104.395 96.300 104.875 ;
        RECT 96.510 104.565 96.715 104.965 ;
        RECT 96.885 104.395 97.220 104.795 ;
        RECT 97.395 104.565 97.655 105.135 ;
        RECT 97.825 104.965 98.635 105.135 ;
        RECT 97.825 104.395 98.210 104.795 ;
        RECT 98.380 104.565 98.635 104.965 ;
        RECT 98.825 104.565 99.070 105.135 ;
        RECT 99.240 104.965 100.050 105.135 ;
        RECT 99.240 104.395 99.625 104.795 ;
        RECT 99.795 104.565 100.050 104.965 ;
        RECT 100.240 104.565 100.665 105.135 ;
        RECT 100.835 104.965 101.825 105.135 ;
        RECT 100.835 104.395 101.220 104.795 ;
        RECT 101.390 104.565 101.825 104.965 ;
        RECT 102.000 104.565 102.255 105.135 ;
        RECT 102.425 104.965 103.355 105.135 ;
        RECT 103.525 105.925 104.535 106.095 ;
        RECT 103.525 105.125 103.695 105.925 ;
        RECT 103.900 105.245 104.175 105.725 ;
        RECT 103.895 105.075 104.175 105.245 ;
        RECT 103.180 104.930 103.355 104.965 ;
        RECT 102.425 104.395 102.755 104.795 ;
        RECT 103.180 104.565 103.710 104.930 ;
        RECT 103.900 104.565 104.175 105.075 ;
        RECT 104.345 104.565 104.535 105.925 ;
        RECT 104.705 105.940 104.875 106.605 ;
        RECT 105.045 106.185 105.215 106.945 ;
        RECT 105.450 106.185 105.965 106.595 ;
        RECT 104.705 105.750 105.455 105.940 ;
        RECT 105.625 105.375 105.965 106.185 ;
        RECT 106.135 105.855 107.345 106.945 ;
        RECT 104.735 105.205 105.965 105.375 ;
        RECT 104.715 104.395 105.225 104.930 ;
        RECT 105.445 104.600 105.690 105.205 ;
        RECT 106.135 105.145 106.655 105.685 ;
        RECT 106.825 105.315 107.345 105.855 ;
        RECT 107.515 105.780 107.805 106.945 ;
        RECT 108.440 105.805 108.775 106.775 ;
        RECT 108.945 105.805 109.115 106.945 ;
        RECT 109.285 106.605 111.315 106.775 ;
        RECT 106.135 104.395 107.345 105.145 ;
        RECT 108.440 105.135 108.610 105.805 ;
        RECT 109.285 105.635 109.455 106.605 ;
        RECT 108.780 105.305 109.035 105.635 ;
        RECT 109.260 105.305 109.455 105.635 ;
        RECT 109.625 106.265 110.750 106.435 ;
        RECT 108.865 105.135 109.035 105.305 ;
        RECT 109.625 105.135 109.795 106.265 ;
        RECT 107.515 104.395 107.805 105.120 ;
        RECT 108.440 104.565 108.695 105.135 ;
        RECT 108.865 104.965 109.795 105.135 ;
        RECT 109.965 105.925 110.975 106.095 ;
        RECT 109.965 105.125 110.135 105.925 ;
        RECT 109.620 104.930 109.795 104.965 ;
        RECT 108.865 104.395 109.195 104.795 ;
        RECT 109.620 104.565 110.150 104.930 ;
        RECT 110.340 104.905 110.615 105.725 ;
        RECT 110.335 104.735 110.615 104.905 ;
        RECT 110.340 104.565 110.615 104.735 ;
        RECT 110.785 104.565 110.975 105.925 ;
        RECT 111.145 105.940 111.315 106.605 ;
        RECT 111.485 106.185 111.655 106.945 ;
        RECT 111.890 106.185 112.405 106.595 ;
        RECT 111.145 105.750 111.895 105.940 ;
        RECT 112.065 105.375 112.405 106.185 ;
        RECT 112.575 105.855 114.245 106.945 ;
        RECT 111.175 105.205 112.405 105.375 ;
        RECT 111.155 104.395 111.665 104.930 ;
        RECT 111.885 104.600 112.130 105.205 ;
        RECT 112.575 105.165 113.325 105.685 ;
        RECT 113.495 105.335 114.245 105.855 ;
        RECT 114.505 105.935 114.675 106.775 ;
        RECT 114.845 106.605 116.015 106.775 ;
        RECT 114.845 106.105 115.175 106.605 ;
        RECT 115.685 106.565 116.015 106.605 ;
        RECT 116.205 106.525 116.560 106.945 ;
        RECT 115.345 106.345 115.575 106.435 ;
        RECT 116.730 106.345 116.980 106.775 ;
        RECT 115.345 106.105 116.980 106.345 ;
        RECT 117.150 106.185 117.480 106.945 ;
        RECT 117.650 106.105 117.905 106.775 ;
        RECT 118.095 106.510 123.440 106.945 ;
        RECT 114.505 105.765 117.565 105.935 ;
        RECT 114.420 105.385 114.770 105.595 ;
        RECT 114.940 105.385 115.385 105.585 ;
        RECT 115.555 105.385 116.030 105.585 ;
        RECT 112.575 104.395 114.245 105.165 ;
        RECT 114.505 105.045 115.570 105.215 ;
        RECT 114.505 104.565 114.675 105.045 ;
        RECT 114.845 104.395 115.175 104.875 ;
        RECT 115.400 104.815 115.570 105.045 ;
        RECT 115.750 104.985 116.030 105.385 ;
        RECT 116.300 105.385 116.630 105.585 ;
        RECT 116.800 105.385 117.165 105.585 ;
        RECT 116.300 104.985 116.585 105.385 ;
        RECT 117.395 105.215 117.565 105.765 ;
        RECT 116.765 105.045 117.565 105.215 ;
        RECT 116.765 104.815 116.935 105.045 ;
        RECT 117.735 104.975 117.905 106.105 ;
        RECT 117.720 104.895 117.905 104.975 ;
        RECT 119.680 104.940 120.020 105.770 ;
        RECT 121.500 105.260 121.850 106.510 ;
        RECT 123.615 105.855 126.205 106.945 ;
        RECT 126.465 106.325 126.635 106.755 ;
        RECT 126.805 106.495 127.135 106.945 ;
        RECT 126.465 106.095 127.140 106.325 ;
        RECT 123.615 105.165 124.825 105.685 ;
        RECT 124.995 105.335 126.205 105.855 ;
        RECT 115.400 104.565 116.935 104.815 ;
        RECT 117.105 104.395 117.435 104.875 ;
        RECT 117.650 104.565 117.905 104.895 ;
        RECT 118.095 104.395 123.440 104.940 ;
        RECT 123.615 104.395 126.205 105.165 ;
        RECT 126.435 105.075 126.735 105.925 ;
        RECT 126.905 105.445 127.140 106.095 ;
        RECT 127.310 105.785 127.595 106.730 ;
        RECT 127.775 106.475 128.460 106.945 ;
        RECT 127.770 105.955 128.465 106.265 ;
        RECT 128.640 105.890 128.945 106.675 ;
        RECT 127.310 105.635 128.170 105.785 ;
        RECT 127.310 105.615 128.595 105.635 ;
        RECT 126.905 105.115 127.440 105.445 ;
        RECT 127.610 105.255 128.595 105.615 ;
        RECT 126.905 104.965 127.125 105.115 ;
        RECT 126.380 104.395 126.715 104.900 ;
        RECT 126.885 104.590 127.125 104.965 ;
        RECT 127.610 104.920 127.780 105.255 ;
        RECT 128.770 105.085 128.945 105.890 ;
        RECT 127.405 104.725 127.780 104.920 ;
        RECT 127.405 104.580 127.575 104.725 ;
        RECT 128.140 104.395 128.535 104.890 ;
        RECT 128.705 104.565 128.945 105.085 ;
        RECT 129.135 105.975 129.405 106.745 ;
        RECT 129.575 106.165 129.905 106.945 ;
        RECT 130.110 106.340 130.295 106.745 ;
        RECT 130.465 106.520 130.800 106.945 ;
        RECT 130.980 106.520 131.315 106.945 ;
        RECT 131.485 106.340 131.670 106.745 ;
        RECT 130.110 106.165 130.775 106.340 ;
        RECT 129.135 105.805 130.265 105.975 ;
        RECT 129.135 104.895 129.305 105.805 ;
        RECT 129.475 105.055 129.835 105.635 ;
        RECT 130.015 105.305 130.265 105.805 ;
        RECT 130.435 105.135 130.775 106.165 ;
        RECT 130.090 104.965 130.775 105.135 ;
        RECT 131.005 106.165 131.670 106.340 ;
        RECT 131.875 106.165 132.205 106.945 ;
        RECT 131.005 105.135 131.345 106.165 ;
        RECT 132.375 105.975 132.645 106.745 ;
        RECT 131.515 105.805 132.645 105.975 ;
        RECT 131.515 105.305 131.765 105.805 ;
        RECT 131.005 104.965 131.690 105.135 ;
        RECT 131.945 105.055 132.305 105.635 ;
        RECT 129.135 104.565 129.395 104.895 ;
        RECT 129.605 104.395 129.880 104.875 ;
        RECT 130.090 104.565 130.295 104.965 ;
        RECT 130.465 104.395 130.800 104.795 ;
        RECT 130.980 104.395 131.315 104.795 ;
        RECT 131.485 104.565 131.690 104.965 ;
        RECT 132.475 104.895 132.645 105.805 ;
        RECT 133.275 105.780 133.565 106.945 ;
        RECT 133.825 106.325 133.995 106.755 ;
        RECT 134.165 106.495 134.495 106.945 ;
        RECT 133.825 106.095 134.500 106.325 ;
        RECT 131.900 104.395 132.175 104.875 ;
        RECT 132.385 104.565 132.645 104.895 ;
        RECT 133.275 104.395 133.565 105.120 ;
        RECT 133.795 105.075 134.095 105.925 ;
        RECT 134.265 105.445 134.500 106.095 ;
        RECT 134.670 105.785 134.955 106.730 ;
        RECT 135.135 106.475 135.820 106.945 ;
        RECT 135.130 105.955 135.825 106.265 ;
        RECT 136.000 105.890 136.305 106.675 ;
        RECT 134.670 105.635 135.530 105.785 ;
        RECT 136.095 105.755 136.305 105.890 ;
        RECT 134.670 105.615 135.955 105.635 ;
        RECT 134.265 105.115 134.800 105.445 ;
        RECT 134.970 105.255 135.955 105.615 ;
        RECT 134.265 104.965 134.485 105.115 ;
        RECT 133.740 104.395 134.075 104.900 ;
        RECT 134.245 104.590 134.485 104.965 ;
        RECT 134.970 104.920 135.140 105.255 ;
        RECT 136.130 105.085 136.305 105.755 ;
        RECT 134.765 104.725 135.140 104.920 ;
        RECT 134.765 104.580 134.935 104.725 ;
        RECT 135.500 104.395 135.895 104.890 ;
        RECT 136.065 104.565 136.305 105.085 ;
        RECT 136.495 106.095 136.755 106.775 ;
        RECT 136.925 106.165 137.175 106.945 ;
        RECT 137.425 106.395 137.675 106.775 ;
        RECT 137.845 106.565 138.200 106.945 ;
        RECT 139.205 106.555 139.540 106.775 ;
        RECT 138.805 106.395 139.035 106.435 ;
        RECT 137.425 106.195 139.035 106.395 ;
        RECT 137.425 106.185 138.260 106.195 ;
        RECT 138.850 106.105 139.035 106.195 ;
        RECT 136.495 104.905 136.665 106.095 ;
        RECT 138.365 105.995 138.695 106.025 ;
        RECT 136.895 105.935 138.695 105.995 ;
        RECT 139.285 105.935 139.540 106.555 ;
        RECT 136.835 105.825 139.540 105.935 ;
        RECT 139.715 105.855 141.385 106.945 ;
        RECT 136.835 105.790 137.035 105.825 ;
        RECT 136.835 105.215 137.005 105.790 ;
        RECT 138.365 105.765 139.540 105.825 ;
        RECT 137.235 105.350 137.645 105.655 ;
        RECT 137.815 105.385 138.145 105.595 ;
        RECT 136.835 105.095 137.105 105.215 ;
        RECT 136.835 105.050 137.680 105.095 ;
        RECT 136.925 104.925 137.680 105.050 ;
        RECT 137.935 104.985 138.145 105.385 ;
        RECT 138.390 105.385 138.865 105.595 ;
        RECT 139.055 105.385 139.545 105.585 ;
        RECT 138.390 104.985 138.610 105.385 ;
        RECT 139.715 105.165 140.465 105.685 ;
        RECT 140.635 105.335 141.385 105.855 ;
        RECT 142.105 106.015 142.275 106.775 ;
        RECT 142.490 106.185 142.820 106.945 ;
        RECT 142.105 105.845 142.820 106.015 ;
        RECT 142.990 105.870 143.245 106.775 ;
        RECT 142.015 105.295 142.370 105.665 ;
        RECT 142.650 105.635 142.820 105.845 ;
        RECT 142.650 105.305 142.905 105.635 ;
        RECT 136.495 104.895 136.725 104.905 ;
        RECT 136.495 104.565 136.755 104.895 ;
        RECT 137.510 104.775 137.680 104.925 ;
        RECT 136.925 104.395 137.255 104.755 ;
        RECT 137.510 104.565 138.810 104.775 ;
        RECT 139.085 104.395 139.540 105.160 ;
        RECT 139.715 104.395 141.385 105.165 ;
        RECT 142.650 105.115 142.820 105.305 ;
        RECT 143.075 105.140 143.245 105.870 ;
        RECT 143.420 105.795 143.680 106.945 ;
        RECT 143.945 106.015 144.115 106.775 ;
        RECT 144.330 106.185 144.660 106.945 ;
        RECT 143.945 105.845 144.660 106.015 ;
        RECT 144.830 105.870 145.085 106.775 ;
        RECT 143.855 105.295 144.210 105.665 ;
        RECT 144.490 105.635 144.660 105.845 ;
        RECT 144.490 105.305 144.745 105.635 ;
        RECT 142.105 104.945 142.820 105.115 ;
        RECT 142.105 104.565 142.275 104.945 ;
        RECT 142.490 104.395 142.820 104.775 ;
        RECT 142.990 104.565 143.245 105.140 ;
        RECT 143.420 104.395 143.680 105.235 ;
        RECT 144.490 105.115 144.660 105.305 ;
        RECT 144.915 105.140 145.085 105.870 ;
        RECT 145.260 105.795 145.520 106.945 ;
        RECT 145.695 105.855 146.905 106.945 ;
        RECT 145.695 105.315 146.215 105.855 ;
        RECT 143.945 104.945 144.660 105.115 ;
        RECT 143.945 104.565 144.115 104.945 ;
        RECT 144.330 104.395 144.660 104.775 ;
        RECT 144.830 104.565 145.085 105.140 ;
        RECT 145.260 104.395 145.520 105.235 ;
        RECT 146.385 105.145 146.905 105.685 ;
        RECT 145.695 104.395 146.905 105.145 ;
        RECT 17.270 104.225 146.990 104.395 ;
        RECT 17.355 103.475 18.565 104.225 ;
        RECT 17.355 102.935 17.875 103.475 ;
        RECT 18.740 103.385 19.000 104.225 ;
        RECT 19.175 103.480 19.430 104.055 ;
        RECT 19.600 103.845 19.930 104.225 ;
        RECT 20.145 103.675 20.315 104.055 ;
        RECT 19.600 103.505 20.315 103.675 ;
        RECT 18.045 102.765 18.565 103.305 ;
        RECT 17.355 101.675 18.565 102.765 ;
        RECT 18.740 101.675 19.000 102.825 ;
        RECT 19.175 102.750 19.345 103.480 ;
        RECT 19.600 103.315 19.770 103.505 ;
        RECT 20.580 103.385 20.840 104.225 ;
        RECT 21.015 103.480 21.270 104.055 ;
        RECT 21.440 103.845 21.770 104.225 ;
        RECT 21.985 103.675 22.155 104.055 ;
        RECT 21.440 103.505 22.155 103.675 ;
        RECT 19.515 102.985 19.770 103.315 ;
        RECT 19.600 102.775 19.770 102.985 ;
        RECT 20.050 102.955 20.405 103.325 ;
        RECT 19.175 101.845 19.430 102.750 ;
        RECT 19.600 102.605 20.315 102.775 ;
        RECT 19.600 101.675 19.930 102.435 ;
        RECT 20.145 101.845 20.315 102.605 ;
        RECT 20.580 101.675 20.840 102.825 ;
        RECT 21.015 102.750 21.185 103.480 ;
        RECT 21.440 103.315 21.610 103.505 ;
        RECT 22.690 103.415 22.935 104.020 ;
        RECT 23.155 103.690 23.665 104.225 ;
        RECT 21.355 102.985 21.610 103.315 ;
        RECT 21.440 102.775 21.610 102.985 ;
        RECT 21.890 102.955 22.245 103.325 ;
        RECT 22.415 103.245 23.645 103.415 ;
        RECT 21.015 101.845 21.270 102.750 ;
        RECT 21.440 102.605 22.155 102.775 ;
        RECT 21.440 101.675 21.770 102.435 ;
        RECT 21.985 101.845 22.155 102.605 ;
        RECT 22.415 102.435 22.755 103.245 ;
        RECT 22.925 102.680 23.675 102.870 ;
        RECT 22.415 102.025 22.930 102.435 ;
        RECT 23.165 101.675 23.335 102.435 ;
        RECT 23.505 102.015 23.675 102.680 ;
        RECT 23.845 102.695 24.035 104.055 ;
        RECT 24.205 103.545 24.480 104.055 ;
        RECT 24.670 103.690 25.200 104.055 ;
        RECT 25.625 103.825 25.955 104.225 ;
        RECT 25.025 103.655 25.200 103.690 ;
        RECT 24.205 103.375 24.485 103.545 ;
        RECT 24.205 102.895 24.480 103.375 ;
        RECT 24.685 102.695 24.855 103.495 ;
        RECT 23.845 102.525 24.855 102.695 ;
        RECT 25.025 103.485 25.955 103.655 ;
        RECT 26.125 103.485 26.380 104.055 ;
        RECT 25.025 102.355 25.195 103.485 ;
        RECT 25.785 103.315 25.955 103.485 ;
        RECT 24.070 102.185 25.195 102.355 ;
        RECT 25.365 102.985 25.560 103.315 ;
        RECT 25.785 102.985 26.040 103.315 ;
        RECT 25.365 102.015 25.535 102.985 ;
        RECT 26.210 102.815 26.380 103.485 ;
        RECT 23.505 101.845 25.535 102.015 ;
        RECT 25.705 101.675 25.875 102.815 ;
        RECT 26.045 101.845 26.380 102.815 ;
        RECT 26.560 103.485 26.815 104.055 ;
        RECT 26.985 103.825 27.315 104.225 ;
        RECT 27.740 103.690 28.270 104.055 ;
        RECT 27.740 103.655 27.915 103.690 ;
        RECT 26.985 103.485 27.915 103.655 ;
        RECT 26.560 102.815 26.730 103.485 ;
        RECT 26.985 103.315 27.155 103.485 ;
        RECT 26.900 102.985 27.155 103.315 ;
        RECT 27.380 102.985 27.575 103.315 ;
        RECT 26.560 101.845 26.895 102.815 ;
        RECT 27.065 101.675 27.235 102.815 ;
        RECT 27.405 102.015 27.575 102.985 ;
        RECT 27.745 102.355 27.915 103.485 ;
        RECT 28.085 102.695 28.255 103.495 ;
        RECT 28.460 103.205 28.735 104.055 ;
        RECT 28.455 103.035 28.735 103.205 ;
        RECT 28.460 102.895 28.735 103.035 ;
        RECT 28.905 102.695 29.095 104.055 ;
        RECT 29.275 103.690 29.785 104.225 ;
        RECT 30.005 103.415 30.250 104.020 ;
        RECT 31.175 103.415 31.415 104.225 ;
        RECT 31.585 103.415 31.915 104.055 ;
        RECT 32.085 103.415 32.355 104.225 ;
        RECT 32.535 103.550 32.810 103.895 ;
        RECT 33.000 103.825 33.380 104.225 ;
        RECT 33.550 103.655 33.720 104.005 ;
        RECT 33.890 103.825 34.220 104.225 ;
        RECT 34.395 103.655 34.565 104.005 ;
        RECT 34.765 103.725 35.095 104.225 ;
        RECT 29.295 103.245 30.525 103.415 ;
        RECT 28.085 102.525 29.095 102.695 ;
        RECT 29.265 102.680 30.015 102.870 ;
        RECT 27.745 102.185 28.870 102.355 ;
        RECT 29.265 102.015 29.435 102.680 ;
        RECT 30.185 102.435 30.525 103.245 ;
        RECT 31.155 102.985 31.505 103.235 ;
        RECT 31.675 102.815 31.845 103.415 ;
        RECT 32.015 102.985 32.365 103.235 ;
        RECT 32.535 102.815 32.705 103.550 ;
        RECT 32.980 103.485 34.565 103.655 ;
        RECT 32.980 103.315 33.150 103.485 ;
        RECT 35.290 103.315 35.535 104.005 ;
        RECT 35.705 103.725 36.045 104.225 ;
        RECT 32.875 102.985 33.150 103.315 ;
        RECT 33.320 102.985 33.700 103.315 ;
        RECT 32.980 102.815 33.150 102.985 ;
        RECT 27.405 101.845 29.435 102.015 ;
        RECT 29.605 101.675 29.775 102.435 ;
        RECT 30.010 102.025 30.525 102.435 ;
        RECT 31.165 102.645 31.845 102.815 ;
        RECT 31.165 101.860 31.495 102.645 ;
        RECT 32.025 101.675 32.355 102.815 ;
        RECT 32.535 101.845 32.810 102.815 ;
        RECT 32.980 102.645 33.640 102.815 ;
        RECT 33.870 102.695 34.610 103.315 ;
        RECT 34.880 102.985 35.535 103.315 ;
        RECT 35.705 102.985 36.045 103.555 ;
        RECT 36.675 103.485 37.115 104.045 ;
        RECT 37.285 103.485 37.735 104.225 ;
        RECT 37.905 103.655 38.075 104.055 ;
        RECT 38.245 103.825 38.665 104.225 ;
        RECT 38.835 103.655 39.065 104.055 ;
        RECT 37.905 103.485 39.065 103.655 ;
        RECT 39.235 103.485 39.725 104.055 ;
        RECT 33.470 102.525 33.640 102.645 ;
        RECT 34.780 102.525 35.100 102.815 ;
        RECT 33.020 101.675 33.300 102.475 ;
        RECT 33.470 102.355 35.100 102.525 ;
        RECT 35.295 102.390 35.535 102.985 ;
        RECT 33.470 101.895 35.520 102.185 ;
        RECT 35.705 101.675 36.045 102.750 ;
        RECT 36.675 102.475 36.985 103.485 ;
        RECT 37.155 102.865 37.325 103.315 ;
        RECT 37.495 103.035 37.885 103.315 ;
        RECT 38.070 102.985 38.315 103.315 ;
        RECT 37.155 102.695 37.945 102.865 ;
        RECT 36.675 101.845 37.115 102.475 ;
        RECT 37.290 101.675 37.605 102.525 ;
        RECT 37.775 102.015 37.945 102.695 ;
        RECT 38.115 102.185 38.315 102.985 ;
        RECT 38.515 102.185 38.765 103.315 ;
        RECT 38.980 102.985 39.385 103.315 ;
        RECT 39.555 102.815 39.725 103.485 ;
        RECT 40.365 103.415 40.635 104.225 ;
        RECT 40.805 103.415 41.135 104.055 ;
        RECT 41.305 103.415 41.545 104.225 ;
        RECT 41.735 103.475 42.945 104.225 ;
        RECT 43.115 103.500 43.405 104.225 ;
        RECT 43.575 103.680 48.920 104.225 ;
        RECT 49.095 103.680 54.440 104.225 ;
        RECT 40.355 102.985 40.705 103.235 ;
        RECT 40.875 102.815 41.045 103.415 ;
        RECT 41.215 102.985 41.565 103.235 ;
        RECT 41.735 102.935 42.255 103.475 ;
        RECT 38.955 102.645 39.725 102.815 ;
        RECT 38.955 102.015 39.205 102.645 ;
        RECT 37.775 101.845 39.205 102.015 ;
        RECT 39.385 101.675 39.715 102.475 ;
        RECT 40.365 101.675 40.695 102.815 ;
        RECT 40.875 102.645 41.555 102.815 ;
        RECT 42.425 102.765 42.945 103.305 ;
        RECT 45.160 102.850 45.500 103.680 ;
        RECT 41.225 101.860 41.555 102.645 ;
        RECT 41.735 101.675 42.945 102.765 ;
        RECT 43.115 101.675 43.405 102.840 ;
        RECT 46.980 102.110 47.330 103.360 ;
        RECT 50.680 102.850 51.020 103.680 ;
        RECT 54.615 103.455 58.125 104.225 ;
        RECT 58.775 103.535 59.015 104.055 ;
        RECT 59.185 103.730 59.580 104.225 ;
        RECT 60.145 103.895 60.315 104.040 ;
        RECT 59.940 103.700 60.315 103.895 ;
        RECT 52.500 102.110 52.850 103.360 ;
        RECT 54.615 102.935 56.265 103.455 ;
        RECT 56.435 102.765 58.125 103.285 ;
        RECT 43.575 101.675 48.920 102.110 ;
        RECT 49.095 101.675 54.440 102.110 ;
        RECT 54.615 101.675 58.125 102.765 ;
        RECT 58.775 102.730 58.950 103.535 ;
        RECT 59.940 103.365 60.110 103.700 ;
        RECT 60.595 103.655 60.835 104.030 ;
        RECT 61.005 103.720 61.340 104.225 ;
        RECT 61.605 103.675 61.775 103.965 ;
        RECT 61.945 103.845 62.275 104.225 ;
        RECT 60.595 103.505 60.815 103.655 ;
        RECT 59.125 103.005 60.110 103.365 ;
        RECT 60.280 103.175 60.815 103.505 ;
        RECT 59.125 102.985 60.410 103.005 ;
        RECT 59.550 102.835 60.410 102.985 ;
        RECT 58.775 101.945 59.080 102.730 ;
        RECT 59.255 102.355 59.950 102.665 ;
        RECT 59.260 101.675 59.945 102.145 ;
        RECT 60.125 101.890 60.410 102.835 ;
        RECT 60.580 102.525 60.815 103.175 ;
        RECT 60.985 102.695 61.285 103.545 ;
        RECT 61.605 103.505 62.270 103.675 ;
        RECT 61.520 102.685 61.870 103.335 ;
        RECT 60.580 102.295 61.255 102.525 ;
        RECT 62.040 102.515 62.270 103.505 ;
        RECT 60.585 101.675 60.915 102.125 ;
        RECT 61.085 101.865 61.255 102.295 ;
        RECT 61.605 102.345 62.270 102.515 ;
        RECT 61.605 101.845 61.775 102.345 ;
        RECT 61.945 101.675 62.275 102.175 ;
        RECT 62.445 101.845 62.630 103.965 ;
        RECT 62.885 103.765 63.135 104.225 ;
        RECT 63.305 103.775 63.640 103.945 ;
        RECT 63.835 103.775 64.510 103.945 ;
        RECT 63.305 103.635 63.475 103.775 ;
        RECT 62.800 102.645 63.080 103.595 ;
        RECT 63.250 103.505 63.475 103.635 ;
        RECT 63.250 102.400 63.420 103.505 ;
        RECT 63.645 103.355 64.170 103.575 ;
        RECT 63.590 102.590 63.830 103.185 ;
        RECT 64.000 102.655 64.170 103.355 ;
        RECT 64.340 102.995 64.510 103.775 ;
        RECT 64.830 103.725 65.200 104.225 ;
        RECT 65.380 103.775 65.785 103.945 ;
        RECT 65.955 103.775 66.740 103.945 ;
        RECT 65.380 103.545 65.550 103.775 ;
        RECT 64.720 103.245 65.550 103.545 ;
        RECT 65.935 103.275 66.400 103.605 ;
        RECT 64.720 103.215 64.920 103.245 ;
        RECT 65.040 102.995 65.210 103.065 ;
        RECT 64.340 102.825 65.210 102.995 ;
        RECT 64.700 102.735 65.210 102.825 ;
        RECT 63.250 102.270 63.555 102.400 ;
        RECT 64.000 102.290 64.530 102.655 ;
        RECT 62.870 101.675 63.135 102.135 ;
        RECT 63.305 101.845 63.555 102.270 ;
        RECT 64.700 102.120 64.870 102.735 ;
        RECT 63.765 101.950 64.870 102.120 ;
        RECT 65.040 101.675 65.210 102.475 ;
        RECT 65.380 102.175 65.550 103.245 ;
        RECT 65.720 102.345 65.910 103.065 ;
        RECT 66.080 102.315 66.400 103.275 ;
        RECT 66.570 103.315 66.740 103.775 ;
        RECT 67.015 103.695 67.225 104.225 ;
        RECT 67.485 103.485 67.815 104.010 ;
        RECT 67.985 103.615 68.155 104.225 ;
        RECT 68.325 103.570 68.655 104.005 ;
        RECT 68.325 103.485 68.705 103.570 ;
        RECT 68.875 103.500 69.165 104.225 ;
        RECT 67.615 103.315 67.815 103.485 ;
        RECT 68.480 103.445 68.705 103.485 ;
        RECT 66.570 102.985 67.445 103.315 ;
        RECT 67.615 102.985 68.365 103.315 ;
        RECT 65.380 101.845 65.630 102.175 ;
        RECT 66.570 102.145 66.740 102.985 ;
        RECT 67.615 102.780 67.805 102.985 ;
        RECT 68.535 102.865 68.705 103.445 ;
        RECT 68.490 102.815 68.705 102.865 ;
        RECT 69.340 103.485 69.595 104.055 ;
        RECT 69.765 103.825 70.095 104.225 ;
        RECT 70.520 103.690 71.050 104.055 ;
        RECT 71.240 103.885 71.515 104.055 ;
        RECT 71.235 103.715 71.515 103.885 ;
        RECT 70.520 103.655 70.695 103.690 ;
        RECT 69.765 103.485 70.695 103.655 ;
        RECT 66.910 102.405 67.805 102.780 ;
        RECT 68.315 102.735 68.705 102.815 ;
        RECT 65.855 101.975 66.740 102.145 ;
        RECT 66.920 101.675 67.235 102.175 ;
        RECT 67.465 101.845 67.805 102.405 ;
        RECT 67.975 101.675 68.145 102.685 ;
        RECT 68.315 101.890 68.645 102.735 ;
        RECT 68.875 101.675 69.165 102.840 ;
        RECT 69.340 102.815 69.510 103.485 ;
        RECT 69.765 103.315 69.935 103.485 ;
        RECT 69.680 102.985 69.935 103.315 ;
        RECT 70.160 102.985 70.355 103.315 ;
        RECT 69.340 101.845 69.675 102.815 ;
        RECT 69.845 101.675 70.015 102.815 ;
        RECT 70.185 102.015 70.355 102.985 ;
        RECT 70.525 102.355 70.695 103.485 ;
        RECT 70.865 102.695 71.035 103.495 ;
        RECT 71.240 102.895 71.515 103.715 ;
        RECT 71.685 102.695 71.875 104.055 ;
        RECT 72.055 103.690 72.565 104.225 ;
        RECT 72.785 103.415 73.030 104.020 ;
        RECT 73.480 103.720 73.815 104.225 ;
        RECT 73.985 103.655 74.225 104.030 ;
        RECT 74.505 103.895 74.675 104.040 ;
        RECT 74.505 103.700 74.880 103.895 ;
        RECT 75.240 103.730 75.635 104.225 ;
        RECT 72.075 103.245 73.305 103.415 ;
        RECT 70.865 102.525 71.875 102.695 ;
        RECT 72.045 102.680 72.795 102.870 ;
        RECT 70.525 102.185 71.650 102.355 ;
        RECT 72.045 102.015 72.215 102.680 ;
        RECT 72.965 102.435 73.305 103.245 ;
        RECT 73.535 102.695 73.835 103.545 ;
        RECT 74.005 103.505 74.225 103.655 ;
        RECT 74.005 103.175 74.540 103.505 ;
        RECT 74.710 103.365 74.880 103.700 ;
        RECT 75.805 103.535 76.045 104.055 ;
        RECT 74.005 102.525 74.240 103.175 ;
        RECT 74.710 103.005 75.695 103.365 ;
        RECT 70.185 101.845 72.215 102.015 ;
        RECT 72.385 101.675 72.555 102.435 ;
        RECT 72.790 102.025 73.305 102.435 ;
        RECT 73.565 102.295 74.240 102.525 ;
        RECT 74.410 102.985 75.695 103.005 ;
        RECT 74.410 102.835 75.270 102.985 ;
        RECT 73.565 101.865 73.735 102.295 ;
        RECT 73.905 101.675 74.235 102.125 ;
        RECT 74.410 101.890 74.695 102.835 ;
        RECT 75.870 102.730 76.045 103.535 ;
        RECT 74.870 102.355 75.565 102.665 ;
        RECT 74.875 101.675 75.560 102.145 ;
        RECT 75.740 101.945 76.045 102.730 ;
        RECT 76.240 103.485 76.495 104.055 ;
        RECT 76.665 103.825 76.995 104.225 ;
        RECT 77.420 103.690 77.950 104.055 ;
        RECT 77.420 103.655 77.595 103.690 ;
        RECT 76.665 103.485 77.595 103.655 ;
        RECT 76.240 102.815 76.410 103.485 ;
        RECT 76.665 103.315 76.835 103.485 ;
        RECT 76.580 102.985 76.835 103.315 ;
        RECT 77.060 102.985 77.255 103.315 ;
        RECT 76.240 101.845 76.575 102.815 ;
        RECT 76.745 101.675 76.915 102.815 ;
        RECT 77.085 102.015 77.255 102.985 ;
        RECT 77.425 102.355 77.595 103.485 ;
        RECT 77.765 102.695 77.935 103.495 ;
        RECT 78.140 103.205 78.415 104.055 ;
        RECT 78.135 103.035 78.415 103.205 ;
        RECT 78.140 102.895 78.415 103.035 ;
        RECT 78.585 102.695 78.775 104.055 ;
        RECT 78.955 103.690 79.465 104.225 ;
        RECT 79.685 103.415 79.930 104.020 ;
        RECT 80.465 103.675 80.635 103.965 ;
        RECT 80.805 103.845 81.135 104.225 ;
        RECT 80.465 103.505 81.130 103.675 ;
        RECT 78.975 103.245 80.205 103.415 ;
        RECT 77.765 102.525 78.775 102.695 ;
        RECT 78.945 102.680 79.695 102.870 ;
        RECT 77.425 102.185 78.550 102.355 ;
        RECT 78.945 102.015 79.115 102.680 ;
        RECT 79.865 102.435 80.205 103.245 ;
        RECT 80.380 102.685 80.730 103.335 ;
        RECT 80.900 102.515 81.130 103.505 ;
        RECT 77.085 101.845 79.115 102.015 ;
        RECT 79.285 101.675 79.455 102.435 ;
        RECT 79.690 102.025 80.205 102.435 ;
        RECT 80.465 102.345 81.130 102.515 ;
        RECT 80.465 101.845 80.635 102.345 ;
        RECT 80.805 101.675 81.135 102.175 ;
        RECT 81.305 101.845 81.490 103.965 ;
        RECT 81.745 103.765 81.995 104.225 ;
        RECT 82.165 103.775 82.500 103.945 ;
        RECT 82.695 103.775 83.370 103.945 ;
        RECT 82.165 103.635 82.335 103.775 ;
        RECT 81.660 102.645 81.940 103.595 ;
        RECT 82.110 103.505 82.335 103.635 ;
        RECT 82.110 102.400 82.280 103.505 ;
        RECT 82.505 103.355 83.030 103.575 ;
        RECT 82.450 102.590 82.690 103.185 ;
        RECT 82.860 102.655 83.030 103.355 ;
        RECT 83.200 102.995 83.370 103.775 ;
        RECT 83.690 103.725 84.060 104.225 ;
        RECT 84.240 103.775 84.645 103.945 ;
        RECT 84.815 103.775 85.600 103.945 ;
        RECT 84.240 103.545 84.410 103.775 ;
        RECT 83.580 103.245 84.410 103.545 ;
        RECT 84.795 103.275 85.260 103.605 ;
        RECT 83.580 103.215 83.780 103.245 ;
        RECT 83.900 102.995 84.070 103.065 ;
        RECT 83.200 102.825 84.070 102.995 ;
        RECT 83.560 102.735 84.070 102.825 ;
        RECT 82.110 102.270 82.415 102.400 ;
        RECT 82.860 102.290 83.390 102.655 ;
        RECT 81.730 101.675 81.995 102.135 ;
        RECT 82.165 101.845 82.415 102.270 ;
        RECT 83.560 102.120 83.730 102.735 ;
        RECT 82.625 101.950 83.730 102.120 ;
        RECT 83.900 101.675 84.070 102.475 ;
        RECT 84.240 102.175 84.410 103.245 ;
        RECT 84.580 102.345 84.770 103.065 ;
        RECT 84.940 102.315 85.260 103.275 ;
        RECT 85.430 103.315 85.600 103.775 ;
        RECT 85.875 103.695 86.085 104.225 ;
        RECT 86.345 103.485 86.675 104.010 ;
        RECT 86.845 103.615 87.015 104.225 ;
        RECT 87.185 103.570 87.515 104.005 ;
        RECT 87.185 103.485 87.565 103.570 ;
        RECT 86.475 103.315 86.675 103.485 ;
        RECT 87.340 103.445 87.565 103.485 ;
        RECT 85.430 102.985 86.305 103.315 ;
        RECT 86.475 102.985 87.225 103.315 ;
        RECT 84.240 101.845 84.490 102.175 ;
        RECT 85.430 102.145 85.600 102.985 ;
        RECT 86.475 102.780 86.665 102.985 ;
        RECT 87.395 102.865 87.565 103.445 ;
        RECT 87.350 102.815 87.565 102.865 ;
        RECT 85.770 102.405 86.665 102.780 ;
        RECT 87.175 102.735 87.565 102.815 ;
        RECT 87.740 103.485 87.995 104.055 ;
        RECT 88.165 103.825 88.495 104.225 ;
        RECT 88.920 103.690 89.450 104.055 ;
        RECT 89.640 103.885 89.915 104.055 ;
        RECT 89.635 103.715 89.915 103.885 ;
        RECT 88.920 103.655 89.095 103.690 ;
        RECT 88.165 103.485 89.095 103.655 ;
        RECT 87.740 102.815 87.910 103.485 ;
        RECT 88.165 103.315 88.335 103.485 ;
        RECT 88.080 102.985 88.335 103.315 ;
        RECT 88.560 102.985 88.755 103.315 ;
        RECT 84.715 101.975 85.600 102.145 ;
        RECT 85.780 101.675 86.095 102.175 ;
        RECT 86.325 101.845 86.665 102.405 ;
        RECT 86.835 101.675 87.005 102.685 ;
        RECT 87.175 101.890 87.505 102.735 ;
        RECT 87.740 101.845 88.075 102.815 ;
        RECT 88.245 101.675 88.415 102.815 ;
        RECT 88.585 102.015 88.755 102.985 ;
        RECT 88.925 102.355 89.095 103.485 ;
        RECT 89.265 102.695 89.435 103.495 ;
        RECT 89.640 102.895 89.915 103.715 ;
        RECT 90.085 102.695 90.275 104.055 ;
        RECT 90.455 103.690 90.965 104.225 ;
        RECT 91.185 103.415 91.430 104.020 ;
        RECT 91.880 103.720 92.215 104.225 ;
        RECT 92.385 103.655 92.625 104.030 ;
        RECT 92.905 103.895 93.075 104.040 ;
        RECT 92.905 103.700 93.280 103.895 ;
        RECT 93.640 103.730 94.035 104.225 ;
        RECT 90.475 103.245 91.705 103.415 ;
        RECT 89.265 102.525 90.275 102.695 ;
        RECT 90.445 102.680 91.195 102.870 ;
        RECT 88.925 102.185 90.050 102.355 ;
        RECT 90.445 102.015 90.615 102.680 ;
        RECT 91.365 102.435 91.705 103.245 ;
        RECT 91.935 102.695 92.235 103.545 ;
        RECT 92.405 103.505 92.625 103.655 ;
        RECT 92.405 103.175 92.940 103.505 ;
        RECT 93.110 103.365 93.280 103.700 ;
        RECT 94.205 103.535 94.445 104.055 ;
        RECT 92.405 102.525 92.640 103.175 ;
        RECT 93.110 103.005 94.095 103.365 ;
        RECT 88.585 101.845 90.615 102.015 ;
        RECT 90.785 101.675 90.955 102.435 ;
        RECT 91.190 102.025 91.705 102.435 ;
        RECT 91.965 102.295 92.640 102.525 ;
        RECT 92.810 102.985 94.095 103.005 ;
        RECT 92.810 102.835 93.670 102.985 ;
        RECT 94.270 102.865 94.445 103.535 ;
        RECT 94.635 103.500 94.925 104.225 ;
        RECT 95.185 103.675 95.355 103.965 ;
        RECT 95.525 103.845 95.855 104.225 ;
        RECT 95.185 103.505 95.850 103.675 ;
        RECT 91.965 101.865 92.135 102.295 ;
        RECT 92.305 101.675 92.635 102.125 ;
        RECT 92.810 101.890 93.095 102.835 ;
        RECT 94.235 102.730 94.445 102.865 ;
        RECT 93.270 102.355 93.965 102.665 ;
        RECT 93.275 101.675 93.960 102.145 ;
        RECT 94.140 101.945 94.445 102.730 ;
        RECT 94.635 101.675 94.925 102.840 ;
        RECT 95.100 102.685 95.450 103.335 ;
        RECT 95.620 102.515 95.850 103.505 ;
        RECT 95.185 102.345 95.850 102.515 ;
        RECT 95.185 101.845 95.355 102.345 ;
        RECT 95.525 101.675 95.855 102.175 ;
        RECT 96.025 101.845 96.210 103.965 ;
        RECT 96.465 103.765 96.715 104.225 ;
        RECT 96.885 103.775 97.220 103.945 ;
        RECT 97.415 103.775 98.090 103.945 ;
        RECT 96.885 103.635 97.055 103.775 ;
        RECT 96.380 102.645 96.660 103.595 ;
        RECT 96.830 103.505 97.055 103.635 ;
        RECT 96.830 102.400 97.000 103.505 ;
        RECT 97.225 103.355 97.750 103.575 ;
        RECT 97.170 102.590 97.410 103.185 ;
        RECT 97.580 102.655 97.750 103.355 ;
        RECT 97.920 102.995 98.090 103.775 ;
        RECT 98.410 103.725 98.780 104.225 ;
        RECT 98.960 103.775 99.365 103.945 ;
        RECT 99.535 103.775 100.320 103.945 ;
        RECT 98.960 103.545 99.130 103.775 ;
        RECT 98.300 103.245 99.130 103.545 ;
        RECT 99.515 103.275 99.980 103.605 ;
        RECT 98.300 103.215 98.500 103.245 ;
        RECT 98.620 102.995 98.790 103.065 ;
        RECT 97.920 102.825 98.790 102.995 ;
        RECT 98.280 102.735 98.790 102.825 ;
        RECT 96.830 102.270 97.135 102.400 ;
        RECT 97.580 102.290 98.110 102.655 ;
        RECT 96.450 101.675 96.715 102.135 ;
        RECT 96.885 101.845 97.135 102.270 ;
        RECT 98.280 102.120 98.450 102.735 ;
        RECT 97.345 101.950 98.450 102.120 ;
        RECT 98.620 101.675 98.790 102.475 ;
        RECT 98.960 102.175 99.130 103.245 ;
        RECT 99.300 102.345 99.490 103.065 ;
        RECT 99.660 102.315 99.980 103.275 ;
        RECT 100.150 103.315 100.320 103.775 ;
        RECT 100.595 103.695 100.805 104.225 ;
        RECT 101.065 103.485 101.395 104.010 ;
        RECT 101.565 103.615 101.735 104.225 ;
        RECT 101.905 103.570 102.235 104.005 ;
        RECT 101.905 103.485 102.285 103.570 ;
        RECT 101.195 103.315 101.395 103.485 ;
        RECT 102.060 103.445 102.285 103.485 ;
        RECT 100.150 102.985 101.025 103.315 ;
        RECT 101.195 102.985 101.945 103.315 ;
        RECT 98.960 101.845 99.210 102.175 ;
        RECT 100.150 102.145 100.320 102.985 ;
        RECT 101.195 102.780 101.385 102.985 ;
        RECT 102.115 102.865 102.285 103.445 ;
        RECT 102.070 102.815 102.285 102.865 ;
        RECT 100.490 102.405 101.385 102.780 ;
        RECT 101.895 102.735 102.285 102.815 ;
        RECT 102.460 103.485 102.715 104.055 ;
        RECT 102.885 103.825 103.215 104.225 ;
        RECT 103.640 103.690 104.170 104.055 ;
        RECT 104.360 103.885 104.635 104.055 ;
        RECT 104.355 103.715 104.635 103.885 ;
        RECT 103.640 103.655 103.815 103.690 ;
        RECT 102.885 103.485 103.815 103.655 ;
        RECT 102.460 102.815 102.630 103.485 ;
        RECT 102.885 103.315 103.055 103.485 ;
        RECT 102.800 102.985 103.055 103.315 ;
        RECT 103.280 102.985 103.475 103.315 ;
        RECT 99.435 101.975 100.320 102.145 ;
        RECT 100.500 101.675 100.815 102.175 ;
        RECT 101.045 101.845 101.385 102.405 ;
        RECT 101.555 101.675 101.725 102.685 ;
        RECT 101.895 101.890 102.225 102.735 ;
        RECT 102.460 101.845 102.795 102.815 ;
        RECT 102.965 101.675 103.135 102.815 ;
        RECT 103.305 102.015 103.475 102.985 ;
        RECT 103.645 102.355 103.815 103.485 ;
        RECT 103.985 102.695 104.155 103.495 ;
        RECT 104.360 102.895 104.635 103.715 ;
        RECT 104.805 102.695 104.995 104.055 ;
        RECT 105.175 103.690 105.685 104.225 ;
        RECT 105.905 103.415 106.150 104.020 ;
        RECT 107.145 103.675 107.315 103.965 ;
        RECT 107.485 103.845 107.815 104.225 ;
        RECT 107.145 103.505 107.810 103.675 ;
        RECT 105.195 103.245 106.425 103.415 ;
        RECT 103.985 102.525 104.995 102.695 ;
        RECT 105.165 102.680 105.915 102.870 ;
        RECT 103.645 102.185 104.770 102.355 ;
        RECT 105.165 102.015 105.335 102.680 ;
        RECT 106.085 102.435 106.425 103.245 ;
        RECT 107.060 102.685 107.410 103.335 ;
        RECT 107.580 102.515 107.810 103.505 ;
        RECT 103.305 101.845 105.335 102.015 ;
        RECT 105.505 101.675 105.675 102.435 ;
        RECT 105.910 102.025 106.425 102.435 ;
        RECT 107.145 102.345 107.810 102.515 ;
        RECT 107.145 101.845 107.315 102.345 ;
        RECT 107.485 101.675 107.815 102.175 ;
        RECT 107.985 101.845 108.170 103.965 ;
        RECT 108.425 103.765 108.675 104.225 ;
        RECT 108.845 103.775 109.180 103.945 ;
        RECT 109.375 103.775 110.050 103.945 ;
        RECT 108.845 103.635 109.015 103.775 ;
        RECT 108.340 102.645 108.620 103.595 ;
        RECT 108.790 103.505 109.015 103.635 ;
        RECT 108.790 102.400 108.960 103.505 ;
        RECT 109.185 103.355 109.710 103.575 ;
        RECT 109.130 102.590 109.370 103.185 ;
        RECT 109.540 102.655 109.710 103.355 ;
        RECT 109.880 102.995 110.050 103.775 ;
        RECT 110.370 103.725 110.740 104.225 ;
        RECT 110.920 103.775 111.325 103.945 ;
        RECT 111.495 103.775 112.280 103.945 ;
        RECT 110.920 103.545 111.090 103.775 ;
        RECT 110.260 103.245 111.090 103.545 ;
        RECT 111.475 103.275 111.940 103.605 ;
        RECT 110.260 103.215 110.460 103.245 ;
        RECT 110.580 102.995 110.750 103.065 ;
        RECT 109.880 102.825 110.750 102.995 ;
        RECT 110.240 102.735 110.750 102.825 ;
        RECT 108.790 102.270 109.095 102.400 ;
        RECT 109.540 102.290 110.070 102.655 ;
        RECT 108.410 101.675 108.675 102.135 ;
        RECT 108.845 101.845 109.095 102.270 ;
        RECT 110.240 102.120 110.410 102.735 ;
        RECT 109.305 101.950 110.410 102.120 ;
        RECT 110.580 101.675 110.750 102.475 ;
        RECT 110.920 102.175 111.090 103.245 ;
        RECT 111.260 102.345 111.450 103.065 ;
        RECT 111.620 102.315 111.940 103.275 ;
        RECT 112.110 103.315 112.280 103.775 ;
        RECT 112.555 103.695 112.765 104.225 ;
        RECT 113.025 103.485 113.355 104.010 ;
        RECT 113.525 103.615 113.695 104.225 ;
        RECT 113.865 103.570 114.195 104.005 ;
        RECT 113.865 103.485 114.245 103.570 ;
        RECT 113.155 103.315 113.355 103.485 ;
        RECT 114.020 103.445 114.245 103.485 ;
        RECT 112.110 102.985 112.985 103.315 ;
        RECT 113.155 102.985 113.905 103.315 ;
        RECT 110.920 101.845 111.170 102.175 ;
        RECT 112.110 102.145 112.280 102.985 ;
        RECT 113.155 102.780 113.345 102.985 ;
        RECT 114.075 102.865 114.245 103.445 ;
        RECT 114.030 102.815 114.245 102.865 ;
        RECT 112.450 102.405 113.345 102.780 ;
        RECT 113.855 102.735 114.245 102.815 ;
        RECT 114.420 103.485 114.675 104.055 ;
        RECT 114.845 103.825 115.175 104.225 ;
        RECT 115.600 103.690 116.130 104.055 ;
        RECT 115.600 103.655 115.775 103.690 ;
        RECT 114.845 103.485 115.775 103.655 ;
        RECT 116.320 103.545 116.595 104.055 ;
        RECT 114.420 102.815 114.590 103.485 ;
        RECT 114.845 103.315 115.015 103.485 ;
        RECT 114.760 102.985 115.015 103.315 ;
        RECT 115.240 102.985 115.435 103.315 ;
        RECT 111.395 101.975 112.280 102.145 ;
        RECT 112.460 101.675 112.775 102.175 ;
        RECT 113.005 101.845 113.345 102.405 ;
        RECT 113.515 101.675 113.685 102.685 ;
        RECT 113.855 101.890 114.185 102.735 ;
        RECT 114.420 101.845 114.755 102.815 ;
        RECT 114.925 101.675 115.095 102.815 ;
        RECT 115.265 102.015 115.435 102.985 ;
        RECT 115.605 102.355 115.775 103.485 ;
        RECT 115.945 102.695 116.115 103.495 ;
        RECT 116.315 103.375 116.595 103.545 ;
        RECT 116.320 102.895 116.595 103.375 ;
        RECT 116.765 102.695 116.955 104.055 ;
        RECT 117.135 103.690 117.645 104.225 ;
        RECT 117.865 103.415 118.110 104.020 ;
        RECT 118.555 103.455 120.225 104.225 ;
        RECT 120.395 103.500 120.685 104.225 ;
        RECT 120.860 103.485 121.115 104.055 ;
        RECT 121.285 103.825 121.615 104.225 ;
        RECT 122.040 103.690 122.570 104.055 ;
        RECT 122.760 103.885 123.035 104.055 ;
        RECT 122.755 103.715 123.035 103.885 ;
        RECT 122.040 103.655 122.215 103.690 ;
        RECT 121.285 103.485 122.215 103.655 ;
        RECT 117.155 103.245 118.385 103.415 ;
        RECT 115.945 102.525 116.955 102.695 ;
        RECT 117.125 102.680 117.875 102.870 ;
        RECT 115.605 102.185 116.730 102.355 ;
        RECT 117.125 102.015 117.295 102.680 ;
        RECT 118.045 102.435 118.385 103.245 ;
        RECT 118.555 102.935 119.305 103.455 ;
        RECT 119.475 102.765 120.225 103.285 ;
        RECT 115.265 101.845 117.295 102.015 ;
        RECT 117.465 101.675 117.635 102.435 ;
        RECT 117.870 102.025 118.385 102.435 ;
        RECT 118.555 101.675 120.225 102.765 ;
        RECT 120.395 101.675 120.685 102.840 ;
        RECT 120.860 102.815 121.030 103.485 ;
        RECT 121.285 103.315 121.455 103.485 ;
        RECT 121.200 102.985 121.455 103.315 ;
        RECT 121.680 102.985 121.875 103.315 ;
        RECT 120.860 101.845 121.195 102.815 ;
        RECT 121.365 101.675 121.535 102.815 ;
        RECT 121.705 102.015 121.875 102.985 ;
        RECT 122.045 102.355 122.215 103.485 ;
        RECT 122.385 102.695 122.555 103.495 ;
        RECT 122.760 102.895 123.035 103.715 ;
        RECT 123.205 102.695 123.395 104.055 ;
        RECT 123.575 103.690 124.085 104.225 ;
        RECT 124.305 103.415 124.550 104.020 ;
        RECT 124.995 103.475 126.205 104.225 ;
        RECT 126.465 103.675 126.635 103.965 ;
        RECT 126.805 103.845 127.135 104.225 ;
        RECT 126.465 103.505 127.130 103.675 ;
        RECT 123.595 103.245 124.825 103.415 ;
        RECT 122.385 102.525 123.395 102.695 ;
        RECT 123.565 102.680 124.315 102.870 ;
        RECT 122.045 102.185 123.170 102.355 ;
        RECT 123.565 102.015 123.735 102.680 ;
        RECT 124.485 102.435 124.825 103.245 ;
        RECT 124.995 102.935 125.515 103.475 ;
        RECT 125.685 102.765 126.205 103.305 ;
        RECT 121.705 101.845 123.735 102.015 ;
        RECT 123.905 101.675 124.075 102.435 ;
        RECT 124.310 102.025 124.825 102.435 ;
        RECT 124.995 101.675 126.205 102.765 ;
        RECT 126.380 102.685 126.730 103.335 ;
        RECT 126.900 102.515 127.130 103.505 ;
        RECT 126.465 102.345 127.130 102.515 ;
        RECT 126.465 101.845 126.635 102.345 ;
        RECT 126.805 101.675 127.135 102.175 ;
        RECT 127.305 101.845 127.490 103.965 ;
        RECT 127.745 103.765 127.995 104.225 ;
        RECT 128.165 103.775 128.500 103.945 ;
        RECT 128.695 103.775 129.370 103.945 ;
        RECT 128.165 103.635 128.335 103.775 ;
        RECT 127.660 102.645 127.940 103.595 ;
        RECT 128.110 103.505 128.335 103.635 ;
        RECT 128.110 102.400 128.280 103.505 ;
        RECT 128.505 103.355 129.030 103.575 ;
        RECT 128.450 102.590 128.690 103.185 ;
        RECT 128.860 102.655 129.030 103.355 ;
        RECT 129.200 102.995 129.370 103.775 ;
        RECT 129.690 103.725 130.060 104.225 ;
        RECT 130.240 103.775 130.645 103.945 ;
        RECT 130.815 103.775 131.600 103.945 ;
        RECT 130.240 103.545 130.410 103.775 ;
        RECT 129.580 103.245 130.410 103.545 ;
        RECT 130.795 103.275 131.260 103.605 ;
        RECT 129.580 103.215 129.780 103.245 ;
        RECT 129.900 102.995 130.070 103.065 ;
        RECT 129.200 102.825 130.070 102.995 ;
        RECT 129.560 102.735 130.070 102.825 ;
        RECT 128.110 102.270 128.415 102.400 ;
        RECT 128.860 102.290 129.390 102.655 ;
        RECT 127.730 101.675 127.995 102.135 ;
        RECT 128.165 101.845 128.415 102.270 ;
        RECT 129.560 102.120 129.730 102.735 ;
        RECT 128.625 101.950 129.730 102.120 ;
        RECT 129.900 101.675 130.070 102.475 ;
        RECT 130.240 102.175 130.410 103.245 ;
        RECT 130.580 102.345 130.770 103.065 ;
        RECT 130.940 102.315 131.260 103.275 ;
        RECT 131.430 103.315 131.600 103.775 ;
        RECT 131.875 103.695 132.085 104.225 ;
        RECT 132.345 103.485 132.675 104.010 ;
        RECT 132.845 103.615 133.015 104.225 ;
        RECT 133.185 103.570 133.515 104.005 ;
        RECT 133.735 103.725 133.995 104.055 ;
        RECT 134.205 103.745 134.480 104.225 ;
        RECT 133.185 103.485 133.565 103.570 ;
        RECT 132.475 103.315 132.675 103.485 ;
        RECT 133.340 103.445 133.565 103.485 ;
        RECT 131.430 102.985 132.305 103.315 ;
        RECT 132.475 102.985 133.225 103.315 ;
        RECT 130.240 101.845 130.490 102.175 ;
        RECT 131.430 102.145 131.600 102.985 ;
        RECT 132.475 102.780 132.665 102.985 ;
        RECT 133.395 102.865 133.565 103.445 ;
        RECT 133.350 102.815 133.565 102.865 ;
        RECT 131.770 102.405 132.665 102.780 ;
        RECT 133.175 102.735 133.565 102.815 ;
        RECT 133.735 102.815 133.905 103.725 ;
        RECT 134.690 103.655 134.895 104.055 ;
        RECT 135.065 103.825 135.400 104.225 ;
        RECT 134.075 102.985 134.435 103.565 ;
        RECT 134.690 103.485 135.375 103.655 ;
        RECT 134.615 102.815 134.865 103.315 ;
        RECT 130.715 101.975 131.600 102.145 ;
        RECT 131.780 101.675 132.095 102.175 ;
        RECT 132.325 101.845 132.665 102.405 ;
        RECT 132.835 101.675 133.005 102.685 ;
        RECT 133.175 101.890 133.505 102.735 ;
        RECT 133.735 102.645 134.865 102.815 ;
        RECT 133.735 101.875 134.005 102.645 ;
        RECT 135.035 102.455 135.375 103.485 ;
        RECT 134.175 101.675 134.505 102.455 ;
        RECT 134.710 102.280 135.375 102.455 ;
        RECT 136.040 103.485 136.295 104.055 ;
        RECT 136.465 103.825 136.795 104.225 ;
        RECT 137.220 103.690 137.750 104.055 ;
        RECT 137.940 103.885 138.215 104.055 ;
        RECT 137.935 103.715 138.215 103.885 ;
        RECT 137.220 103.655 137.395 103.690 ;
        RECT 136.465 103.485 137.395 103.655 ;
        RECT 136.040 102.815 136.210 103.485 ;
        RECT 136.465 103.315 136.635 103.485 ;
        RECT 136.380 102.985 136.635 103.315 ;
        RECT 136.860 102.985 137.055 103.315 ;
        RECT 134.710 101.875 134.895 102.280 ;
        RECT 135.065 101.675 135.400 102.100 ;
        RECT 136.040 101.845 136.375 102.815 ;
        RECT 136.545 101.675 136.715 102.815 ;
        RECT 136.885 102.015 137.055 102.985 ;
        RECT 137.225 102.355 137.395 103.485 ;
        RECT 137.565 102.695 137.735 103.495 ;
        RECT 137.940 102.895 138.215 103.715 ;
        RECT 138.385 102.695 138.575 104.055 ;
        RECT 138.755 103.690 139.265 104.225 ;
        RECT 139.485 103.415 139.730 104.020 ;
        RECT 140.175 103.725 140.435 104.055 ;
        RECT 140.605 103.865 140.935 104.225 ;
        RECT 141.190 103.845 142.490 104.055 ;
        RECT 138.775 103.245 140.005 103.415 ;
        RECT 137.565 102.525 138.575 102.695 ;
        RECT 138.745 102.680 139.495 102.870 ;
        RECT 137.225 102.185 138.350 102.355 ;
        RECT 138.745 102.015 138.915 102.680 ;
        RECT 139.665 102.435 140.005 103.245 ;
        RECT 136.885 101.845 138.915 102.015 ;
        RECT 139.085 101.675 139.255 102.435 ;
        RECT 139.490 102.025 140.005 102.435 ;
        RECT 140.175 102.525 140.345 103.725 ;
        RECT 141.190 103.695 141.360 103.845 ;
        RECT 140.605 103.570 141.360 103.695 ;
        RECT 140.515 103.525 141.360 103.570 ;
        RECT 140.515 103.405 140.785 103.525 ;
        RECT 140.515 102.830 140.685 103.405 ;
        RECT 140.915 102.965 141.325 103.270 ;
        RECT 141.615 103.235 141.825 103.635 ;
        RECT 141.495 103.025 141.825 103.235 ;
        RECT 142.070 103.235 142.290 103.635 ;
        RECT 142.765 103.460 143.220 104.225 ;
        RECT 143.945 103.675 144.115 104.055 ;
        RECT 144.330 103.845 144.660 104.225 ;
        RECT 143.945 103.505 144.660 103.675 ;
        RECT 142.070 103.025 142.545 103.235 ;
        RECT 142.735 103.035 143.225 103.235 ;
        RECT 143.855 102.955 144.210 103.325 ;
        RECT 144.490 103.315 144.660 103.505 ;
        RECT 144.830 103.480 145.085 104.055 ;
        RECT 144.490 102.985 144.745 103.315 ;
        RECT 140.515 102.795 140.715 102.830 ;
        RECT 142.045 102.795 143.220 102.855 ;
        RECT 140.515 102.685 143.220 102.795 ;
        RECT 144.490 102.775 144.660 102.985 ;
        RECT 140.575 102.625 142.375 102.685 ;
        RECT 142.045 102.595 142.375 102.625 ;
        RECT 140.175 101.845 140.435 102.525 ;
        RECT 140.605 101.675 140.855 102.455 ;
        RECT 141.105 102.425 141.940 102.435 ;
        RECT 142.530 102.425 142.715 102.515 ;
        RECT 141.105 102.225 142.715 102.425 ;
        RECT 141.105 101.845 141.355 102.225 ;
        RECT 142.485 102.185 142.715 102.225 ;
        RECT 142.965 102.065 143.220 102.685 ;
        RECT 141.525 101.675 141.880 102.055 ;
        RECT 142.885 101.845 143.220 102.065 ;
        RECT 143.945 102.605 144.660 102.775 ;
        RECT 144.915 102.750 145.085 103.480 ;
        RECT 145.260 103.385 145.520 104.225 ;
        RECT 145.695 103.475 146.905 104.225 ;
        RECT 143.945 101.845 144.115 102.605 ;
        RECT 144.330 101.675 144.660 102.435 ;
        RECT 144.830 101.845 145.085 102.750 ;
        RECT 145.260 101.675 145.520 102.825 ;
        RECT 145.695 102.765 146.215 103.305 ;
        RECT 146.385 102.935 146.905 103.475 ;
        RECT 145.695 101.675 146.905 102.765 ;
        RECT 17.270 101.505 146.990 101.675 ;
        RECT 17.355 100.415 18.565 101.505 ;
        RECT 18.735 100.415 21.325 101.505 ;
        RECT 21.585 100.835 21.755 101.335 ;
        RECT 21.925 101.005 22.255 101.505 ;
        RECT 21.585 100.665 22.250 100.835 ;
        RECT 17.355 99.705 17.875 100.245 ;
        RECT 18.045 99.875 18.565 100.415 ;
        RECT 18.735 99.725 19.945 100.245 ;
        RECT 20.115 99.895 21.325 100.415 ;
        RECT 21.500 99.845 21.850 100.495 ;
        RECT 17.355 98.955 18.565 99.705 ;
        RECT 18.735 98.955 21.325 99.725 ;
        RECT 22.020 99.675 22.250 100.665 ;
        RECT 21.585 99.505 22.250 99.675 ;
        RECT 21.585 99.215 21.755 99.505 ;
        RECT 21.925 98.955 22.255 99.335 ;
        RECT 22.425 99.215 22.610 101.335 ;
        RECT 22.850 101.045 23.115 101.505 ;
        RECT 23.285 100.910 23.535 101.335 ;
        RECT 23.745 101.060 24.850 101.230 ;
        RECT 23.230 100.780 23.535 100.910 ;
        RECT 22.780 99.585 23.060 100.535 ;
        RECT 23.230 99.675 23.400 100.780 ;
        RECT 23.570 99.995 23.810 100.590 ;
        RECT 23.980 100.525 24.510 100.890 ;
        RECT 23.980 99.825 24.150 100.525 ;
        RECT 24.680 100.445 24.850 101.060 ;
        RECT 25.020 100.705 25.190 101.505 ;
        RECT 25.360 101.005 25.610 101.335 ;
        RECT 25.835 101.035 26.720 101.205 ;
        RECT 24.680 100.355 25.190 100.445 ;
        RECT 23.230 99.545 23.455 99.675 ;
        RECT 23.625 99.605 24.150 99.825 ;
        RECT 24.320 100.185 25.190 100.355 ;
        RECT 22.865 98.955 23.115 99.415 ;
        RECT 23.285 99.405 23.455 99.545 ;
        RECT 24.320 99.405 24.490 100.185 ;
        RECT 25.020 100.115 25.190 100.185 ;
        RECT 24.700 99.935 24.900 99.965 ;
        RECT 25.360 99.935 25.530 101.005 ;
        RECT 25.700 100.115 25.890 100.835 ;
        RECT 24.700 99.635 25.530 99.935 ;
        RECT 26.060 99.905 26.380 100.865 ;
        RECT 23.285 99.235 23.620 99.405 ;
        RECT 23.815 99.235 24.490 99.405 ;
        RECT 24.810 98.955 25.180 99.455 ;
        RECT 25.360 99.405 25.530 99.635 ;
        RECT 25.915 99.575 26.380 99.905 ;
        RECT 26.550 100.195 26.720 101.035 ;
        RECT 26.900 101.005 27.215 101.505 ;
        RECT 27.445 100.775 27.785 101.335 ;
        RECT 26.890 100.400 27.785 100.775 ;
        RECT 27.955 100.495 28.125 101.505 ;
        RECT 27.595 100.195 27.785 100.400 ;
        RECT 28.295 100.445 28.625 101.290 ;
        RECT 28.295 100.365 28.685 100.445 ;
        RECT 28.865 100.365 29.195 101.505 ;
        RECT 29.725 100.535 30.055 101.320 ;
        RECT 29.375 100.365 30.055 100.535 ;
        RECT 28.470 100.315 28.685 100.365 ;
        RECT 26.550 99.865 27.425 100.195 ;
        RECT 27.595 99.865 28.345 100.195 ;
        RECT 26.550 99.405 26.720 99.865 ;
        RECT 27.595 99.695 27.795 99.865 ;
        RECT 28.515 99.735 28.685 100.315 ;
        RECT 28.855 99.945 29.205 100.195 ;
        RECT 29.375 99.765 29.545 100.365 ;
        RECT 30.235 100.340 30.525 101.505 ;
        RECT 31.615 100.350 31.955 101.335 ;
        RECT 32.125 101.075 32.535 101.505 ;
        RECT 33.280 101.085 33.610 101.505 ;
        RECT 33.780 100.905 34.105 101.335 ;
        RECT 32.125 100.735 34.105 100.905 ;
        RECT 29.715 99.945 30.065 100.195 ;
        RECT 28.460 99.695 28.685 99.735 ;
        RECT 25.360 99.235 25.765 99.405 ;
        RECT 25.935 99.235 26.720 99.405 ;
        RECT 26.995 98.955 27.205 99.485 ;
        RECT 27.465 99.170 27.795 99.695 ;
        RECT 28.305 99.610 28.685 99.695 ;
        RECT 27.965 98.955 28.135 99.565 ;
        RECT 28.305 99.175 28.635 99.610 ;
        RECT 28.865 98.955 29.135 99.765 ;
        RECT 29.305 99.125 29.635 99.765 ;
        RECT 29.805 98.955 30.045 99.765 ;
        RECT 31.615 99.695 31.870 100.350 ;
        RECT 32.125 100.195 32.390 100.735 ;
        RECT 32.605 100.395 33.230 100.565 ;
        RECT 32.040 99.865 32.390 100.195 ;
        RECT 32.560 99.865 32.890 100.195 ;
        RECT 33.060 99.695 33.230 100.395 ;
        RECT 30.235 98.955 30.525 99.680 ;
        RECT 31.615 99.320 31.975 99.695 ;
        RECT 32.240 98.955 32.410 99.695 ;
        RECT 32.690 99.525 33.230 99.695 ;
        RECT 33.400 100.325 34.105 100.735 ;
        RECT 34.580 100.405 34.910 101.505 ;
        RECT 35.295 100.350 35.635 101.335 ;
        RECT 35.805 101.075 36.215 101.505 ;
        RECT 36.960 101.085 37.290 101.505 ;
        RECT 37.460 100.905 37.785 101.335 ;
        RECT 35.805 100.735 37.785 100.905 ;
        RECT 32.690 99.320 32.860 99.525 ;
        RECT 33.400 99.125 33.570 100.325 ;
        RECT 33.740 99.945 34.310 100.155 ;
        RECT 34.480 99.945 35.125 100.155 ;
        RECT 33.800 99.605 34.970 99.775 ;
        RECT 33.800 99.125 34.130 99.605 ;
        RECT 34.300 98.955 34.470 99.425 ;
        RECT 34.640 99.140 34.970 99.605 ;
        RECT 35.295 99.695 35.550 100.350 ;
        RECT 35.805 100.195 36.070 100.735 ;
        RECT 36.285 100.395 36.910 100.565 ;
        RECT 35.720 99.865 36.070 100.195 ;
        RECT 36.240 99.865 36.570 100.195 ;
        RECT 36.740 99.695 36.910 100.395 ;
        RECT 35.295 99.320 35.655 99.695 ;
        RECT 35.355 99.295 35.525 99.320 ;
        RECT 35.920 98.955 36.090 99.695 ;
        RECT 36.370 99.525 36.910 99.695 ;
        RECT 37.080 100.325 37.785 100.735 ;
        RECT 38.260 100.405 38.590 101.505 ;
        RECT 38.975 100.350 39.315 101.335 ;
        RECT 39.485 101.075 39.895 101.505 ;
        RECT 40.640 101.085 40.970 101.505 ;
        RECT 41.140 100.905 41.465 101.335 ;
        RECT 39.485 100.735 41.465 100.905 ;
        RECT 36.370 99.320 36.540 99.525 ;
        RECT 37.080 99.125 37.250 100.325 ;
        RECT 37.420 99.945 37.990 100.155 ;
        RECT 38.160 99.945 38.805 100.155 ;
        RECT 37.480 99.605 38.650 99.775 ;
        RECT 37.480 99.125 37.810 99.605 ;
        RECT 37.980 98.955 38.150 99.425 ;
        RECT 38.320 99.140 38.650 99.605 ;
        RECT 38.975 99.695 39.230 100.350 ;
        RECT 39.485 100.195 39.750 100.735 ;
        RECT 39.965 100.395 40.590 100.565 ;
        RECT 39.400 99.865 39.750 100.195 ;
        RECT 39.920 99.865 40.250 100.195 ;
        RECT 40.420 99.695 40.590 100.395 ;
        RECT 38.975 99.320 39.335 99.695 ;
        RECT 39.600 98.955 39.770 99.695 ;
        RECT 40.050 99.525 40.590 99.695 ;
        RECT 40.760 100.325 41.465 100.735 ;
        RECT 41.940 100.405 42.270 101.505 ;
        RECT 42.655 100.350 42.995 101.335 ;
        RECT 43.165 101.075 43.575 101.505 ;
        RECT 44.320 101.085 44.650 101.505 ;
        RECT 44.820 100.905 45.145 101.335 ;
        RECT 43.165 100.735 45.145 100.905 ;
        RECT 40.050 99.320 40.220 99.525 ;
        RECT 40.760 99.125 40.930 100.325 ;
        RECT 41.100 99.945 41.670 100.155 ;
        RECT 41.840 99.945 42.485 100.155 ;
        RECT 41.160 99.605 42.330 99.775 ;
        RECT 41.160 99.125 41.490 99.605 ;
        RECT 41.660 98.955 41.830 99.425 ;
        RECT 42.000 99.140 42.330 99.605 ;
        RECT 42.655 99.695 42.910 100.350 ;
        RECT 43.165 100.195 43.430 100.735 ;
        RECT 43.645 100.395 44.270 100.565 ;
        RECT 43.080 99.865 43.430 100.195 ;
        RECT 43.600 99.865 43.930 100.195 ;
        RECT 44.100 99.695 44.270 100.395 ;
        RECT 42.655 99.320 43.015 99.695 ;
        RECT 43.280 98.955 43.450 99.695 ;
        RECT 43.730 99.525 44.270 99.695 ;
        RECT 44.440 100.325 45.145 100.735 ;
        RECT 45.620 100.405 45.950 101.505 ;
        RECT 46.425 100.885 46.595 101.315 ;
        RECT 46.765 101.055 47.095 101.505 ;
        RECT 46.425 100.655 47.100 100.885 ;
        RECT 43.730 99.320 43.900 99.525 ;
        RECT 44.440 99.125 44.610 100.325 ;
        RECT 44.780 99.945 45.350 100.155 ;
        RECT 45.520 99.945 46.165 100.155 ;
        RECT 44.840 99.605 46.010 99.775 ;
        RECT 46.395 99.635 46.695 100.485 ;
        RECT 46.865 100.005 47.100 100.655 ;
        RECT 47.270 100.345 47.555 101.290 ;
        RECT 47.735 101.035 48.420 101.505 ;
        RECT 47.730 100.515 48.425 100.825 ;
        RECT 48.600 100.450 48.905 101.235 ;
        RECT 49.095 101.070 54.440 101.505 ;
        RECT 47.270 100.195 48.130 100.345 ;
        RECT 48.695 100.315 48.905 100.450 ;
        RECT 47.270 100.175 48.555 100.195 ;
        RECT 46.865 99.675 47.400 100.005 ;
        RECT 47.570 99.815 48.555 100.175 ;
        RECT 44.840 99.125 45.170 99.605 ;
        RECT 45.340 98.955 45.510 99.425 ;
        RECT 45.680 99.140 46.010 99.605 ;
        RECT 46.865 99.525 47.085 99.675 ;
        RECT 46.340 98.955 46.675 99.460 ;
        RECT 46.845 99.150 47.085 99.525 ;
        RECT 47.570 99.480 47.740 99.815 ;
        RECT 48.730 99.645 48.905 100.315 ;
        RECT 47.365 99.285 47.740 99.480 ;
        RECT 47.365 99.140 47.535 99.285 ;
        RECT 48.100 98.955 48.495 99.450 ;
        RECT 48.665 99.125 48.905 99.645 ;
        RECT 50.680 99.500 51.020 100.330 ;
        RECT 52.500 99.820 52.850 101.070 ;
        RECT 54.615 100.415 55.825 101.505 ;
        RECT 54.615 99.705 55.135 100.245 ;
        RECT 55.305 99.875 55.825 100.415 ;
        RECT 55.995 100.340 56.285 101.505 ;
        RECT 56.455 100.415 57.665 101.505 ;
        RECT 57.925 100.835 58.095 101.335 ;
        RECT 58.265 101.005 58.595 101.505 ;
        RECT 57.925 100.665 58.590 100.835 ;
        RECT 56.455 99.705 56.975 100.245 ;
        RECT 57.145 99.875 57.665 100.415 ;
        RECT 57.840 99.845 58.190 100.495 ;
        RECT 49.095 98.955 54.440 99.500 ;
        RECT 54.615 98.955 55.825 99.705 ;
        RECT 55.995 98.955 56.285 99.680 ;
        RECT 56.455 98.955 57.665 99.705 ;
        RECT 58.360 99.675 58.590 100.665 ;
        RECT 57.925 99.505 58.590 99.675 ;
        RECT 57.925 99.215 58.095 99.505 ;
        RECT 58.265 98.955 58.595 99.335 ;
        RECT 58.765 99.215 58.950 101.335 ;
        RECT 59.190 101.045 59.455 101.505 ;
        RECT 59.625 100.910 59.875 101.335 ;
        RECT 60.085 101.060 61.190 101.230 ;
        RECT 59.570 100.780 59.875 100.910 ;
        RECT 59.120 99.585 59.400 100.535 ;
        RECT 59.570 99.675 59.740 100.780 ;
        RECT 59.910 99.995 60.150 100.590 ;
        RECT 60.320 100.525 60.850 100.890 ;
        RECT 60.320 99.825 60.490 100.525 ;
        RECT 61.020 100.445 61.190 101.060 ;
        RECT 61.360 100.705 61.530 101.505 ;
        RECT 61.700 101.005 61.950 101.335 ;
        RECT 62.175 101.035 63.060 101.205 ;
        RECT 61.020 100.355 61.530 100.445 ;
        RECT 59.570 99.545 59.795 99.675 ;
        RECT 59.965 99.605 60.490 99.825 ;
        RECT 60.660 100.185 61.530 100.355 ;
        RECT 59.205 98.955 59.455 99.415 ;
        RECT 59.625 99.405 59.795 99.545 ;
        RECT 60.660 99.405 60.830 100.185 ;
        RECT 61.360 100.115 61.530 100.185 ;
        RECT 61.040 99.935 61.240 99.965 ;
        RECT 61.700 99.935 61.870 101.005 ;
        RECT 62.040 100.115 62.230 100.835 ;
        RECT 61.040 99.635 61.870 99.935 ;
        RECT 62.400 99.905 62.720 100.865 ;
        RECT 59.625 99.235 59.960 99.405 ;
        RECT 60.155 99.235 60.830 99.405 ;
        RECT 61.150 98.955 61.520 99.455 ;
        RECT 61.700 99.405 61.870 99.635 ;
        RECT 62.255 99.575 62.720 99.905 ;
        RECT 62.890 100.195 63.060 101.035 ;
        RECT 63.240 101.005 63.555 101.505 ;
        RECT 63.785 100.775 64.125 101.335 ;
        RECT 63.230 100.400 64.125 100.775 ;
        RECT 64.295 100.495 64.465 101.505 ;
        RECT 63.935 100.195 64.125 100.400 ;
        RECT 64.635 100.445 64.965 101.290 ;
        RECT 65.285 100.835 65.455 101.335 ;
        RECT 65.625 101.005 65.955 101.505 ;
        RECT 65.285 100.665 65.950 100.835 ;
        RECT 64.635 100.365 65.025 100.445 ;
        RECT 64.810 100.315 65.025 100.365 ;
        RECT 62.890 99.865 63.765 100.195 ;
        RECT 63.935 99.865 64.685 100.195 ;
        RECT 62.890 99.405 63.060 99.865 ;
        RECT 63.935 99.695 64.135 99.865 ;
        RECT 64.855 99.735 65.025 100.315 ;
        RECT 65.200 99.845 65.550 100.495 ;
        RECT 64.800 99.695 65.025 99.735 ;
        RECT 61.700 99.235 62.105 99.405 ;
        RECT 62.275 99.235 63.060 99.405 ;
        RECT 63.335 98.955 63.545 99.485 ;
        RECT 63.805 99.170 64.135 99.695 ;
        RECT 64.645 99.610 65.025 99.695 ;
        RECT 65.720 99.675 65.950 100.665 ;
        RECT 64.305 98.955 64.475 99.565 ;
        RECT 64.645 99.175 64.975 99.610 ;
        RECT 65.285 99.505 65.950 99.675 ;
        RECT 65.285 99.215 65.455 99.505 ;
        RECT 65.625 98.955 65.955 99.335 ;
        RECT 66.125 99.215 66.310 101.335 ;
        RECT 66.550 101.045 66.815 101.505 ;
        RECT 66.985 100.910 67.235 101.335 ;
        RECT 67.445 101.060 68.550 101.230 ;
        RECT 66.930 100.780 67.235 100.910 ;
        RECT 66.480 99.585 66.760 100.535 ;
        RECT 66.930 99.675 67.100 100.780 ;
        RECT 67.270 99.995 67.510 100.590 ;
        RECT 67.680 100.525 68.210 100.890 ;
        RECT 67.680 99.825 67.850 100.525 ;
        RECT 68.380 100.445 68.550 101.060 ;
        RECT 68.720 100.705 68.890 101.505 ;
        RECT 69.060 101.005 69.310 101.335 ;
        RECT 69.535 101.035 70.420 101.205 ;
        RECT 68.380 100.355 68.890 100.445 ;
        RECT 66.930 99.545 67.155 99.675 ;
        RECT 67.325 99.605 67.850 99.825 ;
        RECT 68.020 100.185 68.890 100.355 ;
        RECT 66.565 98.955 66.815 99.415 ;
        RECT 66.985 99.405 67.155 99.545 ;
        RECT 68.020 99.405 68.190 100.185 ;
        RECT 68.720 100.115 68.890 100.185 ;
        RECT 68.400 99.935 68.600 99.965 ;
        RECT 69.060 99.935 69.230 101.005 ;
        RECT 69.400 100.115 69.590 100.835 ;
        RECT 68.400 99.635 69.230 99.935 ;
        RECT 69.760 99.905 70.080 100.865 ;
        RECT 66.985 99.235 67.320 99.405 ;
        RECT 67.515 99.235 68.190 99.405 ;
        RECT 68.510 98.955 68.880 99.455 ;
        RECT 69.060 99.405 69.230 99.635 ;
        RECT 69.615 99.575 70.080 99.905 ;
        RECT 70.250 100.195 70.420 101.035 ;
        RECT 70.600 101.005 70.915 101.505 ;
        RECT 71.145 100.775 71.485 101.335 ;
        RECT 70.590 100.400 71.485 100.775 ;
        RECT 71.655 100.495 71.825 101.505 ;
        RECT 71.295 100.195 71.485 100.400 ;
        RECT 71.995 100.445 72.325 101.290 ;
        RECT 72.645 100.575 72.815 101.335 ;
        RECT 73.030 100.745 73.360 101.505 ;
        RECT 71.995 100.365 72.385 100.445 ;
        RECT 72.645 100.405 73.360 100.575 ;
        RECT 73.530 100.430 73.785 101.335 ;
        RECT 72.170 100.315 72.385 100.365 ;
        RECT 70.250 99.865 71.125 100.195 ;
        RECT 71.295 99.865 72.045 100.195 ;
        RECT 70.250 99.405 70.420 99.865 ;
        RECT 71.295 99.695 71.495 99.865 ;
        RECT 72.215 99.735 72.385 100.315 ;
        RECT 72.555 99.855 72.910 100.225 ;
        RECT 73.190 100.195 73.360 100.405 ;
        RECT 73.190 99.865 73.445 100.195 ;
        RECT 72.160 99.695 72.385 99.735 ;
        RECT 69.060 99.235 69.465 99.405 ;
        RECT 69.635 99.235 70.420 99.405 ;
        RECT 70.695 98.955 70.905 99.485 ;
        RECT 71.165 99.170 71.495 99.695 ;
        RECT 72.005 99.610 72.385 99.695 ;
        RECT 73.190 99.675 73.360 99.865 ;
        RECT 73.615 99.700 73.785 100.430 ;
        RECT 73.960 100.355 74.220 101.505 ;
        RECT 74.485 100.835 74.655 101.335 ;
        RECT 74.825 101.005 75.155 101.505 ;
        RECT 74.485 100.665 75.150 100.835 ;
        RECT 74.400 99.845 74.750 100.495 ;
        RECT 71.665 98.955 71.835 99.565 ;
        RECT 72.005 99.175 72.335 99.610 ;
        RECT 72.645 99.505 73.360 99.675 ;
        RECT 72.645 99.125 72.815 99.505 ;
        RECT 73.030 98.955 73.360 99.335 ;
        RECT 73.530 99.125 73.785 99.700 ;
        RECT 73.960 98.955 74.220 99.795 ;
        RECT 74.920 99.675 75.150 100.665 ;
        RECT 74.485 99.505 75.150 99.675 ;
        RECT 74.485 99.215 74.655 99.505 ;
        RECT 74.825 98.955 75.155 99.335 ;
        RECT 75.325 99.215 75.510 101.335 ;
        RECT 75.750 101.045 76.015 101.505 ;
        RECT 76.185 100.910 76.435 101.335 ;
        RECT 76.645 101.060 77.750 101.230 ;
        RECT 76.130 100.780 76.435 100.910 ;
        RECT 75.680 99.585 75.960 100.535 ;
        RECT 76.130 99.675 76.300 100.780 ;
        RECT 76.470 99.995 76.710 100.590 ;
        RECT 76.880 100.525 77.410 100.890 ;
        RECT 76.880 99.825 77.050 100.525 ;
        RECT 77.580 100.445 77.750 101.060 ;
        RECT 77.920 100.705 78.090 101.505 ;
        RECT 78.260 101.005 78.510 101.335 ;
        RECT 78.735 101.035 79.620 101.205 ;
        RECT 77.580 100.355 78.090 100.445 ;
        RECT 76.130 99.545 76.355 99.675 ;
        RECT 76.525 99.605 77.050 99.825 ;
        RECT 77.220 100.185 78.090 100.355 ;
        RECT 75.765 98.955 76.015 99.415 ;
        RECT 76.185 99.405 76.355 99.545 ;
        RECT 77.220 99.405 77.390 100.185 ;
        RECT 77.920 100.115 78.090 100.185 ;
        RECT 77.600 99.935 77.800 99.965 ;
        RECT 78.260 99.935 78.430 101.005 ;
        RECT 78.600 100.115 78.790 100.835 ;
        RECT 77.600 99.635 78.430 99.935 ;
        RECT 78.960 99.905 79.280 100.865 ;
        RECT 76.185 99.235 76.520 99.405 ;
        RECT 76.715 99.235 77.390 99.405 ;
        RECT 77.710 98.955 78.080 99.455 ;
        RECT 78.260 99.405 78.430 99.635 ;
        RECT 78.815 99.575 79.280 99.905 ;
        RECT 79.450 100.195 79.620 101.035 ;
        RECT 79.800 101.005 80.115 101.505 ;
        RECT 80.345 100.775 80.685 101.335 ;
        RECT 79.790 100.400 80.685 100.775 ;
        RECT 80.855 100.495 81.025 101.505 ;
        RECT 80.495 100.195 80.685 100.400 ;
        RECT 81.195 100.445 81.525 101.290 ;
        RECT 81.195 100.365 81.585 100.445 ;
        RECT 81.370 100.315 81.585 100.365 ;
        RECT 81.755 100.340 82.045 101.505 ;
        RECT 82.220 101.115 82.555 101.335 ;
        RECT 83.560 101.125 83.915 101.505 ;
        RECT 82.220 100.495 82.475 101.115 ;
        RECT 82.725 100.955 82.955 100.995 ;
        RECT 84.085 100.955 84.335 101.335 ;
        RECT 82.725 100.755 84.335 100.955 ;
        RECT 82.725 100.665 82.910 100.755 ;
        RECT 83.500 100.745 84.335 100.755 ;
        RECT 84.585 100.725 84.835 101.505 ;
        RECT 85.005 100.655 85.265 101.335 ;
        RECT 83.065 100.555 83.395 100.585 ;
        RECT 83.065 100.495 84.865 100.555 ;
        RECT 82.220 100.385 84.925 100.495 ;
        RECT 82.220 100.325 83.395 100.385 ;
        RECT 84.725 100.350 84.925 100.385 ;
        RECT 79.450 99.865 80.325 100.195 ;
        RECT 80.495 99.865 81.245 100.195 ;
        RECT 79.450 99.405 79.620 99.865 ;
        RECT 80.495 99.695 80.695 99.865 ;
        RECT 81.415 99.735 81.585 100.315 ;
        RECT 82.215 99.945 82.705 100.145 ;
        RECT 82.895 99.945 83.370 100.155 ;
        RECT 81.360 99.695 81.585 99.735 ;
        RECT 78.260 99.235 78.665 99.405 ;
        RECT 78.835 99.235 79.620 99.405 ;
        RECT 79.895 98.955 80.105 99.485 ;
        RECT 80.365 99.170 80.695 99.695 ;
        RECT 81.205 99.610 81.585 99.695 ;
        RECT 80.865 98.955 81.035 99.565 ;
        RECT 81.205 99.175 81.535 99.610 ;
        RECT 81.755 98.955 82.045 99.680 ;
        RECT 82.220 98.955 82.675 99.720 ;
        RECT 83.150 99.545 83.370 99.945 ;
        RECT 83.615 99.945 83.945 100.155 ;
        RECT 83.615 99.545 83.825 99.945 ;
        RECT 84.115 99.910 84.525 100.215 ;
        RECT 84.755 99.775 84.925 100.350 ;
        RECT 84.655 99.655 84.925 99.775 ;
        RECT 84.080 99.610 84.925 99.655 ;
        RECT 84.080 99.485 84.835 99.610 ;
        RECT 84.080 99.335 84.250 99.485 ;
        RECT 85.095 99.455 85.265 100.655 ;
        RECT 85.435 100.415 87.105 101.505 ;
        RECT 87.365 100.835 87.535 101.335 ;
        RECT 87.705 101.005 88.035 101.505 ;
        RECT 87.365 100.665 88.030 100.835 ;
        RECT 82.950 99.125 84.250 99.335 ;
        RECT 84.505 98.955 84.835 99.315 ;
        RECT 85.005 99.125 85.265 99.455 ;
        RECT 85.435 99.725 86.185 100.245 ;
        RECT 86.355 99.895 87.105 100.415 ;
        RECT 87.280 99.845 87.630 100.495 ;
        RECT 85.435 98.955 87.105 99.725 ;
        RECT 87.800 99.675 88.030 100.665 ;
        RECT 87.365 99.505 88.030 99.675 ;
        RECT 87.365 99.215 87.535 99.505 ;
        RECT 87.705 98.955 88.035 99.335 ;
        RECT 88.205 99.215 88.390 101.335 ;
        RECT 88.630 101.045 88.895 101.505 ;
        RECT 89.065 100.910 89.315 101.335 ;
        RECT 89.525 101.060 90.630 101.230 ;
        RECT 89.010 100.780 89.315 100.910 ;
        RECT 88.560 99.585 88.840 100.535 ;
        RECT 89.010 99.675 89.180 100.780 ;
        RECT 89.350 99.995 89.590 100.590 ;
        RECT 89.760 100.525 90.290 100.890 ;
        RECT 89.760 99.825 89.930 100.525 ;
        RECT 90.460 100.445 90.630 101.060 ;
        RECT 90.800 100.705 90.970 101.505 ;
        RECT 91.140 101.005 91.390 101.335 ;
        RECT 91.615 101.035 92.500 101.205 ;
        RECT 90.460 100.355 90.970 100.445 ;
        RECT 89.010 99.545 89.235 99.675 ;
        RECT 89.405 99.605 89.930 99.825 ;
        RECT 90.100 100.185 90.970 100.355 ;
        RECT 88.645 98.955 88.895 99.415 ;
        RECT 89.065 99.405 89.235 99.545 ;
        RECT 90.100 99.405 90.270 100.185 ;
        RECT 90.800 100.115 90.970 100.185 ;
        RECT 90.480 99.935 90.680 99.965 ;
        RECT 91.140 99.935 91.310 101.005 ;
        RECT 91.480 100.115 91.670 100.835 ;
        RECT 90.480 99.635 91.310 99.935 ;
        RECT 91.840 99.905 92.160 100.865 ;
        RECT 89.065 99.235 89.400 99.405 ;
        RECT 89.595 99.235 90.270 99.405 ;
        RECT 90.590 98.955 90.960 99.455 ;
        RECT 91.140 99.405 91.310 99.635 ;
        RECT 91.695 99.575 92.160 99.905 ;
        RECT 92.330 100.195 92.500 101.035 ;
        RECT 92.680 101.005 92.995 101.505 ;
        RECT 93.225 100.775 93.565 101.335 ;
        RECT 92.670 100.400 93.565 100.775 ;
        RECT 93.735 100.495 93.905 101.505 ;
        RECT 93.375 100.195 93.565 100.400 ;
        RECT 94.075 100.445 94.405 101.290 ;
        RECT 94.075 100.365 94.465 100.445 ;
        RECT 94.250 100.315 94.465 100.365 ;
        RECT 92.330 99.865 93.205 100.195 ;
        RECT 93.375 99.865 94.125 100.195 ;
        RECT 92.330 99.405 92.500 99.865 ;
        RECT 93.375 99.695 93.575 99.865 ;
        RECT 94.295 99.735 94.465 100.315 ;
        RECT 94.240 99.695 94.465 99.735 ;
        RECT 91.140 99.235 91.545 99.405 ;
        RECT 91.715 99.235 92.500 99.405 ;
        RECT 92.775 98.955 92.985 99.485 ;
        RECT 93.245 99.170 93.575 99.695 ;
        RECT 94.085 99.610 94.465 99.695 ;
        RECT 94.635 100.430 94.905 101.335 ;
        RECT 95.075 100.745 95.405 101.505 ;
        RECT 95.585 100.575 95.765 101.335 ;
        RECT 96.105 100.835 96.275 101.335 ;
        RECT 96.445 101.005 96.775 101.505 ;
        RECT 96.105 100.665 96.770 100.835 ;
        RECT 94.635 99.630 94.815 100.430 ;
        RECT 95.090 100.405 95.765 100.575 ;
        RECT 95.090 100.260 95.260 100.405 ;
        RECT 94.985 99.930 95.260 100.260 ;
        RECT 95.090 99.675 95.260 99.930 ;
        RECT 95.485 99.855 95.825 100.225 ;
        RECT 96.020 99.845 96.370 100.495 ;
        RECT 96.540 99.675 96.770 100.665 ;
        RECT 93.745 98.955 93.915 99.565 ;
        RECT 94.085 99.175 94.415 99.610 ;
        RECT 94.635 99.125 94.895 99.630 ;
        RECT 95.090 99.505 95.755 99.675 ;
        RECT 95.075 98.955 95.405 99.335 ;
        RECT 95.585 99.125 95.755 99.505 ;
        RECT 96.105 99.505 96.770 99.675 ;
        RECT 96.105 99.215 96.275 99.505 ;
        RECT 96.445 98.955 96.775 99.335 ;
        RECT 96.945 99.215 97.130 101.335 ;
        RECT 97.370 101.045 97.635 101.505 ;
        RECT 97.805 100.910 98.055 101.335 ;
        RECT 98.265 101.060 99.370 101.230 ;
        RECT 97.750 100.780 98.055 100.910 ;
        RECT 97.300 99.585 97.580 100.535 ;
        RECT 97.750 99.675 97.920 100.780 ;
        RECT 98.090 99.995 98.330 100.590 ;
        RECT 98.500 100.525 99.030 100.890 ;
        RECT 98.500 99.825 98.670 100.525 ;
        RECT 99.200 100.445 99.370 101.060 ;
        RECT 99.540 100.705 99.710 101.505 ;
        RECT 99.880 101.005 100.130 101.335 ;
        RECT 100.355 101.035 101.240 101.205 ;
        RECT 99.200 100.355 99.710 100.445 ;
        RECT 97.750 99.545 97.975 99.675 ;
        RECT 98.145 99.605 98.670 99.825 ;
        RECT 98.840 100.185 99.710 100.355 ;
        RECT 97.385 98.955 97.635 99.415 ;
        RECT 97.805 99.405 97.975 99.545 ;
        RECT 98.840 99.405 99.010 100.185 ;
        RECT 99.540 100.115 99.710 100.185 ;
        RECT 99.220 99.935 99.420 99.965 ;
        RECT 99.880 99.935 100.050 101.005 ;
        RECT 100.220 100.115 100.410 100.835 ;
        RECT 99.220 99.635 100.050 99.935 ;
        RECT 100.580 99.905 100.900 100.865 ;
        RECT 97.805 99.235 98.140 99.405 ;
        RECT 98.335 99.235 99.010 99.405 ;
        RECT 99.330 98.955 99.700 99.455 ;
        RECT 99.880 99.405 100.050 99.635 ;
        RECT 100.435 99.575 100.900 99.905 ;
        RECT 101.070 100.195 101.240 101.035 ;
        RECT 101.420 101.005 101.735 101.505 ;
        RECT 101.965 100.775 102.305 101.335 ;
        RECT 101.410 100.400 102.305 100.775 ;
        RECT 102.475 100.495 102.645 101.505 ;
        RECT 102.115 100.195 102.305 100.400 ;
        RECT 102.815 100.445 103.145 101.290 ;
        RECT 103.465 100.495 103.635 101.335 ;
        RECT 103.805 101.165 104.975 101.335 ;
        RECT 103.805 100.665 104.135 101.165 ;
        RECT 104.645 101.125 104.975 101.165 ;
        RECT 105.165 101.085 105.520 101.505 ;
        RECT 104.305 100.905 104.535 100.995 ;
        RECT 105.690 100.905 105.940 101.335 ;
        RECT 104.305 100.665 105.940 100.905 ;
        RECT 106.110 100.745 106.440 101.505 ;
        RECT 106.610 100.665 106.865 101.335 ;
        RECT 102.815 100.365 103.205 100.445 ;
        RECT 102.990 100.315 103.205 100.365 ;
        RECT 103.465 100.325 106.525 100.495 ;
        RECT 101.070 99.865 101.945 100.195 ;
        RECT 102.115 99.865 102.865 100.195 ;
        RECT 101.070 99.405 101.240 99.865 ;
        RECT 102.115 99.695 102.315 99.865 ;
        RECT 103.035 99.735 103.205 100.315 ;
        RECT 103.380 99.945 103.730 100.155 ;
        RECT 103.900 99.945 104.345 100.145 ;
        RECT 104.515 99.945 104.990 100.145 ;
        RECT 102.980 99.695 103.205 99.735 ;
        RECT 99.880 99.235 100.285 99.405 ;
        RECT 100.455 99.235 101.240 99.405 ;
        RECT 101.515 98.955 101.725 99.485 ;
        RECT 101.985 99.170 102.315 99.695 ;
        RECT 102.825 99.610 103.205 99.695 ;
        RECT 102.485 98.955 102.655 99.565 ;
        RECT 102.825 99.175 103.155 99.610 ;
        RECT 103.465 99.605 104.530 99.775 ;
        RECT 103.465 99.125 103.635 99.605 ;
        RECT 103.805 98.955 104.135 99.435 ;
        RECT 104.360 99.375 104.530 99.605 ;
        RECT 104.710 99.545 104.990 99.945 ;
        RECT 105.260 99.945 105.590 100.145 ;
        RECT 105.760 99.945 106.125 100.145 ;
        RECT 105.260 99.545 105.545 99.945 ;
        RECT 106.355 99.775 106.525 100.325 ;
        RECT 105.725 99.605 106.525 99.775 ;
        RECT 105.725 99.375 105.895 99.605 ;
        RECT 106.695 99.535 106.865 100.665 ;
        RECT 107.515 100.340 107.805 101.505 ;
        RECT 108.065 100.835 108.235 101.335 ;
        RECT 108.405 101.005 108.735 101.505 ;
        RECT 108.065 100.665 108.730 100.835 ;
        RECT 107.980 99.845 108.330 100.495 ;
        RECT 106.680 99.455 106.865 99.535 ;
        RECT 104.360 99.125 105.895 99.375 ;
        RECT 106.065 98.955 106.395 99.435 ;
        RECT 106.610 99.125 106.865 99.455 ;
        RECT 107.515 98.955 107.805 99.680 ;
        RECT 108.500 99.675 108.730 100.665 ;
        RECT 108.065 99.505 108.730 99.675 ;
        RECT 108.065 99.215 108.235 99.505 ;
        RECT 108.405 98.955 108.735 99.335 ;
        RECT 108.905 99.215 109.090 101.335 ;
        RECT 109.330 101.045 109.595 101.505 ;
        RECT 109.765 100.910 110.015 101.335 ;
        RECT 110.225 101.060 111.330 101.230 ;
        RECT 109.710 100.780 110.015 100.910 ;
        RECT 109.260 99.585 109.540 100.535 ;
        RECT 109.710 99.675 109.880 100.780 ;
        RECT 110.050 99.995 110.290 100.590 ;
        RECT 110.460 100.525 110.990 100.890 ;
        RECT 110.460 99.825 110.630 100.525 ;
        RECT 111.160 100.445 111.330 101.060 ;
        RECT 111.500 100.705 111.670 101.505 ;
        RECT 111.840 101.005 112.090 101.335 ;
        RECT 112.315 101.035 113.200 101.205 ;
        RECT 111.160 100.355 111.670 100.445 ;
        RECT 109.710 99.545 109.935 99.675 ;
        RECT 110.105 99.605 110.630 99.825 ;
        RECT 110.800 100.185 111.670 100.355 ;
        RECT 109.345 98.955 109.595 99.415 ;
        RECT 109.765 99.405 109.935 99.545 ;
        RECT 110.800 99.405 110.970 100.185 ;
        RECT 111.500 100.115 111.670 100.185 ;
        RECT 111.180 99.935 111.380 99.965 ;
        RECT 111.840 99.935 112.010 101.005 ;
        RECT 112.180 100.115 112.370 100.835 ;
        RECT 111.180 99.635 112.010 99.935 ;
        RECT 112.540 99.905 112.860 100.865 ;
        RECT 109.765 99.235 110.100 99.405 ;
        RECT 110.295 99.235 110.970 99.405 ;
        RECT 111.290 98.955 111.660 99.455 ;
        RECT 111.840 99.405 112.010 99.635 ;
        RECT 112.395 99.575 112.860 99.905 ;
        RECT 113.030 100.195 113.200 101.035 ;
        RECT 113.380 101.005 113.695 101.505 ;
        RECT 113.925 100.775 114.265 101.335 ;
        RECT 113.370 100.400 114.265 100.775 ;
        RECT 114.435 100.495 114.605 101.505 ;
        RECT 114.075 100.195 114.265 100.400 ;
        RECT 114.775 100.445 115.105 101.290 ;
        RECT 115.425 100.835 115.595 101.335 ;
        RECT 115.765 101.005 116.095 101.505 ;
        RECT 115.425 100.665 116.090 100.835 ;
        RECT 114.775 100.365 115.165 100.445 ;
        RECT 114.950 100.315 115.165 100.365 ;
        RECT 113.030 99.865 113.905 100.195 ;
        RECT 114.075 99.865 114.825 100.195 ;
        RECT 113.030 99.405 113.200 99.865 ;
        RECT 114.075 99.695 114.275 99.865 ;
        RECT 114.995 99.735 115.165 100.315 ;
        RECT 115.340 99.845 115.690 100.495 ;
        RECT 114.940 99.695 115.165 99.735 ;
        RECT 111.840 99.235 112.245 99.405 ;
        RECT 112.415 99.235 113.200 99.405 ;
        RECT 113.475 98.955 113.685 99.485 ;
        RECT 113.945 99.170 114.275 99.695 ;
        RECT 114.785 99.610 115.165 99.695 ;
        RECT 115.860 99.675 116.090 100.665 ;
        RECT 114.445 98.955 114.615 99.565 ;
        RECT 114.785 99.175 115.115 99.610 ;
        RECT 115.425 99.505 116.090 99.675 ;
        RECT 115.425 99.215 115.595 99.505 ;
        RECT 115.765 98.955 116.095 99.335 ;
        RECT 116.265 99.215 116.450 101.335 ;
        RECT 116.690 101.045 116.955 101.505 ;
        RECT 117.125 100.910 117.375 101.335 ;
        RECT 117.585 101.060 118.690 101.230 ;
        RECT 117.070 100.780 117.375 100.910 ;
        RECT 116.620 99.585 116.900 100.535 ;
        RECT 117.070 99.675 117.240 100.780 ;
        RECT 117.410 99.995 117.650 100.590 ;
        RECT 117.820 100.525 118.350 100.890 ;
        RECT 117.820 99.825 117.990 100.525 ;
        RECT 118.520 100.445 118.690 101.060 ;
        RECT 118.860 100.705 119.030 101.505 ;
        RECT 119.200 101.005 119.450 101.335 ;
        RECT 119.675 101.035 120.560 101.205 ;
        RECT 118.520 100.355 119.030 100.445 ;
        RECT 117.070 99.545 117.295 99.675 ;
        RECT 117.465 99.605 117.990 99.825 ;
        RECT 118.160 100.185 119.030 100.355 ;
        RECT 116.705 98.955 116.955 99.415 ;
        RECT 117.125 99.405 117.295 99.545 ;
        RECT 118.160 99.405 118.330 100.185 ;
        RECT 118.860 100.115 119.030 100.185 ;
        RECT 118.540 99.935 118.740 99.965 ;
        RECT 119.200 99.935 119.370 101.005 ;
        RECT 119.540 100.115 119.730 100.835 ;
        RECT 118.540 99.635 119.370 99.935 ;
        RECT 119.900 99.905 120.220 100.865 ;
        RECT 117.125 99.235 117.460 99.405 ;
        RECT 117.655 99.235 118.330 99.405 ;
        RECT 118.650 98.955 119.020 99.455 ;
        RECT 119.200 99.405 119.370 99.635 ;
        RECT 119.755 99.575 120.220 99.905 ;
        RECT 120.390 100.195 120.560 101.035 ;
        RECT 120.740 101.005 121.055 101.505 ;
        RECT 121.285 100.775 121.625 101.335 ;
        RECT 120.730 100.400 121.625 100.775 ;
        RECT 121.795 100.495 121.965 101.505 ;
        RECT 121.435 100.195 121.625 100.400 ;
        RECT 122.135 100.445 122.465 101.290 ;
        RECT 122.785 100.835 122.955 101.335 ;
        RECT 123.125 101.005 123.455 101.505 ;
        RECT 122.785 100.665 123.450 100.835 ;
        RECT 122.135 100.365 122.525 100.445 ;
        RECT 122.310 100.315 122.525 100.365 ;
        RECT 120.390 99.865 121.265 100.195 ;
        RECT 121.435 99.865 122.185 100.195 ;
        RECT 120.390 99.405 120.560 99.865 ;
        RECT 121.435 99.695 121.635 99.865 ;
        RECT 122.355 99.735 122.525 100.315 ;
        RECT 122.700 99.845 123.050 100.495 ;
        RECT 122.300 99.695 122.525 99.735 ;
        RECT 119.200 99.235 119.605 99.405 ;
        RECT 119.775 99.235 120.560 99.405 ;
        RECT 120.835 98.955 121.045 99.485 ;
        RECT 121.305 99.170 121.635 99.695 ;
        RECT 122.145 99.610 122.525 99.695 ;
        RECT 123.220 99.675 123.450 100.665 ;
        RECT 121.805 98.955 121.975 99.565 ;
        RECT 122.145 99.175 122.475 99.610 ;
        RECT 122.785 99.505 123.450 99.675 ;
        RECT 122.785 99.215 122.955 99.505 ;
        RECT 123.125 98.955 123.455 99.335 ;
        RECT 123.625 99.215 123.810 101.335 ;
        RECT 124.050 101.045 124.315 101.505 ;
        RECT 124.485 100.910 124.735 101.335 ;
        RECT 124.945 101.060 126.050 101.230 ;
        RECT 124.430 100.780 124.735 100.910 ;
        RECT 123.980 99.585 124.260 100.535 ;
        RECT 124.430 99.675 124.600 100.780 ;
        RECT 124.770 99.995 125.010 100.590 ;
        RECT 125.180 100.525 125.710 100.890 ;
        RECT 125.180 99.825 125.350 100.525 ;
        RECT 125.880 100.445 126.050 101.060 ;
        RECT 126.220 100.705 126.390 101.505 ;
        RECT 126.560 101.005 126.810 101.335 ;
        RECT 127.035 101.035 127.920 101.205 ;
        RECT 125.880 100.355 126.390 100.445 ;
        RECT 124.430 99.545 124.655 99.675 ;
        RECT 124.825 99.605 125.350 99.825 ;
        RECT 125.520 100.185 126.390 100.355 ;
        RECT 124.065 98.955 124.315 99.415 ;
        RECT 124.485 99.405 124.655 99.545 ;
        RECT 125.520 99.405 125.690 100.185 ;
        RECT 126.220 100.115 126.390 100.185 ;
        RECT 125.900 99.935 126.100 99.965 ;
        RECT 126.560 99.935 126.730 101.005 ;
        RECT 126.900 100.115 127.090 100.835 ;
        RECT 125.900 99.635 126.730 99.935 ;
        RECT 127.260 99.905 127.580 100.865 ;
        RECT 124.485 99.235 124.820 99.405 ;
        RECT 125.015 99.235 125.690 99.405 ;
        RECT 126.010 98.955 126.380 99.455 ;
        RECT 126.560 99.405 126.730 99.635 ;
        RECT 127.115 99.575 127.580 99.905 ;
        RECT 127.750 100.195 127.920 101.035 ;
        RECT 128.100 101.005 128.415 101.505 ;
        RECT 128.645 100.775 128.985 101.335 ;
        RECT 128.090 100.400 128.985 100.775 ;
        RECT 129.155 100.495 129.325 101.505 ;
        RECT 128.795 100.195 128.985 100.400 ;
        RECT 129.495 100.445 129.825 101.290 ;
        RECT 130.075 100.450 130.380 101.235 ;
        RECT 130.560 101.035 131.245 101.505 ;
        RECT 130.555 100.515 131.250 100.825 ;
        RECT 129.495 100.365 129.885 100.445 ;
        RECT 129.670 100.315 129.885 100.365 ;
        RECT 127.750 99.865 128.625 100.195 ;
        RECT 128.795 99.865 129.545 100.195 ;
        RECT 127.750 99.405 127.920 99.865 ;
        RECT 128.795 99.695 128.995 99.865 ;
        RECT 129.715 99.735 129.885 100.315 ;
        RECT 129.660 99.695 129.885 99.735 ;
        RECT 126.560 99.235 126.965 99.405 ;
        RECT 127.135 99.235 127.920 99.405 ;
        RECT 128.195 98.955 128.405 99.485 ;
        RECT 128.665 99.170 128.995 99.695 ;
        RECT 129.505 99.610 129.885 99.695 ;
        RECT 130.075 99.645 130.250 100.450 ;
        RECT 131.425 100.345 131.710 101.290 ;
        RECT 131.885 101.055 132.215 101.505 ;
        RECT 132.385 100.885 132.555 101.315 ;
        RECT 130.850 100.195 131.710 100.345 ;
        RECT 130.425 100.175 131.710 100.195 ;
        RECT 131.880 100.655 132.555 100.885 ;
        RECT 130.425 99.815 131.410 100.175 ;
        RECT 131.880 100.005 132.115 100.655 ;
        RECT 129.165 98.955 129.335 99.565 ;
        RECT 129.505 99.175 129.835 99.610 ;
        RECT 130.075 99.125 130.315 99.645 ;
        RECT 131.240 99.480 131.410 99.815 ;
        RECT 131.580 99.675 132.115 100.005 ;
        RECT 131.895 99.525 132.115 99.675 ;
        RECT 132.285 99.635 132.585 100.485 ;
        RECT 133.275 100.340 133.565 101.505 ;
        RECT 134.285 100.835 134.455 101.335 ;
        RECT 134.625 101.005 134.955 101.505 ;
        RECT 134.285 100.665 134.950 100.835 ;
        RECT 134.200 99.845 134.550 100.495 ;
        RECT 130.485 98.955 130.880 99.450 ;
        RECT 131.240 99.285 131.615 99.480 ;
        RECT 131.445 99.140 131.615 99.285 ;
        RECT 131.895 99.150 132.135 99.525 ;
        RECT 132.305 98.955 132.640 99.460 ;
        RECT 133.275 98.955 133.565 99.680 ;
        RECT 134.720 99.675 134.950 100.665 ;
        RECT 134.285 99.505 134.950 99.675 ;
        RECT 134.285 99.215 134.455 99.505 ;
        RECT 134.625 98.955 134.955 99.335 ;
        RECT 135.125 99.215 135.310 101.335 ;
        RECT 135.550 101.045 135.815 101.505 ;
        RECT 135.985 100.910 136.235 101.335 ;
        RECT 136.445 101.060 137.550 101.230 ;
        RECT 135.930 100.780 136.235 100.910 ;
        RECT 135.480 99.585 135.760 100.535 ;
        RECT 135.930 99.675 136.100 100.780 ;
        RECT 136.270 99.995 136.510 100.590 ;
        RECT 136.680 100.525 137.210 100.890 ;
        RECT 136.680 99.825 136.850 100.525 ;
        RECT 137.380 100.445 137.550 101.060 ;
        RECT 137.720 100.705 137.890 101.505 ;
        RECT 138.060 101.005 138.310 101.335 ;
        RECT 138.535 101.035 139.420 101.205 ;
        RECT 137.380 100.355 137.890 100.445 ;
        RECT 135.930 99.545 136.155 99.675 ;
        RECT 136.325 99.605 136.850 99.825 ;
        RECT 137.020 100.185 137.890 100.355 ;
        RECT 135.565 98.955 135.815 99.415 ;
        RECT 135.985 99.405 136.155 99.545 ;
        RECT 137.020 99.405 137.190 100.185 ;
        RECT 137.720 100.115 137.890 100.185 ;
        RECT 137.400 99.935 137.600 99.965 ;
        RECT 138.060 99.935 138.230 101.005 ;
        RECT 138.400 100.115 138.590 100.835 ;
        RECT 137.400 99.635 138.230 99.935 ;
        RECT 138.760 99.905 139.080 100.865 ;
        RECT 135.985 99.235 136.320 99.405 ;
        RECT 136.515 99.235 137.190 99.405 ;
        RECT 137.510 98.955 137.880 99.455 ;
        RECT 138.060 99.405 138.230 99.635 ;
        RECT 138.615 99.575 139.080 99.905 ;
        RECT 139.250 100.195 139.420 101.035 ;
        RECT 139.600 101.005 139.915 101.505 ;
        RECT 140.145 100.775 140.485 101.335 ;
        RECT 139.590 100.400 140.485 100.775 ;
        RECT 140.655 100.495 140.825 101.505 ;
        RECT 140.295 100.195 140.485 100.400 ;
        RECT 140.995 100.445 141.325 101.290 ;
        RECT 140.995 100.365 141.385 100.445 ;
        RECT 141.170 100.315 141.385 100.365 ;
        RECT 139.250 99.865 140.125 100.195 ;
        RECT 140.295 99.865 141.045 100.195 ;
        RECT 139.250 99.405 139.420 99.865 ;
        RECT 140.295 99.695 140.495 99.865 ;
        RECT 141.215 99.735 141.385 100.315 ;
        RECT 141.160 99.695 141.385 99.735 ;
        RECT 138.060 99.235 138.465 99.405 ;
        RECT 138.635 99.235 139.420 99.405 ;
        RECT 139.695 98.955 139.905 99.485 ;
        RECT 140.165 99.170 140.495 99.695 ;
        RECT 141.005 99.610 141.385 99.695 ;
        RECT 141.560 100.365 141.895 101.335 ;
        RECT 142.065 100.365 142.235 101.505 ;
        RECT 142.405 101.165 144.435 101.335 ;
        RECT 141.560 99.695 141.730 100.365 ;
        RECT 142.405 100.195 142.575 101.165 ;
        RECT 141.900 99.865 142.155 100.195 ;
        RECT 142.380 99.865 142.575 100.195 ;
        RECT 142.745 100.825 143.870 100.995 ;
        RECT 141.985 99.695 142.155 99.865 ;
        RECT 142.745 99.695 142.915 100.825 ;
        RECT 140.665 98.955 140.835 99.565 ;
        RECT 141.005 99.175 141.335 99.610 ;
        RECT 141.560 99.125 141.815 99.695 ;
        RECT 141.985 99.525 142.915 99.695 ;
        RECT 143.085 100.485 144.095 100.655 ;
        RECT 143.085 99.685 143.255 100.485 ;
        RECT 143.460 99.805 143.735 100.285 ;
        RECT 143.455 99.635 143.735 99.805 ;
        RECT 142.740 99.490 142.915 99.525 ;
        RECT 141.985 98.955 142.315 99.355 ;
        RECT 142.740 99.125 143.270 99.490 ;
        RECT 143.460 99.125 143.735 99.635 ;
        RECT 143.905 99.125 144.095 100.485 ;
        RECT 144.265 100.500 144.435 101.165 ;
        RECT 144.605 100.745 144.775 101.505 ;
        RECT 145.010 100.745 145.525 101.155 ;
        RECT 144.265 100.310 145.015 100.500 ;
        RECT 145.185 99.935 145.525 100.745 ;
        RECT 144.295 99.765 145.525 99.935 ;
        RECT 145.695 100.415 146.905 101.505 ;
        RECT 145.695 99.875 146.215 100.415 ;
        RECT 144.275 98.955 144.785 99.490 ;
        RECT 145.005 99.160 145.250 99.765 ;
        RECT 146.385 99.705 146.905 100.245 ;
        RECT 145.695 98.955 146.905 99.705 ;
        RECT 17.270 98.785 146.990 98.955 ;
        RECT 17.355 98.035 18.565 98.785 ;
        RECT 19.245 98.130 19.575 98.565 ;
        RECT 19.745 98.175 19.915 98.785 ;
        RECT 19.195 98.045 19.575 98.130 ;
        RECT 20.085 98.045 20.415 98.570 ;
        RECT 20.675 98.255 20.885 98.785 ;
        RECT 21.160 98.335 21.945 98.505 ;
        RECT 22.115 98.335 22.520 98.505 ;
        RECT 17.355 97.495 17.875 98.035 ;
        RECT 19.195 98.005 19.420 98.045 ;
        RECT 18.045 97.325 18.565 97.865 ;
        RECT 17.355 96.235 18.565 97.325 ;
        RECT 19.195 97.425 19.365 98.005 ;
        RECT 20.085 97.875 20.285 98.045 ;
        RECT 21.160 97.875 21.330 98.335 ;
        RECT 19.535 97.545 20.285 97.875 ;
        RECT 20.455 97.545 21.330 97.875 ;
        RECT 19.195 97.375 19.410 97.425 ;
        RECT 19.195 97.295 19.585 97.375 ;
        RECT 19.255 96.450 19.585 97.295 ;
        RECT 20.095 97.340 20.285 97.545 ;
        RECT 19.755 96.235 19.925 97.245 ;
        RECT 20.095 96.965 20.990 97.340 ;
        RECT 20.095 96.405 20.435 96.965 ;
        RECT 20.665 96.235 20.980 96.735 ;
        RECT 21.160 96.705 21.330 97.545 ;
        RECT 21.500 97.835 21.965 98.165 ;
        RECT 22.350 98.105 22.520 98.335 ;
        RECT 22.700 98.285 23.070 98.785 ;
        RECT 23.390 98.335 24.065 98.505 ;
        RECT 24.260 98.335 24.595 98.505 ;
        RECT 21.500 96.875 21.820 97.835 ;
        RECT 22.350 97.805 23.180 98.105 ;
        RECT 21.990 96.905 22.180 97.625 ;
        RECT 22.350 96.735 22.520 97.805 ;
        RECT 22.980 97.775 23.180 97.805 ;
        RECT 22.690 97.555 22.860 97.625 ;
        RECT 23.390 97.555 23.560 98.335 ;
        RECT 24.425 98.195 24.595 98.335 ;
        RECT 24.765 98.325 25.015 98.785 ;
        RECT 22.690 97.385 23.560 97.555 ;
        RECT 23.730 97.915 24.255 98.135 ;
        RECT 24.425 98.065 24.650 98.195 ;
        RECT 22.690 97.295 23.200 97.385 ;
        RECT 21.160 96.535 22.045 96.705 ;
        RECT 22.270 96.405 22.520 96.735 ;
        RECT 22.690 96.235 22.860 97.035 ;
        RECT 23.030 96.680 23.200 97.295 ;
        RECT 23.730 97.215 23.900 97.915 ;
        RECT 23.370 96.850 23.900 97.215 ;
        RECT 24.070 97.150 24.310 97.745 ;
        RECT 24.480 96.960 24.650 98.065 ;
        RECT 24.820 97.205 25.100 98.155 ;
        RECT 24.345 96.830 24.650 96.960 ;
        RECT 23.030 96.510 24.135 96.680 ;
        RECT 24.345 96.405 24.595 96.830 ;
        RECT 24.765 96.235 25.030 96.695 ;
        RECT 25.270 96.405 25.455 98.525 ;
        RECT 25.625 98.405 25.955 98.785 ;
        RECT 26.125 98.235 26.295 98.525 ;
        RECT 25.630 98.065 26.295 98.235 ;
        RECT 25.630 97.075 25.860 98.065 ;
        RECT 26.560 98.045 26.815 98.615 ;
        RECT 26.985 98.385 27.315 98.785 ;
        RECT 27.740 98.250 28.270 98.615 ;
        RECT 28.460 98.445 28.735 98.615 ;
        RECT 28.455 98.275 28.735 98.445 ;
        RECT 27.740 98.215 27.915 98.250 ;
        RECT 26.985 98.045 27.915 98.215 ;
        RECT 26.030 97.245 26.380 97.895 ;
        RECT 26.560 97.375 26.730 98.045 ;
        RECT 26.985 97.875 27.155 98.045 ;
        RECT 26.900 97.545 27.155 97.875 ;
        RECT 27.380 97.545 27.575 97.875 ;
        RECT 25.630 96.905 26.295 97.075 ;
        RECT 25.625 96.235 25.955 96.735 ;
        RECT 26.125 96.405 26.295 96.905 ;
        RECT 26.560 96.405 26.895 97.375 ;
        RECT 27.065 96.235 27.235 97.375 ;
        RECT 27.405 96.575 27.575 97.545 ;
        RECT 27.745 96.915 27.915 98.045 ;
        RECT 28.085 97.255 28.255 98.055 ;
        RECT 28.460 97.455 28.735 98.275 ;
        RECT 28.905 97.255 29.095 98.615 ;
        RECT 29.275 98.250 29.785 98.785 ;
        RECT 30.005 97.975 30.250 98.580 ;
        RECT 31.625 98.060 31.955 98.570 ;
        RECT 32.125 98.385 32.455 98.785 ;
        RECT 33.505 98.215 33.835 98.555 ;
        RECT 34.005 98.385 34.335 98.785 ;
        RECT 29.295 97.805 30.525 97.975 ;
        RECT 28.085 97.085 29.095 97.255 ;
        RECT 29.265 97.240 30.015 97.430 ;
        RECT 27.745 96.745 28.870 96.915 ;
        RECT 29.265 96.575 29.435 97.240 ;
        RECT 30.185 96.995 30.525 97.805 ;
        RECT 27.405 96.405 29.435 96.575 ;
        RECT 29.605 96.235 29.775 96.995 ;
        RECT 30.010 96.585 30.525 96.995 ;
        RECT 31.625 97.295 31.815 98.060 ;
        RECT 32.125 98.045 34.490 98.215 ;
        RECT 32.125 97.875 32.295 98.045 ;
        RECT 31.985 97.545 32.295 97.875 ;
        RECT 32.465 97.545 32.770 97.875 ;
        RECT 31.625 96.445 31.955 97.295 ;
        RECT 32.125 96.235 32.375 97.375 ;
        RECT 32.555 97.215 32.770 97.545 ;
        RECT 32.945 97.215 33.230 97.875 ;
        RECT 33.425 97.215 33.690 97.875 ;
        RECT 33.905 97.215 34.150 97.875 ;
        RECT 34.320 97.045 34.490 98.045 ;
        RECT 32.565 96.875 33.855 97.045 ;
        RECT 32.565 96.455 32.815 96.875 ;
        RECT 33.045 96.235 33.375 96.705 ;
        RECT 33.605 96.455 33.855 96.875 ;
        RECT 34.035 96.875 34.490 97.045 ;
        RECT 34.835 98.045 35.195 98.420 ;
        RECT 35.460 98.045 35.630 98.785 ;
        RECT 35.910 98.215 36.080 98.420 ;
        RECT 35.910 98.045 36.450 98.215 ;
        RECT 34.835 97.390 35.090 98.045 ;
        RECT 35.260 97.545 35.610 97.875 ;
        RECT 35.780 97.545 36.110 97.875 ;
        RECT 34.035 96.445 34.365 96.875 ;
        RECT 34.835 96.405 35.175 97.390 ;
        RECT 35.345 97.005 35.610 97.545 ;
        RECT 36.280 97.345 36.450 98.045 ;
        RECT 35.825 97.175 36.450 97.345 ;
        RECT 36.620 97.415 36.790 98.615 ;
        RECT 37.020 98.135 37.350 98.615 ;
        RECT 37.520 98.315 37.690 98.785 ;
        RECT 37.860 98.135 38.190 98.600 ;
        RECT 37.020 97.965 38.190 98.135 ;
        RECT 38.515 98.110 38.785 98.455 ;
        RECT 38.975 98.385 39.355 98.785 ;
        RECT 39.525 98.215 39.695 98.565 ;
        RECT 39.865 98.385 40.195 98.785 ;
        RECT 40.395 98.215 40.565 98.565 ;
        RECT 40.765 98.285 41.095 98.785 ;
        RECT 36.960 97.585 37.530 97.795 ;
        RECT 37.700 97.585 38.345 97.795 ;
        RECT 36.620 97.005 37.325 97.415 ;
        RECT 38.515 97.375 38.685 98.110 ;
        RECT 38.955 98.045 40.565 98.215 ;
        RECT 38.955 97.875 39.125 98.045 ;
        RECT 38.855 97.545 39.125 97.875 ;
        RECT 39.295 97.545 39.700 97.875 ;
        RECT 38.955 97.375 39.125 97.545 ;
        RECT 35.345 96.835 37.325 97.005 ;
        RECT 35.345 96.235 35.755 96.665 ;
        RECT 36.500 96.235 36.830 96.655 ;
        RECT 37.000 96.405 37.325 96.835 ;
        RECT 37.800 96.235 38.130 97.335 ;
        RECT 38.515 96.405 38.785 97.375 ;
        RECT 38.955 97.205 39.680 97.375 ;
        RECT 39.870 97.255 40.580 97.875 ;
        RECT 40.750 97.545 41.100 98.115 ;
        RECT 41.295 97.975 41.535 98.785 ;
        RECT 41.705 97.975 42.035 98.615 ;
        RECT 42.205 97.975 42.475 98.785 ;
        RECT 43.115 98.060 43.405 98.785 ;
        RECT 41.275 97.545 41.625 97.795 ;
        RECT 41.795 97.375 41.965 97.975 ;
        RECT 43.575 97.840 43.915 98.615 ;
        RECT 44.085 98.325 44.255 98.785 ;
        RECT 44.495 98.350 44.855 98.615 ;
        RECT 44.495 98.345 44.850 98.350 ;
        RECT 44.495 98.335 44.845 98.345 ;
        RECT 44.495 98.330 44.840 98.335 ;
        RECT 44.495 98.320 44.835 98.330 ;
        RECT 45.485 98.325 45.655 98.785 ;
        RECT 44.495 98.315 44.830 98.320 ;
        RECT 44.495 98.305 44.820 98.315 ;
        RECT 44.495 98.295 44.810 98.305 ;
        RECT 44.495 98.155 44.795 98.295 ;
        RECT 44.085 97.965 44.795 98.155 ;
        RECT 44.985 98.155 45.315 98.235 ;
        RECT 45.825 98.155 46.165 98.615 ;
        RECT 46.335 98.240 51.680 98.785 ;
        RECT 51.855 98.240 57.200 98.785 ;
        RECT 44.985 97.965 46.165 98.155 ;
        RECT 42.135 97.545 42.485 97.795 ;
        RECT 39.510 97.085 39.680 97.205 ;
        RECT 40.780 97.085 41.100 97.375 ;
        RECT 38.995 96.235 39.275 97.035 ;
        RECT 39.510 96.915 41.100 97.085 ;
        RECT 41.285 97.205 41.965 97.375 ;
        RECT 39.445 96.455 41.100 96.745 ;
        RECT 41.285 96.420 41.615 97.205 ;
        RECT 42.145 96.235 42.475 97.375 ;
        RECT 43.115 96.235 43.405 97.400 ;
        RECT 43.575 96.405 43.855 97.840 ;
        RECT 44.085 97.395 44.370 97.965 ;
        RECT 44.555 97.565 45.025 97.795 ;
        RECT 45.195 97.775 45.525 97.795 ;
        RECT 45.195 97.595 45.645 97.775 ;
        RECT 45.835 97.595 46.165 97.795 ;
        RECT 44.085 97.180 45.235 97.395 ;
        RECT 44.025 96.235 44.735 97.010 ;
        RECT 44.905 96.405 45.235 97.180 ;
        RECT 45.430 96.480 45.645 97.595 ;
        RECT 45.935 97.255 46.165 97.595 ;
        RECT 47.920 97.410 48.260 98.240 ;
        RECT 45.825 96.235 46.155 96.955 ;
        RECT 49.740 96.670 50.090 97.920 ;
        RECT 53.440 97.410 53.780 98.240 ;
        RECT 57.375 98.110 57.635 98.615 ;
        RECT 57.815 98.405 58.145 98.785 ;
        RECT 58.325 98.235 58.495 98.615 ;
        RECT 55.260 96.670 55.610 97.920 ;
        RECT 57.375 97.310 57.545 98.110 ;
        RECT 57.830 98.065 58.495 98.235 ;
        RECT 57.830 97.810 58.000 98.065 ;
        RECT 58.755 98.015 60.425 98.785 ;
        RECT 60.685 98.235 60.855 98.525 ;
        RECT 61.025 98.405 61.355 98.785 ;
        RECT 60.685 98.065 61.350 98.235 ;
        RECT 57.715 97.480 58.000 97.810 ;
        RECT 58.235 97.515 58.565 97.885 ;
        RECT 58.755 97.495 59.505 98.015 ;
        RECT 57.830 97.335 58.000 97.480 ;
        RECT 46.335 96.235 51.680 96.670 ;
        RECT 51.855 96.235 57.200 96.670 ;
        RECT 57.375 96.405 57.645 97.310 ;
        RECT 57.830 97.165 58.495 97.335 ;
        RECT 59.675 97.325 60.425 97.845 ;
        RECT 57.815 96.235 58.145 96.995 ;
        RECT 58.325 96.405 58.495 97.165 ;
        RECT 58.755 96.235 60.425 97.325 ;
        RECT 60.600 97.245 60.950 97.895 ;
        RECT 61.120 97.075 61.350 98.065 ;
        RECT 60.685 96.905 61.350 97.075 ;
        RECT 60.685 96.405 60.855 96.905 ;
        RECT 61.025 96.235 61.355 96.735 ;
        RECT 61.525 96.405 61.710 98.525 ;
        RECT 61.965 98.325 62.215 98.785 ;
        RECT 62.385 98.335 62.720 98.505 ;
        RECT 62.915 98.335 63.590 98.505 ;
        RECT 62.385 98.195 62.555 98.335 ;
        RECT 61.880 97.205 62.160 98.155 ;
        RECT 62.330 98.065 62.555 98.195 ;
        RECT 62.330 96.960 62.500 98.065 ;
        RECT 62.725 97.915 63.250 98.135 ;
        RECT 62.670 97.150 62.910 97.745 ;
        RECT 63.080 97.215 63.250 97.915 ;
        RECT 63.420 97.555 63.590 98.335 ;
        RECT 63.910 98.285 64.280 98.785 ;
        RECT 64.460 98.335 64.865 98.505 ;
        RECT 65.035 98.335 65.820 98.505 ;
        RECT 64.460 98.105 64.630 98.335 ;
        RECT 63.800 97.805 64.630 98.105 ;
        RECT 65.015 97.835 65.480 98.165 ;
        RECT 63.800 97.775 64.000 97.805 ;
        RECT 64.120 97.555 64.290 97.625 ;
        RECT 63.420 97.385 64.290 97.555 ;
        RECT 63.780 97.295 64.290 97.385 ;
        RECT 62.330 96.830 62.635 96.960 ;
        RECT 63.080 96.850 63.610 97.215 ;
        RECT 61.950 96.235 62.215 96.695 ;
        RECT 62.385 96.405 62.635 96.830 ;
        RECT 63.780 96.680 63.950 97.295 ;
        RECT 62.845 96.510 63.950 96.680 ;
        RECT 64.120 96.235 64.290 97.035 ;
        RECT 64.460 96.735 64.630 97.805 ;
        RECT 64.800 96.905 64.990 97.625 ;
        RECT 65.160 96.875 65.480 97.835 ;
        RECT 65.650 97.875 65.820 98.335 ;
        RECT 66.095 98.255 66.305 98.785 ;
        RECT 66.565 98.045 66.895 98.570 ;
        RECT 67.065 98.175 67.235 98.785 ;
        RECT 67.405 98.130 67.735 98.565 ;
        RECT 67.405 98.045 67.785 98.130 ;
        RECT 68.875 98.060 69.165 98.785 ;
        RECT 66.695 97.875 66.895 98.045 ;
        RECT 67.560 98.005 67.785 98.045 ;
        RECT 65.650 97.545 66.525 97.875 ;
        RECT 66.695 97.545 67.445 97.875 ;
        RECT 64.460 96.405 64.710 96.735 ;
        RECT 65.650 96.705 65.820 97.545 ;
        RECT 66.695 97.340 66.885 97.545 ;
        RECT 67.615 97.425 67.785 98.005 ;
        RECT 67.570 97.375 67.785 97.425 ;
        RECT 69.340 98.045 69.595 98.615 ;
        RECT 69.765 98.385 70.095 98.785 ;
        RECT 70.520 98.250 71.050 98.615 ;
        RECT 70.520 98.215 70.695 98.250 ;
        RECT 69.765 98.045 70.695 98.215 ;
        RECT 65.990 96.965 66.885 97.340 ;
        RECT 67.395 97.295 67.785 97.375 ;
        RECT 64.935 96.535 65.820 96.705 ;
        RECT 66.000 96.235 66.315 96.735 ;
        RECT 66.545 96.405 66.885 96.965 ;
        RECT 67.055 96.235 67.225 97.245 ;
        RECT 67.395 96.450 67.725 97.295 ;
        RECT 68.875 96.235 69.165 97.400 ;
        RECT 69.340 97.375 69.510 98.045 ;
        RECT 69.765 97.875 69.935 98.045 ;
        RECT 69.680 97.545 69.935 97.875 ;
        RECT 70.160 97.545 70.355 97.875 ;
        RECT 69.340 96.405 69.675 97.375 ;
        RECT 69.845 96.235 70.015 97.375 ;
        RECT 70.185 96.575 70.355 97.545 ;
        RECT 70.525 96.915 70.695 98.045 ;
        RECT 70.865 97.255 71.035 98.055 ;
        RECT 71.240 97.765 71.515 98.615 ;
        RECT 71.235 97.595 71.515 97.765 ;
        RECT 71.240 97.455 71.515 97.595 ;
        RECT 71.685 97.255 71.875 98.615 ;
        RECT 72.055 98.250 72.565 98.785 ;
        RECT 72.785 97.975 73.030 98.580 ;
        RECT 73.480 98.020 73.935 98.785 ;
        RECT 74.210 98.405 75.510 98.615 ;
        RECT 75.765 98.425 76.095 98.785 ;
        RECT 75.340 98.255 75.510 98.405 ;
        RECT 76.265 98.285 76.525 98.615 ;
        RECT 76.295 98.275 76.525 98.285 ;
        RECT 72.075 97.805 73.305 97.975 ;
        RECT 70.865 97.085 71.875 97.255 ;
        RECT 72.045 97.240 72.795 97.430 ;
        RECT 70.525 96.745 71.650 96.915 ;
        RECT 72.045 96.575 72.215 97.240 ;
        RECT 72.965 96.995 73.305 97.805 ;
        RECT 74.410 97.795 74.630 98.195 ;
        RECT 73.475 97.595 73.965 97.795 ;
        RECT 74.155 97.585 74.630 97.795 ;
        RECT 74.875 97.795 75.085 98.195 ;
        RECT 75.340 98.130 76.095 98.255 ;
        RECT 75.340 98.085 76.185 98.130 ;
        RECT 75.915 97.965 76.185 98.085 ;
        RECT 74.875 97.585 75.205 97.795 ;
        RECT 75.375 97.525 75.785 97.830 ;
        RECT 70.185 96.405 72.215 96.575 ;
        RECT 72.385 96.235 72.555 96.995 ;
        RECT 72.790 96.585 73.305 96.995 ;
        RECT 73.480 97.355 74.655 97.415 ;
        RECT 76.015 97.390 76.185 97.965 ;
        RECT 75.985 97.355 76.185 97.390 ;
        RECT 73.480 97.245 76.185 97.355 ;
        RECT 73.480 96.625 73.735 97.245 ;
        RECT 74.325 97.185 76.125 97.245 ;
        RECT 74.325 97.155 74.655 97.185 ;
        RECT 76.355 97.085 76.525 98.275 ;
        RECT 76.695 98.240 82.040 98.785 ;
        RECT 78.280 97.410 78.620 98.240 ;
        RECT 82.215 98.035 83.425 98.785 ;
        RECT 83.685 98.235 83.855 98.525 ;
        RECT 84.025 98.405 84.355 98.785 ;
        RECT 83.685 98.065 84.350 98.235 ;
        RECT 73.985 96.985 74.170 97.075 ;
        RECT 74.760 96.985 75.595 96.995 ;
        RECT 73.985 96.785 75.595 96.985 ;
        RECT 73.985 96.745 74.215 96.785 ;
        RECT 73.480 96.405 73.815 96.625 ;
        RECT 74.820 96.235 75.175 96.615 ;
        RECT 75.345 96.405 75.595 96.785 ;
        RECT 75.845 96.235 76.095 97.015 ;
        RECT 76.265 96.405 76.525 97.085 ;
        RECT 80.100 96.670 80.450 97.920 ;
        RECT 82.215 97.495 82.735 98.035 ;
        RECT 82.905 97.325 83.425 97.865 ;
        RECT 76.695 96.235 82.040 96.670 ;
        RECT 82.215 96.235 83.425 97.325 ;
        RECT 83.600 97.245 83.950 97.895 ;
        RECT 84.120 97.075 84.350 98.065 ;
        RECT 83.685 96.905 84.350 97.075 ;
        RECT 83.685 96.405 83.855 96.905 ;
        RECT 84.025 96.235 84.355 96.735 ;
        RECT 84.525 96.405 84.710 98.525 ;
        RECT 84.965 98.325 85.215 98.785 ;
        RECT 85.385 98.335 85.720 98.505 ;
        RECT 85.915 98.335 86.590 98.505 ;
        RECT 85.385 98.195 85.555 98.335 ;
        RECT 84.880 97.205 85.160 98.155 ;
        RECT 85.330 98.065 85.555 98.195 ;
        RECT 85.330 96.960 85.500 98.065 ;
        RECT 85.725 97.915 86.250 98.135 ;
        RECT 85.670 97.150 85.910 97.745 ;
        RECT 86.080 97.215 86.250 97.915 ;
        RECT 86.420 97.555 86.590 98.335 ;
        RECT 86.910 98.285 87.280 98.785 ;
        RECT 87.460 98.335 87.865 98.505 ;
        RECT 88.035 98.335 88.820 98.505 ;
        RECT 87.460 98.105 87.630 98.335 ;
        RECT 86.800 97.805 87.630 98.105 ;
        RECT 88.015 97.835 88.480 98.165 ;
        RECT 86.800 97.775 87.000 97.805 ;
        RECT 87.120 97.555 87.290 97.625 ;
        RECT 86.420 97.385 87.290 97.555 ;
        RECT 86.780 97.295 87.290 97.385 ;
        RECT 85.330 96.830 85.635 96.960 ;
        RECT 86.080 96.850 86.610 97.215 ;
        RECT 84.950 96.235 85.215 96.695 ;
        RECT 85.385 96.405 85.635 96.830 ;
        RECT 86.780 96.680 86.950 97.295 ;
        RECT 85.845 96.510 86.950 96.680 ;
        RECT 87.120 96.235 87.290 97.035 ;
        RECT 87.460 96.735 87.630 97.805 ;
        RECT 87.800 96.905 87.990 97.625 ;
        RECT 88.160 96.875 88.480 97.835 ;
        RECT 88.650 97.875 88.820 98.335 ;
        RECT 89.095 98.255 89.305 98.785 ;
        RECT 89.565 98.045 89.895 98.570 ;
        RECT 90.065 98.175 90.235 98.785 ;
        RECT 90.405 98.130 90.735 98.565 ;
        RECT 91.045 98.135 91.215 98.615 ;
        RECT 91.385 98.305 91.715 98.785 ;
        RECT 91.940 98.365 93.475 98.615 ;
        RECT 91.940 98.135 92.110 98.365 ;
        RECT 90.405 98.045 90.785 98.130 ;
        RECT 89.695 97.875 89.895 98.045 ;
        RECT 90.560 98.005 90.785 98.045 ;
        RECT 88.650 97.545 89.525 97.875 ;
        RECT 89.695 97.545 90.445 97.875 ;
        RECT 87.460 96.405 87.710 96.735 ;
        RECT 88.650 96.705 88.820 97.545 ;
        RECT 89.695 97.340 89.885 97.545 ;
        RECT 90.615 97.425 90.785 98.005 ;
        RECT 91.045 97.965 92.110 98.135 ;
        RECT 92.290 97.795 92.570 98.195 ;
        RECT 90.960 97.585 91.310 97.795 ;
        RECT 91.480 97.595 91.925 97.795 ;
        RECT 92.095 97.595 92.570 97.795 ;
        RECT 92.840 97.795 93.125 98.195 ;
        RECT 93.305 98.135 93.475 98.365 ;
        RECT 93.645 98.305 93.975 98.785 ;
        RECT 94.190 98.285 94.445 98.615 ;
        RECT 94.235 98.275 94.445 98.285 ;
        RECT 94.260 98.205 94.445 98.275 ;
        RECT 93.305 97.965 94.105 98.135 ;
        RECT 92.840 97.595 93.170 97.795 ;
        RECT 93.340 97.595 93.705 97.795 ;
        RECT 90.570 97.375 90.785 97.425 ;
        RECT 93.935 97.415 94.105 97.965 ;
        RECT 88.990 96.965 89.885 97.340 ;
        RECT 90.395 97.295 90.785 97.375 ;
        RECT 87.935 96.535 88.820 96.705 ;
        RECT 89.000 96.235 89.315 96.735 ;
        RECT 89.545 96.405 89.885 96.965 ;
        RECT 90.055 96.235 90.225 97.245 ;
        RECT 90.395 96.450 90.725 97.295 ;
        RECT 91.045 97.245 94.105 97.415 ;
        RECT 91.045 96.405 91.215 97.245 ;
        RECT 94.275 97.075 94.445 98.205 ;
        RECT 94.635 98.060 94.925 98.785 ;
        RECT 95.100 98.045 95.355 98.615 ;
        RECT 95.525 98.385 95.855 98.785 ;
        RECT 96.280 98.250 96.810 98.615 ;
        RECT 96.280 98.215 96.455 98.250 ;
        RECT 95.525 98.045 96.455 98.215 ;
        RECT 91.385 96.575 91.715 97.075 ;
        RECT 91.885 96.835 93.520 97.075 ;
        RECT 91.885 96.745 92.115 96.835 ;
        RECT 92.225 96.575 92.555 96.615 ;
        RECT 91.385 96.405 92.555 96.575 ;
        RECT 92.745 96.235 93.100 96.655 ;
        RECT 93.270 96.405 93.520 96.835 ;
        RECT 93.690 96.235 94.020 96.995 ;
        RECT 94.190 96.405 94.445 97.075 ;
        RECT 94.635 96.235 94.925 97.400 ;
        RECT 95.100 97.375 95.270 98.045 ;
        RECT 95.525 97.875 95.695 98.045 ;
        RECT 95.440 97.545 95.695 97.875 ;
        RECT 95.920 97.545 96.115 97.875 ;
        RECT 95.100 96.405 95.435 97.375 ;
        RECT 95.605 96.235 95.775 97.375 ;
        RECT 95.945 96.575 96.115 97.545 ;
        RECT 96.285 96.915 96.455 98.045 ;
        RECT 96.625 97.255 96.795 98.055 ;
        RECT 97.000 97.765 97.275 98.615 ;
        RECT 96.995 97.595 97.275 97.765 ;
        RECT 97.000 97.455 97.275 97.595 ;
        RECT 97.445 97.255 97.635 98.615 ;
        RECT 97.815 98.250 98.325 98.785 ;
        RECT 98.545 97.975 98.790 98.580 ;
        RECT 99.240 98.280 99.575 98.785 ;
        RECT 99.745 98.215 99.985 98.590 ;
        RECT 100.265 98.455 100.435 98.600 ;
        RECT 100.265 98.260 100.640 98.455 ;
        RECT 101.000 98.290 101.395 98.785 ;
        RECT 97.835 97.805 99.065 97.975 ;
        RECT 96.625 97.085 97.635 97.255 ;
        RECT 97.805 97.240 98.555 97.430 ;
        RECT 96.285 96.745 97.410 96.915 ;
        RECT 97.805 96.575 97.975 97.240 ;
        RECT 98.725 96.995 99.065 97.805 ;
        RECT 99.295 97.255 99.595 98.105 ;
        RECT 99.765 98.065 99.985 98.215 ;
        RECT 99.765 97.735 100.300 98.065 ;
        RECT 100.470 97.925 100.640 98.260 ;
        RECT 101.565 98.095 101.805 98.615 ;
        RECT 99.765 97.085 100.000 97.735 ;
        RECT 100.470 97.565 101.455 97.925 ;
        RECT 95.945 96.405 97.975 96.575 ;
        RECT 98.145 96.235 98.315 96.995 ;
        RECT 98.550 96.585 99.065 96.995 ;
        RECT 99.325 96.855 100.000 97.085 ;
        RECT 100.170 97.545 101.455 97.565 ;
        RECT 100.170 97.395 101.030 97.545 ;
        RECT 99.325 96.425 99.495 96.855 ;
        RECT 99.665 96.235 99.995 96.685 ;
        RECT 100.170 96.450 100.455 97.395 ;
        RECT 101.630 97.290 101.805 98.095 ;
        RECT 101.995 98.015 104.585 98.785 ;
        RECT 104.760 98.280 105.095 98.785 ;
        RECT 105.265 98.215 105.505 98.590 ;
        RECT 105.785 98.455 105.955 98.600 ;
        RECT 105.785 98.260 106.160 98.455 ;
        RECT 106.520 98.290 106.915 98.785 ;
        RECT 101.995 97.495 103.205 98.015 ;
        RECT 103.375 97.325 104.585 97.845 ;
        RECT 100.630 96.915 101.325 97.225 ;
        RECT 100.635 96.235 101.320 96.705 ;
        RECT 101.500 96.505 101.805 97.290 ;
        RECT 101.995 96.235 104.585 97.325 ;
        RECT 104.815 97.255 105.115 98.105 ;
        RECT 105.285 98.065 105.505 98.215 ;
        RECT 105.285 97.735 105.820 98.065 ;
        RECT 105.990 97.925 106.160 98.260 ;
        RECT 107.085 98.095 107.325 98.615 ;
        RECT 105.285 97.085 105.520 97.735 ;
        RECT 105.990 97.565 106.975 97.925 ;
        RECT 104.845 96.855 105.520 97.085 ;
        RECT 105.690 97.545 106.975 97.565 ;
        RECT 105.690 97.395 106.550 97.545 ;
        RECT 104.845 96.425 105.015 96.855 ;
        RECT 105.185 96.235 105.515 96.685 ;
        RECT 105.690 96.450 105.975 97.395 ;
        RECT 107.150 97.290 107.325 98.095 ;
        RECT 107.515 98.015 111.025 98.785 ;
        RECT 111.195 98.035 112.405 98.785 ;
        RECT 112.580 98.280 112.915 98.785 ;
        RECT 113.085 98.215 113.325 98.590 ;
        RECT 113.605 98.455 113.775 98.600 ;
        RECT 113.605 98.260 113.980 98.455 ;
        RECT 114.340 98.290 114.735 98.785 ;
        RECT 107.515 97.495 109.165 98.015 ;
        RECT 109.335 97.325 111.025 97.845 ;
        RECT 111.195 97.495 111.715 98.035 ;
        RECT 111.885 97.325 112.405 97.865 ;
        RECT 106.150 96.915 106.845 97.225 ;
        RECT 106.155 96.235 106.840 96.705 ;
        RECT 107.020 96.505 107.325 97.290 ;
        RECT 107.515 96.235 111.025 97.325 ;
        RECT 111.195 96.235 112.405 97.325 ;
        RECT 112.635 97.255 112.935 98.105 ;
        RECT 113.105 98.065 113.325 98.215 ;
        RECT 113.105 97.735 113.640 98.065 ;
        RECT 113.810 97.925 113.980 98.260 ;
        RECT 114.905 98.095 115.145 98.615 ;
        RECT 113.105 97.085 113.340 97.735 ;
        RECT 113.810 97.565 114.795 97.925 ;
        RECT 112.665 96.855 113.340 97.085 ;
        RECT 113.510 97.545 114.795 97.565 ;
        RECT 113.510 97.395 114.370 97.545 ;
        RECT 112.665 96.425 112.835 96.855 ;
        RECT 113.005 96.235 113.335 96.685 ;
        RECT 113.510 96.450 113.795 97.395 ;
        RECT 114.970 97.290 115.145 98.095 ;
        RECT 113.970 96.915 114.665 97.225 ;
        RECT 113.975 96.235 114.660 96.705 ;
        RECT 114.840 96.505 115.145 97.290 ;
        RECT 115.800 98.045 116.055 98.615 ;
        RECT 116.225 98.385 116.555 98.785 ;
        RECT 116.980 98.250 117.510 98.615 ;
        RECT 117.700 98.445 117.975 98.615 ;
        RECT 117.695 98.275 117.975 98.445 ;
        RECT 116.980 98.215 117.155 98.250 ;
        RECT 116.225 98.045 117.155 98.215 ;
        RECT 115.800 97.375 115.970 98.045 ;
        RECT 116.225 97.875 116.395 98.045 ;
        RECT 116.140 97.545 116.395 97.875 ;
        RECT 116.620 97.545 116.815 97.875 ;
        RECT 115.800 96.405 116.135 97.375 ;
        RECT 116.305 96.235 116.475 97.375 ;
        RECT 116.645 96.575 116.815 97.545 ;
        RECT 116.985 96.915 117.155 98.045 ;
        RECT 117.325 97.255 117.495 98.055 ;
        RECT 117.700 97.455 117.975 98.275 ;
        RECT 118.145 97.255 118.335 98.615 ;
        RECT 118.515 98.250 119.025 98.785 ;
        RECT 119.245 97.975 119.490 98.580 ;
        RECT 120.395 98.060 120.685 98.785 ;
        RECT 120.855 98.015 123.445 98.785 ;
        RECT 123.705 98.235 123.875 98.525 ;
        RECT 124.045 98.405 124.375 98.785 ;
        RECT 123.705 98.065 124.370 98.235 ;
        RECT 118.535 97.805 119.765 97.975 ;
        RECT 117.325 97.085 118.335 97.255 ;
        RECT 118.505 97.240 119.255 97.430 ;
        RECT 116.985 96.745 118.110 96.915 ;
        RECT 118.505 96.575 118.675 97.240 ;
        RECT 119.425 96.995 119.765 97.805 ;
        RECT 120.855 97.495 122.065 98.015 ;
        RECT 116.645 96.405 118.675 96.575 ;
        RECT 118.845 96.235 119.015 96.995 ;
        RECT 119.250 96.585 119.765 96.995 ;
        RECT 120.395 96.235 120.685 97.400 ;
        RECT 122.235 97.325 123.445 97.845 ;
        RECT 120.855 96.235 123.445 97.325 ;
        RECT 123.620 97.245 123.970 97.895 ;
        RECT 124.140 97.075 124.370 98.065 ;
        RECT 123.705 96.905 124.370 97.075 ;
        RECT 123.705 96.405 123.875 96.905 ;
        RECT 124.045 96.235 124.375 96.735 ;
        RECT 124.545 96.405 124.730 98.525 ;
        RECT 124.985 98.325 125.235 98.785 ;
        RECT 125.405 98.335 125.740 98.505 ;
        RECT 125.935 98.335 126.610 98.505 ;
        RECT 125.405 98.195 125.575 98.335 ;
        RECT 124.900 97.205 125.180 98.155 ;
        RECT 125.350 98.065 125.575 98.195 ;
        RECT 125.350 96.960 125.520 98.065 ;
        RECT 125.745 97.915 126.270 98.135 ;
        RECT 125.690 97.150 125.930 97.745 ;
        RECT 126.100 97.215 126.270 97.915 ;
        RECT 126.440 97.555 126.610 98.335 ;
        RECT 126.930 98.285 127.300 98.785 ;
        RECT 127.480 98.335 127.885 98.505 ;
        RECT 128.055 98.335 128.840 98.505 ;
        RECT 127.480 98.105 127.650 98.335 ;
        RECT 126.820 97.805 127.650 98.105 ;
        RECT 128.035 97.835 128.500 98.165 ;
        RECT 126.820 97.775 127.020 97.805 ;
        RECT 127.140 97.555 127.310 97.625 ;
        RECT 126.440 97.385 127.310 97.555 ;
        RECT 126.800 97.295 127.310 97.385 ;
        RECT 125.350 96.830 125.655 96.960 ;
        RECT 126.100 96.850 126.630 97.215 ;
        RECT 124.970 96.235 125.235 96.695 ;
        RECT 125.405 96.405 125.655 96.830 ;
        RECT 126.800 96.680 126.970 97.295 ;
        RECT 125.865 96.510 126.970 96.680 ;
        RECT 127.140 96.235 127.310 97.035 ;
        RECT 127.480 96.735 127.650 97.805 ;
        RECT 127.820 96.905 128.010 97.625 ;
        RECT 128.180 96.875 128.500 97.835 ;
        RECT 128.670 97.875 128.840 98.335 ;
        RECT 129.115 98.255 129.325 98.785 ;
        RECT 129.585 98.045 129.915 98.570 ;
        RECT 130.085 98.175 130.255 98.785 ;
        RECT 130.425 98.130 130.755 98.565 ;
        RECT 130.425 98.045 130.805 98.130 ;
        RECT 129.715 97.875 129.915 98.045 ;
        RECT 130.580 98.005 130.805 98.045 ;
        RECT 128.670 97.545 129.545 97.875 ;
        RECT 129.715 97.545 130.465 97.875 ;
        RECT 127.480 96.405 127.730 96.735 ;
        RECT 128.670 96.705 128.840 97.545 ;
        RECT 129.715 97.340 129.905 97.545 ;
        RECT 130.635 97.425 130.805 98.005 ;
        RECT 130.590 97.375 130.805 97.425 ;
        RECT 129.010 96.965 129.905 97.340 ;
        RECT 130.415 97.295 130.805 97.375 ;
        RECT 130.980 98.045 131.235 98.615 ;
        RECT 131.405 98.385 131.735 98.785 ;
        RECT 132.160 98.250 132.690 98.615 ;
        RECT 132.880 98.445 133.155 98.615 ;
        RECT 132.875 98.275 133.155 98.445 ;
        RECT 132.160 98.215 132.335 98.250 ;
        RECT 131.405 98.045 132.335 98.215 ;
        RECT 130.980 97.375 131.150 98.045 ;
        RECT 131.405 97.875 131.575 98.045 ;
        RECT 131.320 97.545 131.575 97.875 ;
        RECT 131.800 97.545 131.995 97.875 ;
        RECT 127.955 96.535 128.840 96.705 ;
        RECT 129.020 96.235 129.335 96.735 ;
        RECT 129.565 96.405 129.905 96.965 ;
        RECT 130.075 96.235 130.245 97.245 ;
        RECT 130.415 96.450 130.745 97.295 ;
        RECT 130.980 96.405 131.315 97.375 ;
        RECT 131.485 96.235 131.655 97.375 ;
        RECT 131.825 96.575 131.995 97.545 ;
        RECT 132.165 96.915 132.335 98.045 ;
        RECT 132.505 97.255 132.675 98.055 ;
        RECT 132.880 97.455 133.155 98.275 ;
        RECT 133.325 97.255 133.515 98.615 ;
        RECT 133.695 98.250 134.205 98.785 ;
        RECT 134.425 97.975 134.670 98.580 ;
        RECT 135.115 98.110 135.375 98.615 ;
        RECT 135.555 98.405 135.885 98.785 ;
        RECT 136.065 98.235 136.235 98.615 ;
        RECT 133.715 97.805 134.945 97.975 ;
        RECT 132.505 97.085 133.515 97.255 ;
        RECT 133.685 97.240 134.435 97.430 ;
        RECT 132.165 96.745 133.290 96.915 ;
        RECT 133.685 96.575 133.855 97.240 ;
        RECT 134.605 96.995 134.945 97.805 ;
        RECT 131.825 96.405 133.855 96.575 ;
        RECT 134.025 96.235 134.195 96.995 ;
        RECT 134.430 96.585 134.945 96.995 ;
        RECT 135.115 97.310 135.295 98.110 ;
        RECT 135.570 98.065 136.235 98.235 ;
        RECT 136.585 98.235 136.755 98.525 ;
        RECT 136.925 98.405 137.255 98.785 ;
        RECT 136.585 98.065 137.250 98.235 ;
        RECT 135.570 97.810 135.740 98.065 ;
        RECT 135.465 97.480 135.740 97.810 ;
        RECT 135.965 97.515 136.305 97.885 ;
        RECT 135.570 97.335 135.740 97.480 ;
        RECT 135.115 96.405 135.385 97.310 ;
        RECT 135.570 97.165 136.245 97.335 ;
        RECT 136.500 97.245 136.850 97.895 ;
        RECT 135.555 96.235 135.885 96.995 ;
        RECT 136.065 96.405 136.245 97.165 ;
        RECT 137.020 97.075 137.250 98.065 ;
        RECT 136.585 96.905 137.250 97.075 ;
        RECT 136.585 96.405 136.755 96.905 ;
        RECT 136.925 96.235 137.255 96.735 ;
        RECT 137.425 96.405 137.610 98.525 ;
        RECT 137.865 98.325 138.115 98.785 ;
        RECT 138.285 98.335 138.620 98.505 ;
        RECT 138.815 98.335 139.490 98.505 ;
        RECT 138.285 98.195 138.455 98.335 ;
        RECT 137.780 97.205 138.060 98.155 ;
        RECT 138.230 98.065 138.455 98.195 ;
        RECT 138.230 96.960 138.400 98.065 ;
        RECT 138.625 97.915 139.150 98.135 ;
        RECT 138.570 97.150 138.810 97.745 ;
        RECT 138.980 97.215 139.150 97.915 ;
        RECT 139.320 97.555 139.490 98.335 ;
        RECT 139.810 98.285 140.180 98.785 ;
        RECT 140.360 98.335 140.765 98.505 ;
        RECT 140.935 98.335 141.720 98.505 ;
        RECT 140.360 98.105 140.530 98.335 ;
        RECT 139.700 97.805 140.530 98.105 ;
        RECT 140.915 97.835 141.380 98.165 ;
        RECT 139.700 97.775 139.900 97.805 ;
        RECT 140.020 97.555 140.190 97.625 ;
        RECT 139.320 97.385 140.190 97.555 ;
        RECT 139.680 97.295 140.190 97.385 ;
        RECT 138.230 96.830 138.535 96.960 ;
        RECT 138.980 96.850 139.510 97.215 ;
        RECT 137.850 96.235 138.115 96.695 ;
        RECT 138.285 96.405 138.535 96.830 ;
        RECT 139.680 96.680 139.850 97.295 ;
        RECT 138.745 96.510 139.850 96.680 ;
        RECT 140.020 96.235 140.190 97.035 ;
        RECT 140.360 96.735 140.530 97.805 ;
        RECT 140.700 96.905 140.890 97.625 ;
        RECT 141.060 96.875 141.380 97.835 ;
        RECT 141.550 97.875 141.720 98.335 ;
        RECT 141.995 98.255 142.205 98.785 ;
        RECT 142.465 98.045 142.795 98.570 ;
        RECT 142.965 98.175 143.135 98.785 ;
        RECT 143.305 98.130 143.635 98.565 ;
        RECT 143.945 98.235 144.115 98.615 ;
        RECT 144.330 98.405 144.660 98.785 ;
        RECT 143.305 98.045 143.685 98.130 ;
        RECT 143.945 98.065 144.660 98.235 ;
        RECT 142.595 97.875 142.795 98.045 ;
        RECT 143.460 98.005 143.685 98.045 ;
        RECT 141.550 97.545 142.425 97.875 ;
        RECT 142.595 97.545 143.345 97.875 ;
        RECT 140.360 96.405 140.610 96.735 ;
        RECT 141.550 96.705 141.720 97.545 ;
        RECT 142.595 97.340 142.785 97.545 ;
        RECT 143.515 97.425 143.685 98.005 ;
        RECT 143.855 97.515 144.210 97.885 ;
        RECT 144.490 97.875 144.660 98.065 ;
        RECT 144.830 98.040 145.085 98.615 ;
        RECT 144.490 97.545 144.745 97.875 ;
        RECT 143.470 97.375 143.685 97.425 ;
        RECT 141.890 96.965 142.785 97.340 ;
        RECT 143.295 97.295 143.685 97.375 ;
        RECT 144.490 97.335 144.660 97.545 ;
        RECT 140.835 96.535 141.720 96.705 ;
        RECT 141.900 96.235 142.215 96.735 ;
        RECT 142.445 96.405 142.785 96.965 ;
        RECT 142.955 96.235 143.125 97.245 ;
        RECT 143.295 96.450 143.625 97.295 ;
        RECT 143.945 97.165 144.660 97.335 ;
        RECT 144.915 97.310 145.085 98.040 ;
        RECT 145.260 97.945 145.520 98.785 ;
        RECT 145.695 98.035 146.905 98.785 ;
        RECT 143.945 96.405 144.115 97.165 ;
        RECT 144.330 96.235 144.660 96.995 ;
        RECT 144.830 96.405 145.085 97.310 ;
        RECT 145.260 96.235 145.520 97.385 ;
        RECT 145.695 97.325 146.215 97.865 ;
        RECT 146.385 97.495 146.905 98.035 ;
        RECT 145.695 96.235 146.905 97.325 ;
        RECT 17.270 96.065 146.990 96.235 ;
        RECT 17.355 94.975 18.565 96.065 ;
        RECT 17.355 94.265 17.875 94.805 ;
        RECT 18.045 94.435 18.565 94.975 ;
        RECT 18.815 95.135 18.995 95.895 ;
        RECT 19.175 95.305 19.505 96.065 ;
        RECT 18.815 94.965 19.490 95.135 ;
        RECT 19.675 94.990 19.945 95.895 ;
        RECT 19.320 94.820 19.490 94.965 ;
        RECT 18.755 94.415 19.095 94.785 ;
        RECT 19.320 94.490 19.595 94.820 ;
        RECT 17.355 93.515 18.565 94.265 ;
        RECT 19.320 94.235 19.490 94.490 ;
        RECT 18.825 94.065 19.490 94.235 ;
        RECT 19.765 94.190 19.945 94.990 ;
        RECT 20.205 95.135 20.375 95.895 ;
        RECT 20.555 95.305 20.885 96.065 ;
        RECT 20.205 94.965 20.870 95.135 ;
        RECT 21.055 94.990 21.325 95.895 ;
        RECT 20.700 94.820 20.870 94.965 ;
        RECT 20.135 94.415 20.465 94.785 ;
        RECT 20.700 94.490 20.985 94.820 ;
        RECT 20.700 94.235 20.870 94.490 ;
        RECT 18.825 93.685 18.995 94.065 ;
        RECT 19.175 93.515 19.505 93.895 ;
        RECT 19.685 93.685 19.945 94.190 ;
        RECT 20.205 94.065 20.870 94.235 ;
        RECT 21.155 94.190 21.325 94.990 ;
        RECT 21.960 94.915 22.220 96.065 ;
        RECT 22.395 94.990 22.650 95.895 ;
        RECT 22.820 95.305 23.150 96.065 ;
        RECT 23.365 95.135 23.535 95.895 ;
        RECT 20.205 93.685 20.375 94.065 ;
        RECT 20.555 93.515 20.885 93.895 ;
        RECT 21.065 93.685 21.325 94.190 ;
        RECT 21.960 93.515 22.220 94.355 ;
        RECT 22.395 94.260 22.565 94.990 ;
        RECT 22.820 94.965 23.535 95.135 ;
        RECT 23.875 95.135 24.055 95.895 ;
        RECT 24.235 95.305 24.565 96.065 ;
        RECT 23.875 94.965 24.550 95.135 ;
        RECT 24.735 94.990 25.005 95.895 ;
        RECT 22.820 94.755 22.990 94.965 ;
        RECT 24.380 94.820 24.550 94.965 ;
        RECT 22.735 94.425 22.990 94.755 ;
        RECT 22.395 93.685 22.650 94.260 ;
        RECT 22.820 94.235 22.990 94.425 ;
        RECT 23.270 94.415 23.625 94.785 ;
        RECT 23.815 94.415 24.155 94.785 ;
        RECT 24.380 94.490 24.655 94.820 ;
        RECT 24.380 94.235 24.550 94.490 ;
        RECT 22.820 94.065 23.535 94.235 ;
        RECT 22.820 93.515 23.150 93.895 ;
        RECT 23.365 93.685 23.535 94.065 ;
        RECT 23.885 94.065 24.550 94.235 ;
        RECT 24.825 94.190 25.005 94.990 ;
        RECT 25.255 95.135 25.435 95.895 ;
        RECT 25.615 95.305 25.945 96.065 ;
        RECT 25.255 94.965 25.930 95.135 ;
        RECT 26.115 94.990 26.385 95.895 ;
        RECT 25.760 94.820 25.930 94.965 ;
        RECT 25.195 94.415 25.535 94.785 ;
        RECT 25.760 94.490 26.035 94.820 ;
        RECT 25.760 94.235 25.930 94.490 ;
        RECT 23.885 93.685 24.055 94.065 ;
        RECT 24.235 93.515 24.565 93.895 ;
        RECT 24.745 93.685 25.005 94.190 ;
        RECT 25.265 94.065 25.930 94.235 ;
        RECT 26.205 94.190 26.385 94.990 ;
        RECT 26.555 94.975 28.225 96.065 ;
        RECT 25.265 93.685 25.435 94.065 ;
        RECT 25.615 93.515 25.945 93.895 ;
        RECT 26.125 93.685 26.385 94.190 ;
        RECT 26.555 94.285 27.305 94.805 ;
        RECT 27.475 94.455 28.225 94.975 ;
        RECT 28.485 95.135 28.655 95.895 ;
        RECT 28.870 95.305 29.200 96.065 ;
        RECT 28.485 94.965 29.200 95.135 ;
        RECT 29.370 94.990 29.625 95.895 ;
        RECT 28.395 94.415 28.750 94.785 ;
        RECT 29.030 94.755 29.200 94.965 ;
        RECT 29.030 94.425 29.285 94.755 ;
        RECT 26.555 93.515 28.225 94.285 ;
        RECT 29.030 94.235 29.200 94.425 ;
        RECT 29.455 94.260 29.625 94.990 ;
        RECT 29.800 94.915 30.060 96.065 ;
        RECT 30.235 94.900 30.525 96.065 ;
        RECT 30.775 95.135 30.955 95.895 ;
        RECT 31.135 95.305 31.465 96.065 ;
        RECT 30.775 94.965 31.450 95.135 ;
        RECT 31.635 94.990 31.905 95.895 ;
        RECT 31.280 94.820 31.450 94.965 ;
        RECT 30.715 94.415 31.055 94.785 ;
        RECT 31.280 94.490 31.555 94.820 ;
        RECT 28.485 94.065 29.200 94.235 ;
        RECT 28.485 93.685 28.655 94.065 ;
        RECT 28.870 93.515 29.200 93.895 ;
        RECT 29.370 93.685 29.625 94.260 ;
        RECT 29.800 93.515 30.060 94.355 ;
        RECT 30.235 93.515 30.525 94.240 ;
        RECT 31.280 94.235 31.450 94.490 ;
        RECT 30.785 94.065 31.450 94.235 ;
        RECT 31.725 94.190 31.905 94.990 ;
        RECT 30.785 93.685 30.955 94.065 ;
        RECT 31.135 93.515 31.465 93.895 ;
        RECT 31.645 93.685 31.905 94.190 ;
        RECT 32.075 95.265 32.515 95.895 ;
        RECT 32.075 94.255 32.385 95.265 ;
        RECT 32.690 95.215 33.005 96.065 ;
        RECT 33.175 95.725 34.605 95.895 ;
        RECT 33.175 95.045 33.345 95.725 ;
        RECT 32.555 94.875 33.345 95.045 ;
        RECT 32.555 94.425 32.725 94.875 ;
        RECT 33.515 94.755 33.715 95.555 ;
        RECT 32.895 94.425 33.285 94.705 ;
        RECT 33.470 94.425 33.715 94.755 ;
        RECT 33.915 94.425 34.165 95.555 ;
        RECT 34.355 95.095 34.605 95.725 ;
        RECT 34.785 95.265 35.115 96.065 ;
        RECT 35.385 95.135 35.555 95.895 ;
        RECT 35.735 95.305 36.065 96.065 ;
        RECT 34.355 94.925 35.125 95.095 ;
        RECT 35.385 94.965 36.050 95.135 ;
        RECT 36.235 94.990 36.505 95.895 ;
        RECT 34.380 94.425 34.785 94.755 ;
        RECT 34.955 94.255 35.125 94.925 ;
        RECT 35.880 94.820 36.050 94.965 ;
        RECT 35.315 94.415 35.645 94.785 ;
        RECT 35.880 94.490 36.165 94.820 ;
        RECT 32.075 93.695 32.515 94.255 ;
        RECT 32.685 93.515 33.135 94.255 ;
        RECT 33.305 94.085 34.465 94.255 ;
        RECT 33.305 93.685 33.475 94.085 ;
        RECT 33.645 93.515 34.065 93.915 ;
        RECT 34.235 93.685 34.465 94.085 ;
        RECT 34.635 93.685 35.125 94.255 ;
        RECT 35.880 94.235 36.050 94.490 ;
        RECT 35.385 94.065 36.050 94.235 ;
        RECT 36.335 94.190 36.505 94.990 ;
        RECT 36.675 94.975 37.885 96.065 ;
        RECT 35.385 93.685 35.555 94.065 ;
        RECT 35.735 93.515 36.065 93.895 ;
        RECT 36.245 93.685 36.505 94.190 ;
        RECT 36.675 94.265 37.195 94.805 ;
        RECT 37.365 94.435 37.885 94.975 ;
        RECT 38.145 95.135 38.315 95.895 ;
        RECT 38.495 95.305 38.825 96.065 ;
        RECT 38.145 94.965 38.810 95.135 ;
        RECT 38.995 94.990 39.265 95.895 ;
        RECT 38.640 94.820 38.810 94.965 ;
        RECT 38.075 94.415 38.405 94.785 ;
        RECT 38.640 94.490 38.925 94.820 ;
        RECT 36.675 93.515 37.885 94.265 ;
        RECT 38.640 94.235 38.810 94.490 ;
        RECT 38.145 94.065 38.810 94.235 ;
        RECT 39.095 94.190 39.265 94.990 ;
        RECT 39.435 94.975 41.105 96.065 ;
        RECT 38.145 93.685 38.315 94.065 ;
        RECT 38.495 93.515 38.825 93.895 ;
        RECT 39.005 93.685 39.265 94.190 ;
        RECT 39.435 94.285 40.185 94.805 ;
        RECT 40.355 94.455 41.105 94.975 ;
        RECT 41.275 94.990 41.545 95.895 ;
        RECT 41.715 95.305 42.045 96.065 ;
        RECT 42.225 95.135 42.405 95.895 ;
        RECT 39.435 93.515 41.105 94.285 ;
        RECT 41.275 94.190 41.455 94.990 ;
        RECT 41.730 94.965 42.405 95.135 ;
        RECT 41.730 94.820 41.900 94.965 ;
        RECT 43.115 94.900 43.405 96.065 ;
        RECT 44.495 94.990 44.765 95.895 ;
        RECT 44.935 95.305 45.265 96.065 ;
        RECT 45.445 95.135 45.625 95.895 ;
        RECT 41.625 94.490 41.900 94.820 ;
        RECT 41.730 94.235 41.900 94.490 ;
        RECT 42.125 94.415 42.465 94.785 ;
        RECT 41.275 93.685 41.535 94.190 ;
        RECT 41.730 94.065 42.395 94.235 ;
        RECT 41.715 93.515 42.045 93.895 ;
        RECT 42.225 93.685 42.395 94.065 ;
        RECT 43.115 93.515 43.405 94.240 ;
        RECT 44.495 94.190 44.675 94.990 ;
        RECT 44.950 94.965 45.625 95.135 ;
        RECT 45.875 94.975 47.545 96.065 ;
        RECT 44.950 94.820 45.120 94.965 ;
        RECT 44.845 94.490 45.120 94.820 ;
        RECT 44.950 94.235 45.120 94.490 ;
        RECT 45.345 94.415 45.685 94.785 ;
        RECT 45.875 94.285 46.625 94.805 ;
        RECT 46.795 94.455 47.545 94.975 ;
        RECT 47.715 94.990 47.985 95.895 ;
        RECT 48.155 95.305 48.485 96.065 ;
        RECT 48.665 95.135 48.845 95.895 ;
        RECT 44.495 93.685 44.755 94.190 ;
        RECT 44.950 94.065 45.615 94.235 ;
        RECT 44.935 93.515 45.265 93.895 ;
        RECT 45.445 93.685 45.615 94.065 ;
        RECT 45.875 93.515 47.545 94.285 ;
        RECT 47.715 94.190 47.895 94.990 ;
        RECT 48.170 94.965 48.845 95.135 ;
        RECT 49.095 94.975 50.765 96.065 ;
        RECT 48.170 94.820 48.340 94.965 ;
        RECT 48.065 94.490 48.340 94.820 ;
        RECT 48.170 94.235 48.340 94.490 ;
        RECT 48.565 94.415 48.905 94.785 ;
        RECT 49.095 94.285 49.845 94.805 ;
        RECT 50.015 94.455 50.765 94.975 ;
        RECT 50.935 94.990 51.205 95.895 ;
        RECT 51.375 95.305 51.705 96.065 ;
        RECT 51.885 95.135 52.055 95.895 ;
        RECT 47.715 93.685 47.975 94.190 ;
        RECT 48.170 94.065 48.835 94.235 ;
        RECT 48.155 93.515 48.485 93.895 ;
        RECT 48.665 93.685 48.835 94.065 ;
        RECT 49.095 93.515 50.765 94.285 ;
        RECT 50.935 94.190 51.105 94.990 ;
        RECT 51.390 94.965 52.055 95.135 ;
        RECT 52.315 94.975 53.985 96.065 ;
        RECT 51.390 94.820 51.560 94.965 ;
        RECT 51.275 94.490 51.560 94.820 ;
        RECT 51.390 94.235 51.560 94.490 ;
        RECT 51.795 94.415 52.125 94.785 ;
        RECT 52.315 94.285 53.065 94.805 ;
        RECT 53.235 94.455 53.985 94.975 ;
        RECT 54.155 94.990 54.425 95.895 ;
        RECT 54.595 95.305 54.925 96.065 ;
        RECT 55.105 95.135 55.275 95.895 ;
        RECT 50.935 93.685 51.195 94.190 ;
        RECT 51.390 94.065 52.055 94.235 ;
        RECT 51.375 93.515 51.705 93.895 ;
        RECT 51.885 93.685 52.055 94.065 ;
        RECT 52.315 93.515 53.985 94.285 ;
        RECT 54.155 94.190 54.325 94.990 ;
        RECT 54.610 94.965 55.275 95.135 ;
        RECT 54.610 94.820 54.780 94.965 ;
        RECT 55.995 94.900 56.285 96.065 ;
        RECT 56.460 94.915 56.720 96.065 ;
        RECT 56.895 94.990 57.150 95.895 ;
        RECT 57.320 95.305 57.650 96.065 ;
        RECT 57.865 95.135 58.035 95.895 ;
        RECT 54.495 94.490 54.780 94.820 ;
        RECT 54.610 94.235 54.780 94.490 ;
        RECT 55.015 94.415 55.345 94.785 ;
        RECT 54.155 93.685 54.415 94.190 ;
        RECT 54.610 94.065 55.275 94.235 ;
        RECT 54.595 93.515 54.925 93.895 ;
        RECT 55.105 93.685 55.275 94.065 ;
        RECT 55.995 93.515 56.285 94.240 ;
        RECT 56.460 93.515 56.720 94.355 ;
        RECT 56.895 94.260 57.065 94.990 ;
        RECT 57.320 94.965 58.035 95.135 ;
        RECT 57.320 94.755 57.490 94.965 ;
        RECT 58.300 94.915 58.560 96.065 ;
        RECT 58.735 94.990 58.990 95.895 ;
        RECT 59.160 95.305 59.490 96.065 ;
        RECT 59.705 95.135 59.875 95.895 ;
        RECT 57.235 94.425 57.490 94.755 ;
        RECT 56.895 93.685 57.150 94.260 ;
        RECT 57.320 94.235 57.490 94.425 ;
        RECT 57.770 94.415 58.125 94.785 ;
        RECT 57.320 94.065 58.035 94.235 ;
        RECT 57.320 93.515 57.650 93.895 ;
        RECT 57.865 93.685 58.035 94.065 ;
        RECT 58.300 93.515 58.560 94.355 ;
        RECT 58.735 94.260 58.905 94.990 ;
        RECT 59.160 94.965 59.875 95.135 ;
        RECT 59.160 94.755 59.330 94.965 ;
        RECT 60.140 94.915 60.400 96.065 ;
        RECT 60.575 94.990 60.830 95.895 ;
        RECT 61.000 95.305 61.330 96.065 ;
        RECT 61.545 95.135 61.715 95.895 ;
        RECT 59.075 94.425 59.330 94.755 ;
        RECT 58.735 93.685 58.990 94.260 ;
        RECT 59.160 94.235 59.330 94.425 ;
        RECT 59.610 94.415 59.965 94.785 ;
        RECT 59.160 94.065 59.875 94.235 ;
        RECT 59.160 93.515 59.490 93.895 ;
        RECT 59.705 93.685 59.875 94.065 ;
        RECT 60.140 93.515 60.400 94.355 ;
        RECT 60.575 94.260 60.745 94.990 ;
        RECT 61.000 94.965 61.715 95.135 ;
        RECT 61.995 95.010 62.300 95.795 ;
        RECT 62.480 95.595 63.165 96.065 ;
        RECT 62.475 95.075 63.170 95.385 ;
        RECT 61.000 94.755 61.170 94.965 ;
        RECT 60.915 94.425 61.170 94.755 ;
        RECT 60.575 93.685 60.830 94.260 ;
        RECT 61.000 94.235 61.170 94.425 ;
        RECT 61.450 94.415 61.805 94.785 ;
        RECT 61.000 94.065 61.715 94.235 ;
        RECT 61.000 93.515 61.330 93.895 ;
        RECT 61.545 93.685 61.715 94.065 ;
        RECT 61.995 94.205 62.170 95.010 ;
        RECT 63.345 94.905 63.630 95.850 ;
        RECT 63.805 95.615 64.135 96.065 ;
        RECT 64.305 95.445 64.475 95.875 ;
        RECT 62.770 94.755 63.630 94.905 ;
        RECT 62.345 94.735 63.630 94.755 ;
        RECT 63.800 95.215 64.475 95.445 ;
        RECT 65.745 95.445 65.915 95.875 ;
        RECT 66.085 95.615 66.415 96.065 ;
        RECT 65.745 95.215 66.420 95.445 ;
        RECT 62.345 94.375 63.330 94.735 ;
        RECT 63.800 94.565 64.035 95.215 ;
        RECT 61.995 93.685 62.235 94.205 ;
        RECT 63.160 94.040 63.330 94.375 ;
        RECT 63.500 94.235 64.035 94.565 ;
        RECT 63.815 94.085 64.035 94.235 ;
        RECT 64.205 94.195 64.505 95.045 ;
        RECT 65.715 94.195 66.015 95.045 ;
        RECT 66.185 94.565 66.420 95.215 ;
        RECT 66.590 94.905 66.875 95.850 ;
        RECT 67.055 95.595 67.740 96.065 ;
        RECT 67.050 95.075 67.745 95.385 ;
        RECT 67.920 95.010 68.225 95.795 ;
        RECT 66.590 94.755 67.450 94.905 ;
        RECT 66.590 94.735 67.875 94.755 ;
        RECT 66.185 94.235 66.720 94.565 ;
        RECT 66.890 94.375 67.875 94.735 ;
        RECT 66.185 94.085 66.405 94.235 ;
        RECT 62.405 93.515 62.800 94.010 ;
        RECT 63.160 93.845 63.535 94.040 ;
        RECT 63.365 93.700 63.535 93.845 ;
        RECT 63.815 93.710 64.055 94.085 ;
        RECT 64.225 93.515 64.560 94.020 ;
        RECT 65.660 93.515 65.995 94.020 ;
        RECT 66.165 93.710 66.405 94.085 ;
        RECT 66.890 94.040 67.060 94.375 ;
        RECT 68.050 94.205 68.225 95.010 ;
        RECT 68.875 94.900 69.165 96.065 ;
        RECT 69.340 94.925 69.675 95.895 ;
        RECT 69.845 94.925 70.015 96.065 ;
        RECT 70.185 95.725 72.215 95.895 ;
        RECT 69.340 94.255 69.510 94.925 ;
        RECT 70.185 94.755 70.355 95.725 ;
        RECT 69.680 94.425 69.935 94.755 ;
        RECT 70.160 94.425 70.355 94.755 ;
        RECT 70.525 95.385 71.650 95.555 ;
        RECT 69.765 94.255 69.935 94.425 ;
        RECT 70.525 94.255 70.695 95.385 ;
        RECT 66.685 93.845 67.060 94.040 ;
        RECT 66.685 93.700 66.855 93.845 ;
        RECT 67.420 93.515 67.815 94.010 ;
        RECT 67.985 93.685 68.225 94.205 ;
        RECT 68.875 93.515 69.165 94.240 ;
        RECT 69.340 93.685 69.595 94.255 ;
        RECT 69.765 94.085 70.695 94.255 ;
        RECT 70.865 95.045 71.875 95.215 ;
        RECT 70.865 94.245 71.035 95.045 ;
        RECT 71.240 94.705 71.515 94.845 ;
        RECT 71.235 94.535 71.515 94.705 ;
        RECT 70.520 94.050 70.695 94.085 ;
        RECT 69.765 93.515 70.095 93.915 ;
        RECT 70.520 93.685 71.050 94.050 ;
        RECT 71.240 93.685 71.515 94.535 ;
        RECT 71.685 93.685 71.875 95.045 ;
        RECT 72.045 95.060 72.215 95.725 ;
        RECT 72.385 95.305 72.555 96.065 ;
        RECT 72.790 95.305 73.305 95.715 ;
        RECT 72.045 94.870 72.795 95.060 ;
        RECT 72.965 94.495 73.305 95.305 ;
        RECT 73.565 95.135 73.735 95.895 ;
        RECT 73.950 95.305 74.280 96.065 ;
        RECT 73.565 94.965 74.280 95.135 ;
        RECT 74.450 94.990 74.705 95.895 ;
        RECT 72.075 94.325 73.305 94.495 ;
        RECT 73.475 94.415 73.830 94.785 ;
        RECT 74.110 94.755 74.280 94.965 ;
        RECT 74.110 94.425 74.365 94.755 ;
        RECT 72.055 93.515 72.565 94.050 ;
        RECT 72.785 93.720 73.030 94.325 ;
        RECT 74.110 94.235 74.280 94.425 ;
        RECT 74.535 94.260 74.705 94.990 ;
        RECT 74.880 94.915 75.140 96.065 ;
        RECT 76.240 94.915 76.500 96.065 ;
        RECT 76.675 94.990 76.930 95.895 ;
        RECT 77.100 95.305 77.430 96.065 ;
        RECT 77.645 95.135 77.815 95.895 ;
        RECT 73.565 94.065 74.280 94.235 ;
        RECT 73.565 93.685 73.735 94.065 ;
        RECT 73.950 93.515 74.280 93.895 ;
        RECT 74.450 93.685 74.705 94.260 ;
        RECT 74.880 93.515 75.140 94.355 ;
        RECT 76.240 93.515 76.500 94.355 ;
        RECT 76.675 94.260 76.845 94.990 ;
        RECT 77.100 94.965 77.815 95.135 ;
        RECT 78.165 95.135 78.335 95.895 ;
        RECT 78.550 95.305 78.880 96.065 ;
        RECT 78.165 94.965 78.880 95.135 ;
        RECT 79.050 94.990 79.305 95.895 ;
        RECT 77.100 94.755 77.270 94.965 ;
        RECT 77.015 94.425 77.270 94.755 ;
        RECT 76.675 93.685 76.930 94.260 ;
        RECT 77.100 94.235 77.270 94.425 ;
        RECT 77.550 94.415 77.905 94.785 ;
        RECT 78.075 94.415 78.430 94.785 ;
        RECT 78.710 94.755 78.880 94.965 ;
        RECT 78.710 94.425 78.965 94.755 ;
        RECT 78.710 94.235 78.880 94.425 ;
        RECT 79.135 94.260 79.305 94.990 ;
        RECT 79.480 94.915 79.740 96.065 ;
        RECT 80.005 95.135 80.175 95.895 ;
        RECT 80.390 95.305 80.720 96.065 ;
        RECT 80.005 94.965 80.720 95.135 ;
        RECT 80.890 94.990 81.145 95.895 ;
        RECT 79.915 94.415 80.270 94.785 ;
        RECT 80.550 94.755 80.720 94.965 ;
        RECT 80.550 94.425 80.805 94.755 ;
        RECT 77.100 94.065 77.815 94.235 ;
        RECT 77.100 93.515 77.430 93.895 ;
        RECT 77.645 93.685 77.815 94.065 ;
        RECT 78.165 94.065 78.880 94.235 ;
        RECT 78.165 93.685 78.335 94.065 ;
        RECT 78.550 93.515 78.880 93.895 ;
        RECT 79.050 93.685 79.305 94.260 ;
        RECT 79.480 93.515 79.740 94.355 ;
        RECT 80.550 94.235 80.720 94.425 ;
        RECT 80.975 94.260 81.145 94.990 ;
        RECT 81.320 94.915 81.580 96.065 ;
        RECT 81.755 94.900 82.045 96.065 ;
        RECT 82.215 94.975 83.425 96.065 ;
        RECT 83.685 95.445 83.855 95.875 ;
        RECT 84.025 95.615 84.355 96.065 ;
        RECT 83.685 95.215 84.360 95.445 ;
        RECT 80.005 94.065 80.720 94.235 ;
        RECT 80.005 93.685 80.175 94.065 ;
        RECT 80.390 93.515 80.720 93.895 ;
        RECT 80.890 93.685 81.145 94.260 ;
        RECT 81.320 93.515 81.580 94.355 ;
        RECT 82.215 94.265 82.735 94.805 ;
        RECT 82.905 94.435 83.425 94.975 ;
        RECT 81.755 93.515 82.045 94.240 ;
        RECT 82.215 93.515 83.425 94.265 ;
        RECT 83.655 94.195 83.955 95.045 ;
        RECT 84.125 94.565 84.360 95.215 ;
        RECT 84.530 94.905 84.815 95.850 ;
        RECT 84.995 95.595 85.680 96.065 ;
        RECT 84.990 95.075 85.685 95.385 ;
        RECT 85.860 95.010 86.165 95.795 ;
        RECT 87.365 95.445 87.535 95.875 ;
        RECT 87.705 95.615 88.035 96.065 ;
        RECT 87.365 95.215 88.040 95.445 ;
        RECT 84.530 94.755 85.390 94.905 ;
        RECT 84.530 94.735 85.815 94.755 ;
        RECT 84.125 94.235 84.660 94.565 ;
        RECT 84.830 94.375 85.815 94.735 ;
        RECT 84.125 94.085 84.345 94.235 ;
        RECT 83.600 93.515 83.935 94.020 ;
        RECT 84.105 93.710 84.345 94.085 ;
        RECT 84.830 94.040 85.000 94.375 ;
        RECT 85.990 94.205 86.165 95.010 ;
        RECT 84.625 93.845 85.000 94.040 ;
        RECT 84.625 93.700 84.795 93.845 ;
        RECT 85.360 93.515 85.755 94.010 ;
        RECT 85.925 93.685 86.165 94.205 ;
        RECT 87.335 94.195 87.635 95.045 ;
        RECT 87.805 94.565 88.040 95.215 ;
        RECT 88.210 94.905 88.495 95.850 ;
        RECT 88.675 95.595 89.360 96.065 ;
        RECT 88.670 95.075 89.365 95.385 ;
        RECT 89.540 95.010 89.845 95.795 ;
        RECT 88.210 94.755 89.070 94.905 ;
        RECT 88.210 94.735 89.495 94.755 ;
        RECT 87.805 94.235 88.340 94.565 ;
        RECT 88.510 94.375 89.495 94.735 ;
        RECT 87.805 94.085 88.025 94.235 ;
        RECT 87.280 93.515 87.615 94.020 ;
        RECT 87.785 93.710 88.025 94.085 ;
        RECT 88.510 94.040 88.680 94.375 ;
        RECT 89.670 94.205 89.845 95.010 ;
        RECT 90.040 94.915 90.300 96.065 ;
        RECT 90.475 94.990 90.730 95.895 ;
        RECT 90.900 95.305 91.230 96.065 ;
        RECT 91.445 95.135 91.615 95.895 ;
        RECT 88.305 93.845 88.680 94.040 ;
        RECT 88.305 93.700 88.475 93.845 ;
        RECT 89.040 93.515 89.435 94.010 ;
        RECT 89.605 93.685 89.845 94.205 ;
        RECT 90.040 93.515 90.300 94.355 ;
        RECT 90.475 94.260 90.645 94.990 ;
        RECT 90.900 94.965 91.615 95.135 ;
        RECT 91.965 95.135 92.135 95.895 ;
        RECT 92.350 95.305 92.680 96.065 ;
        RECT 91.965 94.965 92.680 95.135 ;
        RECT 92.850 94.990 93.105 95.895 ;
        RECT 90.900 94.755 91.070 94.965 ;
        RECT 90.815 94.425 91.070 94.755 ;
        RECT 90.475 93.685 90.730 94.260 ;
        RECT 90.900 94.235 91.070 94.425 ;
        RECT 91.350 94.415 91.705 94.785 ;
        RECT 91.875 94.415 92.230 94.785 ;
        RECT 92.510 94.755 92.680 94.965 ;
        RECT 92.510 94.425 92.765 94.755 ;
        RECT 92.510 94.235 92.680 94.425 ;
        RECT 92.935 94.260 93.105 94.990 ;
        RECT 93.280 94.915 93.540 96.065 ;
        RECT 94.635 94.900 94.925 96.065 ;
        RECT 95.185 95.135 95.355 95.895 ;
        RECT 95.570 95.305 95.900 96.065 ;
        RECT 95.185 94.965 95.900 95.135 ;
        RECT 96.070 94.990 96.325 95.895 ;
        RECT 95.095 94.415 95.450 94.785 ;
        RECT 95.730 94.755 95.900 94.965 ;
        RECT 95.730 94.425 95.985 94.755 ;
        RECT 90.900 94.065 91.615 94.235 ;
        RECT 90.900 93.515 91.230 93.895 ;
        RECT 91.445 93.685 91.615 94.065 ;
        RECT 91.965 94.065 92.680 94.235 ;
        RECT 91.965 93.685 92.135 94.065 ;
        RECT 92.350 93.515 92.680 93.895 ;
        RECT 92.850 93.685 93.105 94.260 ;
        RECT 93.280 93.515 93.540 94.355 ;
        RECT 94.635 93.515 94.925 94.240 ;
        RECT 95.730 94.235 95.900 94.425 ;
        RECT 96.155 94.260 96.325 94.990 ;
        RECT 96.500 94.915 96.760 96.065 ;
        RECT 97.025 95.135 97.195 95.895 ;
        RECT 97.410 95.305 97.740 96.065 ;
        RECT 97.025 94.965 97.740 95.135 ;
        RECT 97.910 94.990 98.165 95.895 ;
        RECT 96.935 94.415 97.290 94.785 ;
        RECT 97.570 94.755 97.740 94.965 ;
        RECT 97.570 94.425 97.825 94.755 ;
        RECT 95.185 94.065 95.900 94.235 ;
        RECT 95.185 93.685 95.355 94.065 ;
        RECT 95.570 93.515 95.900 93.895 ;
        RECT 96.070 93.685 96.325 94.260 ;
        RECT 96.500 93.515 96.760 94.355 ;
        RECT 97.570 94.235 97.740 94.425 ;
        RECT 97.995 94.260 98.165 94.990 ;
        RECT 98.340 94.915 98.600 96.065 ;
        RECT 99.240 94.915 99.500 96.065 ;
        RECT 99.675 94.990 99.930 95.895 ;
        RECT 100.100 95.305 100.430 96.065 ;
        RECT 100.645 95.135 100.815 95.895 ;
        RECT 97.025 94.065 97.740 94.235 ;
        RECT 97.025 93.685 97.195 94.065 ;
        RECT 97.410 93.515 97.740 93.895 ;
        RECT 97.910 93.685 98.165 94.260 ;
        RECT 98.340 93.515 98.600 94.355 ;
        RECT 99.240 93.515 99.500 94.355 ;
        RECT 99.675 94.260 99.845 94.990 ;
        RECT 100.100 94.965 100.815 95.135 ;
        RECT 101.075 94.975 102.285 96.065 ;
        RECT 100.100 94.755 100.270 94.965 ;
        RECT 100.015 94.425 100.270 94.755 ;
        RECT 99.675 93.685 99.930 94.260 ;
        RECT 100.100 94.235 100.270 94.425 ;
        RECT 100.550 94.415 100.905 94.785 ;
        RECT 101.075 94.265 101.595 94.805 ;
        RECT 101.765 94.435 102.285 94.975 ;
        RECT 102.460 94.915 102.720 96.065 ;
        RECT 102.895 94.990 103.150 95.895 ;
        RECT 103.320 95.305 103.650 96.065 ;
        RECT 103.865 95.135 104.035 95.895 ;
        RECT 100.100 94.065 100.815 94.235 ;
        RECT 100.100 93.515 100.430 93.895 ;
        RECT 100.645 93.685 100.815 94.065 ;
        RECT 101.075 93.515 102.285 94.265 ;
        RECT 102.460 93.515 102.720 94.355 ;
        RECT 102.895 94.260 103.065 94.990 ;
        RECT 103.320 94.965 104.035 95.135 ;
        RECT 104.295 94.975 105.505 96.065 ;
        RECT 103.320 94.755 103.490 94.965 ;
        RECT 103.235 94.425 103.490 94.755 ;
        RECT 102.895 93.685 103.150 94.260 ;
        RECT 103.320 94.235 103.490 94.425 ;
        RECT 103.770 94.415 104.125 94.785 ;
        RECT 104.295 94.265 104.815 94.805 ;
        RECT 104.985 94.435 105.505 94.975 ;
        RECT 105.680 94.915 105.940 96.065 ;
        RECT 106.115 94.990 106.370 95.895 ;
        RECT 106.540 95.305 106.870 96.065 ;
        RECT 107.085 95.135 107.255 95.895 ;
        RECT 103.320 94.065 104.035 94.235 ;
        RECT 103.320 93.515 103.650 93.895 ;
        RECT 103.865 93.685 104.035 94.065 ;
        RECT 104.295 93.515 105.505 94.265 ;
        RECT 105.680 93.515 105.940 94.355 ;
        RECT 106.115 94.260 106.285 94.990 ;
        RECT 106.540 94.965 107.255 95.135 ;
        RECT 106.540 94.755 106.710 94.965 ;
        RECT 107.515 94.900 107.805 96.065 ;
        RECT 108.900 94.915 109.160 96.065 ;
        RECT 109.335 94.990 109.590 95.895 ;
        RECT 109.760 95.305 110.090 96.065 ;
        RECT 110.305 95.135 110.475 95.895 ;
        RECT 106.455 94.425 106.710 94.755 ;
        RECT 106.115 93.685 106.370 94.260 ;
        RECT 106.540 94.235 106.710 94.425 ;
        RECT 106.990 94.415 107.345 94.785 ;
        RECT 106.540 94.065 107.255 94.235 ;
        RECT 106.540 93.515 106.870 93.895 ;
        RECT 107.085 93.685 107.255 94.065 ;
        RECT 107.515 93.515 107.805 94.240 ;
        RECT 108.900 93.515 109.160 94.355 ;
        RECT 109.335 94.260 109.505 94.990 ;
        RECT 109.760 94.965 110.475 95.135 ;
        RECT 110.735 94.975 111.945 96.065 ;
        RECT 109.760 94.755 109.930 94.965 ;
        RECT 109.675 94.425 109.930 94.755 ;
        RECT 109.335 93.685 109.590 94.260 ;
        RECT 109.760 94.235 109.930 94.425 ;
        RECT 110.210 94.415 110.565 94.785 ;
        RECT 110.735 94.265 111.255 94.805 ;
        RECT 111.425 94.435 111.945 94.975 ;
        RECT 112.120 94.915 112.380 96.065 ;
        RECT 112.555 94.990 112.810 95.895 ;
        RECT 112.980 95.305 113.310 96.065 ;
        RECT 113.525 95.135 113.695 95.895 ;
        RECT 114.045 95.445 114.215 95.875 ;
        RECT 114.385 95.615 114.715 96.065 ;
        RECT 114.045 95.215 114.720 95.445 ;
        RECT 109.760 94.065 110.475 94.235 ;
        RECT 109.760 93.515 110.090 93.895 ;
        RECT 110.305 93.685 110.475 94.065 ;
        RECT 110.735 93.515 111.945 94.265 ;
        RECT 112.120 93.515 112.380 94.355 ;
        RECT 112.555 94.260 112.725 94.990 ;
        RECT 112.980 94.965 113.695 95.135 ;
        RECT 112.980 94.755 113.150 94.965 ;
        RECT 112.895 94.425 113.150 94.755 ;
        RECT 112.555 93.685 112.810 94.260 ;
        RECT 112.980 94.235 113.150 94.425 ;
        RECT 113.430 94.415 113.785 94.785 ;
        RECT 112.980 94.065 113.695 94.235 ;
        RECT 114.015 94.195 114.315 95.045 ;
        RECT 114.485 94.565 114.720 95.215 ;
        RECT 114.890 94.905 115.175 95.850 ;
        RECT 115.355 95.595 116.040 96.065 ;
        RECT 115.350 95.075 116.045 95.385 ;
        RECT 116.220 95.010 116.525 95.795 ;
        RECT 114.890 94.755 115.750 94.905 ;
        RECT 114.890 94.735 116.175 94.755 ;
        RECT 114.485 94.235 115.020 94.565 ;
        RECT 115.190 94.375 116.175 94.735 ;
        RECT 114.485 94.085 114.705 94.235 ;
        RECT 112.980 93.515 113.310 93.895 ;
        RECT 113.525 93.685 113.695 94.065 ;
        RECT 113.960 93.515 114.295 94.020 ;
        RECT 114.465 93.710 114.705 94.085 ;
        RECT 115.190 94.040 115.360 94.375 ;
        RECT 116.350 94.205 116.525 95.010 ;
        RECT 114.985 93.845 115.360 94.040 ;
        RECT 114.985 93.700 115.155 93.845 ;
        RECT 115.720 93.515 116.115 94.010 ;
        RECT 116.285 93.685 116.525 94.205 ;
        RECT 117.175 95.215 117.435 95.895 ;
        RECT 117.605 95.285 117.855 96.065 ;
        RECT 118.105 95.515 118.355 95.895 ;
        RECT 118.525 95.685 118.880 96.065 ;
        RECT 119.885 95.675 120.220 95.895 ;
        RECT 119.485 95.515 119.715 95.555 ;
        RECT 118.105 95.315 119.715 95.515 ;
        RECT 118.105 95.305 118.940 95.315 ;
        RECT 119.530 95.225 119.715 95.315 ;
        RECT 117.175 94.015 117.345 95.215 ;
        RECT 119.045 95.115 119.375 95.145 ;
        RECT 117.575 95.055 119.375 95.115 ;
        RECT 119.965 95.055 120.220 95.675 ;
        RECT 117.515 94.945 120.220 95.055 ;
        RECT 117.515 94.910 117.715 94.945 ;
        RECT 117.515 94.335 117.685 94.910 ;
        RECT 119.045 94.885 120.220 94.945 ;
        RECT 120.395 94.900 120.685 96.065 ;
        RECT 120.945 95.135 121.115 95.895 ;
        RECT 121.330 95.305 121.660 96.065 ;
        RECT 120.945 94.965 121.660 95.135 ;
        RECT 121.830 94.990 122.085 95.895 ;
        RECT 117.915 94.470 118.325 94.775 ;
        RECT 118.495 94.505 118.825 94.715 ;
        RECT 117.515 94.215 117.785 94.335 ;
        RECT 117.515 94.170 118.360 94.215 ;
        RECT 117.605 94.045 118.360 94.170 ;
        RECT 118.615 94.105 118.825 94.505 ;
        RECT 119.070 94.505 119.545 94.715 ;
        RECT 119.735 94.505 120.225 94.705 ;
        RECT 119.070 94.105 119.290 94.505 ;
        RECT 120.855 94.415 121.210 94.785 ;
        RECT 121.490 94.755 121.660 94.965 ;
        RECT 121.490 94.425 121.745 94.755 ;
        RECT 117.175 93.685 117.435 94.015 ;
        RECT 118.190 93.895 118.360 94.045 ;
        RECT 117.605 93.515 117.935 93.875 ;
        RECT 118.190 93.685 119.490 93.895 ;
        RECT 119.765 93.515 120.220 94.280 ;
        RECT 120.395 93.515 120.685 94.240 ;
        RECT 121.490 94.235 121.660 94.425 ;
        RECT 121.915 94.260 122.085 94.990 ;
        RECT 122.260 94.915 122.520 96.065 ;
        RECT 122.785 95.135 122.955 95.895 ;
        RECT 123.170 95.305 123.500 96.065 ;
        RECT 122.785 94.965 123.500 95.135 ;
        RECT 123.670 94.990 123.925 95.895 ;
        RECT 122.695 94.415 123.050 94.785 ;
        RECT 123.330 94.755 123.500 94.965 ;
        RECT 123.330 94.425 123.585 94.755 ;
        RECT 120.945 94.065 121.660 94.235 ;
        RECT 120.945 93.685 121.115 94.065 ;
        RECT 121.330 93.515 121.660 93.895 ;
        RECT 121.830 93.685 122.085 94.260 ;
        RECT 122.260 93.515 122.520 94.355 ;
        RECT 123.330 94.235 123.500 94.425 ;
        RECT 123.755 94.260 123.925 94.990 ;
        RECT 124.100 94.915 124.360 96.065 ;
        RECT 124.540 94.915 124.800 96.065 ;
        RECT 124.975 94.990 125.230 95.895 ;
        RECT 125.400 95.305 125.730 96.065 ;
        RECT 125.945 95.135 126.115 95.895 ;
        RECT 122.785 94.065 123.500 94.235 ;
        RECT 122.785 93.685 122.955 94.065 ;
        RECT 123.170 93.515 123.500 93.895 ;
        RECT 123.670 93.685 123.925 94.260 ;
        RECT 124.100 93.515 124.360 94.355 ;
        RECT 124.540 93.515 124.800 94.355 ;
        RECT 124.975 94.260 125.145 94.990 ;
        RECT 125.400 94.965 126.115 95.135 ;
        RECT 126.375 95.305 126.890 95.715 ;
        RECT 127.125 95.305 127.295 96.065 ;
        RECT 127.465 95.725 129.495 95.895 ;
        RECT 125.400 94.755 125.570 94.965 ;
        RECT 125.315 94.425 125.570 94.755 ;
        RECT 124.975 93.685 125.230 94.260 ;
        RECT 125.400 94.235 125.570 94.425 ;
        RECT 125.850 94.415 126.205 94.785 ;
        RECT 126.375 94.495 126.715 95.305 ;
        RECT 127.465 95.060 127.635 95.725 ;
        RECT 128.030 95.385 129.155 95.555 ;
        RECT 126.885 94.870 127.635 95.060 ;
        RECT 127.805 95.045 128.815 95.215 ;
        RECT 126.375 94.325 127.605 94.495 ;
        RECT 125.400 94.065 126.115 94.235 ;
        RECT 125.400 93.515 125.730 93.895 ;
        RECT 125.945 93.685 126.115 94.065 ;
        RECT 126.650 93.720 126.895 94.325 ;
        RECT 127.115 93.515 127.625 94.050 ;
        RECT 127.805 93.685 127.995 95.045 ;
        RECT 128.165 94.025 128.440 94.845 ;
        RECT 128.645 94.245 128.815 95.045 ;
        RECT 128.985 94.255 129.155 95.385 ;
        RECT 129.325 94.755 129.495 95.725 ;
        RECT 129.665 94.925 129.835 96.065 ;
        RECT 130.005 94.925 130.340 95.895 ;
        RECT 130.605 95.135 130.775 95.895 ;
        RECT 130.990 95.305 131.320 96.065 ;
        RECT 130.605 94.965 131.320 95.135 ;
        RECT 131.490 94.990 131.745 95.895 ;
        RECT 129.325 94.425 129.520 94.755 ;
        RECT 129.745 94.425 130.000 94.755 ;
        RECT 129.745 94.255 129.915 94.425 ;
        RECT 130.170 94.255 130.340 94.925 ;
        RECT 130.515 94.415 130.870 94.785 ;
        RECT 131.150 94.755 131.320 94.965 ;
        RECT 131.150 94.425 131.405 94.755 ;
        RECT 128.985 94.085 129.915 94.255 ;
        RECT 128.985 94.050 129.160 94.085 ;
        RECT 128.165 93.855 128.445 94.025 ;
        RECT 128.165 93.685 128.440 93.855 ;
        RECT 128.630 93.685 129.160 94.050 ;
        RECT 129.585 93.515 129.915 93.915 ;
        RECT 130.085 93.685 130.340 94.255 ;
        RECT 131.150 94.235 131.320 94.425 ;
        RECT 131.575 94.260 131.745 94.990 ;
        RECT 131.920 94.915 132.180 96.065 ;
        RECT 133.275 94.900 133.565 96.065 ;
        RECT 133.755 95.225 134.010 95.895 ;
        RECT 134.180 95.305 134.510 96.065 ;
        RECT 134.680 95.465 134.930 95.895 ;
        RECT 135.100 95.645 135.455 96.065 ;
        RECT 135.645 95.725 136.815 95.895 ;
        RECT 135.645 95.685 135.975 95.725 ;
        RECT 136.085 95.465 136.315 95.555 ;
        RECT 134.680 95.225 136.315 95.465 ;
        RECT 136.485 95.225 136.815 95.725 ;
        RECT 130.605 94.065 131.320 94.235 ;
        RECT 130.605 93.685 130.775 94.065 ;
        RECT 130.990 93.515 131.320 93.895 ;
        RECT 131.490 93.685 131.745 94.260 ;
        RECT 131.920 93.515 132.180 94.355 ;
        RECT 133.275 93.515 133.565 94.240 ;
        RECT 133.755 94.095 133.925 95.225 ;
        RECT 136.985 95.055 137.155 95.895 ;
        RECT 137.505 95.445 137.675 95.875 ;
        RECT 137.845 95.615 138.175 96.065 ;
        RECT 137.505 95.215 138.180 95.445 ;
        RECT 134.095 94.885 137.155 95.055 ;
        RECT 134.095 94.335 134.265 94.885 ;
        RECT 134.485 94.535 134.860 94.705 ;
        RECT 134.495 94.505 134.860 94.535 ;
        RECT 135.030 94.505 135.360 94.705 ;
        RECT 134.095 94.165 134.895 94.335 ;
        RECT 133.755 94.015 133.940 94.095 ;
        RECT 133.755 93.685 134.010 94.015 ;
        RECT 134.225 93.515 134.555 93.995 ;
        RECT 134.725 93.935 134.895 94.165 ;
        RECT 135.075 94.105 135.360 94.505 ;
        RECT 135.630 94.505 136.105 94.705 ;
        RECT 136.275 94.505 136.720 94.705 ;
        RECT 136.890 94.505 137.240 94.715 ;
        RECT 135.630 94.105 135.910 94.505 ;
        RECT 136.090 94.165 137.155 94.335 ;
        RECT 137.475 94.195 137.775 95.045 ;
        RECT 137.945 94.565 138.180 95.215 ;
        RECT 138.350 94.905 138.635 95.850 ;
        RECT 138.815 95.595 139.500 96.065 ;
        RECT 138.810 95.075 139.505 95.385 ;
        RECT 139.680 95.010 139.985 95.795 ;
        RECT 138.350 94.755 139.210 94.905 ;
        RECT 138.350 94.735 139.635 94.755 ;
        RECT 137.945 94.235 138.480 94.565 ;
        RECT 138.650 94.375 139.635 94.735 ;
        RECT 136.090 93.935 136.260 94.165 ;
        RECT 134.725 93.685 136.260 93.935 ;
        RECT 136.485 93.515 136.815 93.995 ;
        RECT 136.985 93.685 137.155 94.165 ;
        RECT 137.945 94.085 138.165 94.235 ;
        RECT 137.420 93.515 137.755 94.020 ;
        RECT 137.925 93.710 138.165 94.085 ;
        RECT 138.650 94.040 138.820 94.375 ;
        RECT 139.810 94.205 139.985 95.010 ;
        RECT 140.265 95.135 140.435 95.895 ;
        RECT 140.650 95.305 140.980 96.065 ;
        RECT 140.265 94.965 140.980 95.135 ;
        RECT 141.150 94.990 141.405 95.895 ;
        RECT 140.175 94.415 140.530 94.785 ;
        RECT 140.810 94.755 140.980 94.965 ;
        RECT 140.810 94.425 141.065 94.755 ;
        RECT 140.810 94.235 140.980 94.425 ;
        RECT 141.235 94.260 141.405 94.990 ;
        RECT 141.580 94.915 141.840 96.065 ;
        RECT 142.105 95.135 142.275 95.895 ;
        RECT 142.490 95.305 142.820 96.065 ;
        RECT 142.105 94.965 142.820 95.135 ;
        RECT 142.990 94.990 143.245 95.895 ;
        RECT 142.015 94.415 142.370 94.785 ;
        RECT 142.650 94.755 142.820 94.965 ;
        RECT 142.650 94.425 142.905 94.755 ;
        RECT 138.445 93.845 138.820 94.040 ;
        RECT 138.445 93.700 138.615 93.845 ;
        RECT 139.180 93.515 139.575 94.010 ;
        RECT 139.745 93.685 139.985 94.205 ;
        RECT 140.265 94.065 140.980 94.235 ;
        RECT 140.265 93.685 140.435 94.065 ;
        RECT 140.650 93.515 140.980 93.895 ;
        RECT 141.150 93.685 141.405 94.260 ;
        RECT 141.580 93.515 141.840 94.355 ;
        RECT 142.650 94.235 142.820 94.425 ;
        RECT 143.075 94.260 143.245 94.990 ;
        RECT 143.420 94.915 143.680 96.065 ;
        RECT 143.945 95.135 144.115 95.895 ;
        RECT 144.330 95.305 144.660 96.065 ;
        RECT 143.945 94.965 144.660 95.135 ;
        RECT 144.830 94.990 145.085 95.895 ;
        RECT 143.855 94.415 144.210 94.785 ;
        RECT 144.490 94.755 144.660 94.965 ;
        RECT 144.490 94.425 144.745 94.755 ;
        RECT 142.105 94.065 142.820 94.235 ;
        RECT 142.105 93.685 142.275 94.065 ;
        RECT 142.490 93.515 142.820 93.895 ;
        RECT 142.990 93.685 143.245 94.260 ;
        RECT 143.420 93.515 143.680 94.355 ;
        RECT 144.490 94.235 144.660 94.425 ;
        RECT 144.915 94.260 145.085 94.990 ;
        RECT 145.260 94.915 145.520 96.065 ;
        RECT 145.695 94.975 146.905 96.065 ;
        RECT 145.695 94.435 146.215 94.975 ;
        RECT 143.945 94.065 144.660 94.235 ;
        RECT 143.945 93.685 144.115 94.065 ;
        RECT 144.330 93.515 144.660 93.895 ;
        RECT 144.830 93.685 145.085 94.260 ;
        RECT 145.260 93.515 145.520 94.355 ;
        RECT 146.385 94.265 146.905 94.805 ;
        RECT 145.695 93.515 146.905 94.265 ;
        RECT 17.270 93.345 146.990 93.515 ;
        RECT 87.250 76.480 90.620 76.490 ;
        RECT 75.120 76.460 90.620 76.480 ;
        RECT 102.030 76.460 105.400 76.480 ;
        RECT 75.120 76.420 117.910 76.460 ;
        RECT 120.120 76.420 147.910 76.460 ;
        RECT 75.120 76.350 147.910 76.420 ;
        RECT 73.070 76.160 74.720 76.330 ;
        RECT 54.720 75.350 67.430 75.960 ;
        RECT 54.670 75.150 67.480 75.350 ;
        RECT 54.670 68.040 54.840 75.150 ;
        RECT 55.240 68.770 55.410 74.810 ;
        RECT 55.680 68.770 55.850 74.810 ;
        RECT 55.380 68.385 55.710 68.555 ;
        RECT 56.250 68.040 56.420 75.150 ;
        RECT 56.820 68.770 56.990 74.810 ;
        RECT 57.260 68.770 57.430 74.810 ;
        RECT 56.960 68.385 57.290 68.555 ;
        RECT 57.830 68.040 58.000 75.150 ;
        RECT 58.400 68.770 58.570 74.810 ;
        RECT 58.840 68.770 59.010 74.810 ;
        RECT 58.540 68.385 58.870 68.555 ;
        RECT 59.410 68.040 59.580 75.150 ;
        RECT 59.980 68.770 60.150 74.810 ;
        RECT 60.420 68.770 60.590 74.810 ;
        RECT 60.120 68.385 60.450 68.555 ;
        RECT 60.990 68.040 61.160 75.150 ;
        RECT 61.560 68.770 61.730 74.810 ;
        RECT 62.000 68.770 62.170 74.810 ;
        RECT 61.700 68.385 62.030 68.555 ;
        RECT 62.570 68.040 62.740 75.150 ;
        RECT 63.140 68.770 63.310 74.810 ;
        RECT 63.580 68.770 63.750 74.810 ;
        RECT 63.280 68.385 63.610 68.555 ;
        RECT 64.150 68.040 64.320 75.150 ;
        RECT 64.720 68.770 64.890 74.810 ;
        RECT 65.160 68.770 65.330 74.810 ;
        RECT 64.860 68.385 65.190 68.555 ;
        RECT 65.730 68.040 65.900 75.150 ;
        RECT 66.300 68.770 66.470 74.810 ;
        RECT 66.740 68.770 66.910 74.810 ;
        RECT 66.440 68.385 66.770 68.555 ;
        RECT 67.310 68.040 67.480 75.150 ;
        RECT 54.670 67.870 67.480 68.040 ;
        RECT 73.070 70.340 73.240 76.160 ;
        RECT 73.720 73.520 74.070 75.680 ;
        RECT 73.720 70.820 74.070 72.980 ;
        RECT 74.550 70.760 74.720 76.160 ;
        RECT 75.120 75.680 147.920 76.350 ;
        RECT 75.080 75.570 147.920 75.680 ;
        RECT 75.080 75.510 87.930 75.570 ;
        RECT 74.550 70.340 74.730 70.760 ;
        RECT 73.070 70.170 74.730 70.340 ;
        RECT 54.680 66.630 67.490 66.800 ;
        RECT 54.680 63.560 54.850 66.630 ;
        RECT 55.390 66.120 55.720 66.290 ;
        RECT 55.250 63.910 55.420 65.950 ;
        RECT 55.690 63.910 55.860 65.950 ;
        RECT 56.260 63.560 56.430 66.630 ;
        RECT 56.970 66.120 57.300 66.290 ;
        RECT 56.830 63.910 57.000 65.950 ;
        RECT 57.270 63.910 57.440 65.950 ;
        RECT 57.840 63.560 58.010 66.630 ;
        RECT 58.550 66.120 58.880 66.290 ;
        RECT 58.410 63.910 58.580 65.950 ;
        RECT 58.850 63.910 59.020 65.950 ;
        RECT 59.420 63.560 59.590 66.630 ;
        RECT 60.130 66.120 60.460 66.290 ;
        RECT 59.990 63.910 60.160 65.950 ;
        RECT 60.430 63.910 60.600 65.950 ;
        RECT 61.000 63.560 61.170 66.630 ;
        RECT 61.710 66.120 62.040 66.290 ;
        RECT 61.570 63.910 61.740 65.950 ;
        RECT 62.010 63.910 62.180 65.950 ;
        RECT 62.580 63.560 62.750 66.630 ;
        RECT 63.290 66.120 63.620 66.290 ;
        RECT 63.150 63.910 63.320 65.950 ;
        RECT 63.590 63.910 63.760 65.950 ;
        RECT 64.160 63.560 64.330 66.630 ;
        RECT 64.870 66.120 65.200 66.290 ;
        RECT 64.730 63.910 64.900 65.950 ;
        RECT 65.170 63.910 65.340 65.950 ;
        RECT 65.740 63.560 65.910 66.630 ;
        RECT 66.450 66.120 66.780 66.290 ;
        RECT 66.310 63.910 66.480 65.950 ;
        RECT 66.750 63.910 66.920 65.950 ;
        RECT 67.320 63.560 67.490 66.630 ;
        RECT 54.680 63.370 67.490 63.560 ;
        RECT 73.070 64.350 73.240 70.170 ;
        RECT 74.550 69.710 74.730 70.170 ;
        RECT 73.720 67.530 74.070 69.690 ;
        RECT 73.720 64.830 74.070 66.990 ;
        RECT 74.550 64.350 74.720 69.710 ;
        RECT 75.080 66.020 75.250 75.510 ;
        RECT 75.880 75.000 76.880 75.170 ;
        RECT 75.650 66.745 75.820 74.785 ;
        RECT 76.940 66.745 77.110 74.785 ;
        RECT 75.880 66.360 76.880 66.530 ;
        RECT 77.510 66.020 77.680 75.510 ;
        RECT 78.310 75.000 80.310 75.170 ;
        RECT 78.080 66.745 78.250 74.785 ;
        RECT 80.370 66.745 80.540 74.785 ;
        RECT 78.310 66.360 80.310 66.530 ;
        RECT 80.940 66.020 81.110 75.510 ;
        RECT 81.740 75.000 83.740 75.170 ;
        RECT 81.510 66.745 81.680 74.785 ;
        RECT 83.800 66.745 83.970 74.785 ;
        RECT 81.740 66.360 83.740 66.530 ;
        RECT 84.370 66.020 84.540 75.510 ;
        RECT 85.170 75.000 86.170 75.170 ;
        RECT 84.940 66.745 85.110 74.785 ;
        RECT 86.230 66.745 86.400 74.785 ;
        RECT 86.800 69.910 87.930 75.510 ;
        RECT 90.060 75.560 147.920 75.570 ;
        RECT 90.060 75.490 102.910 75.560 ;
        RECT 85.170 66.360 86.170 66.530 ;
        RECT 86.800 66.020 87.950 69.910 ;
        RECT 75.080 65.850 87.950 66.020 ;
        RECT 86.830 65.820 87.950 65.850 ;
        RECT 90.060 66.000 90.230 75.490 ;
        RECT 90.860 74.980 91.860 75.150 ;
        RECT 90.630 66.725 90.800 74.765 ;
        RECT 91.920 66.725 92.090 74.765 ;
        RECT 90.860 66.340 91.860 66.510 ;
        RECT 92.490 66.000 92.660 75.490 ;
        RECT 93.290 74.980 95.290 75.150 ;
        RECT 93.060 66.725 93.230 74.765 ;
        RECT 95.350 66.725 95.520 74.765 ;
        RECT 93.290 66.340 95.290 66.510 ;
        RECT 95.920 66.000 96.090 75.490 ;
        RECT 96.720 74.980 98.720 75.150 ;
        RECT 96.490 66.725 96.660 74.765 ;
        RECT 98.780 66.725 98.950 74.765 ;
        RECT 96.720 66.340 98.720 66.510 ;
        RECT 99.350 66.000 99.520 75.490 ;
        RECT 100.150 74.980 101.150 75.150 ;
        RECT 99.920 66.725 100.090 74.765 ;
        RECT 101.210 66.725 101.380 74.765 ;
        RECT 101.780 69.890 102.910 75.490 ;
        RECT 105.070 75.540 147.920 75.560 ;
        RECT 105.070 75.500 132.930 75.540 ;
        RECT 105.070 75.490 117.920 75.500 ;
        RECT 100.150 66.340 101.150 66.510 ;
        RECT 101.780 66.000 102.930 69.890 ;
        RECT 90.060 65.830 102.930 66.000 ;
        RECT 105.070 66.000 105.240 75.490 ;
        RECT 105.870 74.980 106.870 75.150 ;
        RECT 105.640 66.725 105.810 74.765 ;
        RECT 106.930 66.725 107.100 74.765 ;
        RECT 105.870 66.340 106.870 66.510 ;
        RECT 107.500 66.000 107.670 75.490 ;
        RECT 108.300 74.980 110.300 75.150 ;
        RECT 108.070 66.725 108.240 74.765 ;
        RECT 110.360 66.725 110.530 74.765 ;
        RECT 108.300 66.340 110.300 66.510 ;
        RECT 110.930 66.000 111.100 75.490 ;
        RECT 111.730 74.980 113.730 75.150 ;
        RECT 111.500 66.725 111.670 74.765 ;
        RECT 113.790 66.725 113.960 74.765 ;
        RECT 111.730 66.340 113.730 66.510 ;
        RECT 114.360 66.000 114.530 75.490 ;
        RECT 115.160 74.980 116.160 75.150 ;
        RECT 114.930 66.725 115.100 74.765 ;
        RECT 116.220 66.725 116.390 74.765 ;
        RECT 116.790 69.890 117.920 75.490 ;
        RECT 120.080 75.490 132.930 75.500 ;
        RECT 115.160 66.340 116.160 66.510 ;
        RECT 116.790 66.000 117.940 69.890 ;
        RECT 105.070 65.830 117.940 66.000 ;
        RECT 120.080 66.000 120.250 75.490 ;
        RECT 120.880 74.980 121.880 75.150 ;
        RECT 120.650 66.725 120.820 74.765 ;
        RECT 121.940 66.725 122.110 74.765 ;
        RECT 120.880 66.340 121.880 66.510 ;
        RECT 122.510 66.000 122.680 75.490 ;
        RECT 123.310 74.980 125.310 75.150 ;
        RECT 123.080 66.725 123.250 74.765 ;
        RECT 125.370 66.725 125.540 74.765 ;
        RECT 123.310 66.340 125.310 66.510 ;
        RECT 125.940 66.000 126.110 75.490 ;
        RECT 126.740 74.980 128.740 75.150 ;
        RECT 126.510 66.725 126.680 74.765 ;
        RECT 128.800 66.725 128.970 74.765 ;
        RECT 126.740 66.340 128.740 66.510 ;
        RECT 129.370 66.000 129.540 75.490 ;
        RECT 130.170 74.980 131.170 75.150 ;
        RECT 129.940 66.725 130.110 74.765 ;
        RECT 131.230 66.725 131.400 74.765 ;
        RECT 131.800 69.890 132.930 75.490 ;
        RECT 135.070 75.490 147.920 75.540 ;
        RECT 130.170 66.340 131.170 66.510 ;
        RECT 131.800 66.000 132.950 69.890 ;
        RECT 120.080 65.830 132.950 66.000 ;
        RECT 135.070 66.000 135.240 75.490 ;
        RECT 135.870 74.980 136.870 75.150 ;
        RECT 135.640 66.725 135.810 74.765 ;
        RECT 136.930 66.725 137.100 74.765 ;
        RECT 135.870 66.340 136.870 66.510 ;
        RECT 137.500 66.000 137.670 75.490 ;
        RECT 138.300 74.980 140.300 75.150 ;
        RECT 138.070 66.725 138.240 74.765 ;
        RECT 140.360 66.725 140.530 74.765 ;
        RECT 138.300 66.340 140.300 66.510 ;
        RECT 140.930 66.000 141.100 75.490 ;
        RECT 141.730 74.980 143.730 75.150 ;
        RECT 141.500 66.725 141.670 74.765 ;
        RECT 143.790 66.725 143.960 74.765 ;
        RECT 141.730 66.340 143.730 66.510 ;
        RECT 144.360 66.000 144.530 75.490 ;
        RECT 145.160 74.980 146.160 75.150 ;
        RECT 144.930 66.725 145.100 74.765 ;
        RECT 146.220 66.725 146.390 74.765 ;
        RECT 146.790 69.890 147.920 75.490 ;
        RECT 145.160 66.340 146.160 66.510 ;
        RECT 146.790 66.000 147.940 69.890 ;
        RECT 135.070 65.830 147.940 66.000 ;
        RECT 73.070 64.260 74.720 64.350 ;
        RECT 86.940 64.600 87.940 65.820 ;
        RECT 101.810 65.800 102.930 65.830 ;
        RECT 116.820 65.800 117.940 65.830 ;
        RECT 131.830 65.800 132.950 65.830 ;
        RECT 146.820 65.800 147.940 65.830 ;
        RECT 86.940 64.530 87.960 64.600 ;
        RECT 101.920 64.580 102.920 65.800 ;
        RECT 116.930 64.580 117.930 65.800 ;
        RECT 131.940 64.580 132.940 65.800 ;
        RECT 146.930 64.580 147.930 65.800 ;
        RECT 84.390 64.260 86.630 64.270 ;
        RECT 73.070 64.180 86.630 64.260 ;
        RECT 54.760 62.740 67.450 63.370 ;
        RECT 54.680 62.570 68.170 62.740 ;
        RECT 54.680 56.050 54.850 62.570 ;
        RECT 55.330 59.930 55.680 62.090 ;
        RECT 55.330 56.530 55.680 58.690 ;
        RECT 56.160 56.050 56.330 62.570 ;
        RECT 56.810 59.930 57.160 62.090 ;
        RECT 56.810 56.530 57.160 58.690 ;
        RECT 57.640 56.050 57.810 62.570 ;
        RECT 58.290 59.930 58.640 62.090 ;
        RECT 58.290 56.530 58.640 58.690 ;
        RECT 59.120 56.050 59.290 62.570 ;
        RECT 59.770 59.930 60.120 62.090 ;
        RECT 59.770 56.530 60.120 58.690 ;
        RECT 60.600 56.050 60.770 62.570 ;
        RECT 61.250 59.930 61.600 62.090 ;
        RECT 61.250 56.530 61.600 58.690 ;
        RECT 62.080 56.050 62.250 62.570 ;
        RECT 62.730 59.930 63.080 62.090 ;
        RECT 62.730 56.530 63.080 58.690 ;
        RECT 63.560 56.050 63.730 62.570 ;
        RECT 64.210 59.930 64.560 62.090 ;
        RECT 64.210 56.530 64.560 58.690 ;
        RECT 65.040 56.050 65.210 62.570 ;
        RECT 65.690 59.930 66.040 62.090 ;
        RECT 65.690 56.530 66.040 58.690 ;
        RECT 66.520 56.050 66.690 62.570 ;
        RECT 67.170 59.930 67.520 62.090 ;
        RECT 67.170 56.530 67.520 58.690 ;
        RECT 68.000 56.050 68.170 62.570 ;
        RECT 73.070 58.360 73.240 64.180 ;
        RECT 74.550 64.100 86.630 64.180 ;
        RECT 74.550 64.090 85.050 64.100 ;
        RECT 73.720 61.540 74.070 63.700 ;
        RECT 73.720 58.840 74.070 61.000 ;
        RECT 74.550 58.700 75.260 64.090 ;
        RECT 75.890 63.580 76.890 63.750 ;
        RECT 75.660 59.370 75.830 63.410 ;
        RECT 76.950 59.370 77.120 63.410 ;
        RECT 75.890 59.030 76.890 59.200 ;
        RECT 77.520 58.700 77.690 64.090 ;
        RECT 78.320 63.580 80.320 63.750 ;
        RECT 78.090 59.370 78.260 63.410 ;
        RECT 80.380 59.370 80.550 63.410 ;
        RECT 78.320 59.030 80.320 59.200 ;
        RECT 80.950 58.700 81.120 64.090 ;
        RECT 81.750 63.580 83.750 63.750 ;
        RECT 81.520 59.370 81.690 63.410 ;
        RECT 83.810 59.370 83.980 63.410 ;
        RECT 84.380 63.190 85.050 64.090 ;
        RECT 85.590 63.590 85.920 63.760 ;
        RECT 84.380 62.010 85.070 63.190 ;
        RECT 85.450 62.380 85.620 63.420 ;
        RECT 85.890 62.380 86.060 63.420 ;
        RECT 86.460 62.010 86.630 64.100 ;
        RECT 86.940 64.070 88.740 64.530 ;
        RECT 101.920 64.510 102.940 64.580 ;
        RECT 116.930 64.510 117.950 64.580 ;
        RECT 131.940 64.510 132.960 64.580 ;
        RECT 146.930 64.510 147.950 64.580 ;
        RECT 99.370 64.240 101.610 64.250 ;
        RECT 84.380 61.840 86.630 62.010 ;
        RECT 86.990 64.030 88.740 64.070 ;
        RECT 84.380 61.680 86.240 61.840 ;
        RECT 84.380 61.450 85.150 61.680 ;
        RECT 84.380 59.940 85.140 61.450 ;
        RECT 81.750 59.030 83.750 59.200 ;
        RECT 84.380 58.730 86.410 59.940 ;
        RECT 86.990 59.900 87.160 64.030 ;
        RECT 87.700 63.525 88.030 63.695 ;
        RECT 88.370 63.320 88.740 64.030 ;
        RECT 87.560 60.270 87.730 63.310 ;
        RECT 88.000 60.270 88.170 63.310 ;
        RECT 88.430 60.350 88.740 63.320 ;
        RECT 88.570 59.900 88.740 60.350 ;
        RECT 86.990 59.730 88.740 59.900 ;
        RECT 90.070 64.080 101.610 64.240 ;
        RECT 90.070 64.070 100.030 64.080 ;
        RECT 90.070 58.730 90.240 64.070 ;
        RECT 90.870 63.560 91.870 63.730 ;
        RECT 90.640 59.350 90.810 63.390 ;
        RECT 91.930 59.350 92.100 63.390 ;
        RECT 90.870 59.010 91.870 59.180 ;
        RECT 84.380 58.700 90.950 58.730 ;
        RECT 74.550 58.680 90.950 58.700 ;
        RECT 92.500 58.680 92.670 64.070 ;
        RECT 93.300 63.560 95.300 63.730 ;
        RECT 93.070 59.350 93.240 63.390 ;
        RECT 95.360 59.350 95.530 63.390 ;
        RECT 93.300 59.010 95.300 59.180 ;
        RECT 95.930 58.680 96.100 64.070 ;
        RECT 96.730 63.560 98.730 63.730 ;
        RECT 96.500 59.350 96.670 63.390 ;
        RECT 98.790 59.350 98.960 63.390 ;
        RECT 99.360 63.170 100.030 64.070 ;
        RECT 100.570 63.570 100.900 63.740 ;
        RECT 99.360 61.990 100.050 63.170 ;
        RECT 100.430 62.360 100.600 63.400 ;
        RECT 100.870 62.360 101.040 63.400 ;
        RECT 101.440 61.990 101.610 64.080 ;
        RECT 101.920 64.050 103.720 64.510 ;
        RECT 114.380 64.240 116.620 64.250 ;
        RECT 99.360 61.820 101.610 61.990 ;
        RECT 101.970 64.010 103.720 64.050 ;
        RECT 99.360 61.660 101.220 61.820 ;
        RECT 99.360 61.430 100.130 61.660 ;
        RECT 99.360 59.920 100.120 61.430 ;
        RECT 96.730 59.010 98.730 59.180 ;
        RECT 99.360 58.710 101.390 59.920 ;
        RECT 101.970 59.880 102.140 64.010 ;
        RECT 102.680 63.505 103.010 63.675 ;
        RECT 103.350 63.300 103.720 64.010 ;
        RECT 102.540 60.250 102.710 63.290 ;
        RECT 102.980 60.250 103.150 63.290 ;
        RECT 103.410 60.330 103.720 63.300 ;
        RECT 103.550 59.880 103.720 60.330 ;
        RECT 101.970 59.710 103.720 59.880 ;
        RECT 105.080 64.080 116.620 64.240 ;
        RECT 105.080 64.070 115.040 64.080 ;
        RECT 105.080 58.710 105.250 64.070 ;
        RECT 105.880 63.560 106.880 63.730 ;
        RECT 105.650 59.350 105.820 63.390 ;
        RECT 106.940 59.350 107.110 63.390 ;
        RECT 105.880 59.010 106.880 59.180 ;
        RECT 99.360 58.680 105.920 58.710 ;
        RECT 107.510 58.680 107.680 64.070 ;
        RECT 108.310 63.560 110.310 63.730 ;
        RECT 108.080 59.350 108.250 63.390 ;
        RECT 110.370 59.350 110.540 63.390 ;
        RECT 108.310 59.010 110.310 59.180 ;
        RECT 110.940 58.680 111.110 64.070 ;
        RECT 111.740 63.560 113.740 63.730 ;
        RECT 111.510 59.350 111.680 63.390 ;
        RECT 113.800 59.350 113.970 63.390 ;
        RECT 114.370 63.170 115.040 64.070 ;
        RECT 115.580 63.570 115.910 63.740 ;
        RECT 114.370 61.990 115.060 63.170 ;
        RECT 115.440 62.360 115.610 63.400 ;
        RECT 115.880 62.360 116.050 63.400 ;
        RECT 116.450 61.990 116.620 64.080 ;
        RECT 116.930 64.050 118.730 64.510 ;
        RECT 129.390 64.240 131.630 64.250 ;
        RECT 114.370 61.820 116.620 61.990 ;
        RECT 116.980 64.010 118.730 64.050 ;
        RECT 114.370 61.660 116.230 61.820 ;
        RECT 114.370 61.430 115.140 61.660 ;
        RECT 114.370 59.920 115.130 61.430 ;
        RECT 111.740 59.010 113.740 59.180 ;
        RECT 114.370 58.680 116.400 59.920 ;
        RECT 116.980 59.880 117.150 64.010 ;
        RECT 117.690 63.505 118.020 63.675 ;
        RECT 118.360 63.300 118.730 64.010 ;
        RECT 117.550 60.250 117.720 63.290 ;
        RECT 117.990 60.250 118.160 63.290 ;
        RECT 118.420 60.330 118.730 63.300 ;
        RECT 118.560 59.880 118.730 60.330 ;
        RECT 116.980 59.710 118.730 59.880 ;
        RECT 120.090 64.080 131.630 64.240 ;
        RECT 120.090 64.070 130.050 64.080 ;
        RECT 120.090 58.680 120.260 64.070 ;
        RECT 120.890 63.560 121.890 63.730 ;
        RECT 120.660 59.350 120.830 63.390 ;
        RECT 121.950 59.350 122.120 63.390 ;
        RECT 120.890 59.010 121.890 59.180 ;
        RECT 122.520 58.680 122.690 64.070 ;
        RECT 123.320 63.560 125.320 63.730 ;
        RECT 123.090 59.350 123.260 63.390 ;
        RECT 125.380 59.350 125.550 63.390 ;
        RECT 123.320 59.010 125.320 59.180 ;
        RECT 125.950 58.680 126.120 64.070 ;
        RECT 126.750 63.560 128.750 63.730 ;
        RECT 126.520 59.350 126.690 63.390 ;
        RECT 128.810 59.350 128.980 63.390 ;
        RECT 129.380 63.170 130.050 64.070 ;
        RECT 130.590 63.570 130.920 63.740 ;
        RECT 129.380 61.990 130.070 63.170 ;
        RECT 130.450 62.360 130.620 63.400 ;
        RECT 130.890 62.360 131.060 63.400 ;
        RECT 131.460 61.990 131.630 64.080 ;
        RECT 131.940 64.050 133.740 64.510 ;
        RECT 144.380 64.240 146.620 64.250 ;
        RECT 129.380 61.820 131.630 61.990 ;
        RECT 131.990 64.010 133.740 64.050 ;
        RECT 129.380 61.660 131.240 61.820 ;
        RECT 129.380 61.430 130.150 61.660 ;
        RECT 129.380 59.920 130.140 61.430 ;
        RECT 126.750 59.010 128.750 59.180 ;
        RECT 129.380 58.720 131.410 59.920 ;
        RECT 131.990 59.880 132.160 64.010 ;
        RECT 132.700 63.505 133.030 63.675 ;
        RECT 133.370 63.300 133.740 64.010 ;
        RECT 132.560 60.250 132.730 63.290 ;
        RECT 133.000 60.250 133.170 63.290 ;
        RECT 133.430 60.330 133.740 63.300 ;
        RECT 133.570 59.880 133.740 60.330 ;
        RECT 131.990 59.710 133.740 59.880 ;
        RECT 135.080 64.080 146.620 64.240 ;
        RECT 135.080 64.070 145.040 64.080 ;
        RECT 135.080 58.720 135.250 64.070 ;
        RECT 135.880 63.560 136.880 63.730 ;
        RECT 135.650 59.350 135.820 63.390 ;
        RECT 136.940 59.350 137.110 63.390 ;
        RECT 135.880 59.010 136.880 59.180 ;
        RECT 129.380 58.680 135.620 58.720 ;
        RECT 137.510 58.680 137.680 64.070 ;
        RECT 138.310 63.560 140.310 63.730 ;
        RECT 138.080 59.350 138.250 63.390 ;
        RECT 140.370 59.350 140.540 63.390 ;
        RECT 138.310 59.010 140.310 59.180 ;
        RECT 140.940 58.680 141.110 64.070 ;
        RECT 141.740 63.560 143.740 63.730 ;
        RECT 141.510 59.350 141.680 63.390 ;
        RECT 143.800 59.350 143.970 63.390 ;
        RECT 144.370 63.170 145.040 64.070 ;
        RECT 145.580 63.570 145.910 63.740 ;
        RECT 144.370 61.990 145.060 63.170 ;
        RECT 145.440 62.360 145.610 63.400 ;
        RECT 145.880 62.360 146.050 63.400 ;
        RECT 146.450 61.990 146.620 64.080 ;
        RECT 146.930 64.050 148.730 64.510 ;
        RECT 144.370 61.820 146.620 61.990 ;
        RECT 146.980 64.010 148.730 64.050 ;
        RECT 144.370 61.660 146.230 61.820 ;
        RECT 144.370 61.430 145.140 61.660 ;
        RECT 144.370 59.920 145.130 61.430 ;
        RECT 141.740 59.010 143.740 59.180 ;
        RECT 144.370 58.680 146.400 59.920 ;
        RECT 146.980 59.880 147.150 64.010 ;
        RECT 147.690 63.505 148.020 63.675 ;
        RECT 148.360 63.300 148.730 64.010 ;
        RECT 147.550 60.250 147.720 63.290 ;
        RECT 147.990 60.250 148.160 63.290 ;
        RECT 148.420 60.330 148.730 63.300 ;
        RECT 148.560 59.880 148.730 60.330 ;
        RECT 146.980 59.710 148.730 59.880 ;
        RECT 74.550 58.360 146.400 58.680 ;
        RECT 54.680 55.880 68.170 56.050 ;
        RECT 71.590 58.190 146.400 58.360 ;
        RECT 54.680 50.060 54.850 55.880 ;
        RECT 55.330 53.240 55.680 55.400 ;
        RECT 55.330 50.540 55.680 52.700 ;
        RECT 56.160 50.060 56.330 55.880 ;
        RECT 56.810 53.240 57.160 55.400 ;
        RECT 56.810 50.540 57.160 52.700 ;
        RECT 57.640 50.060 57.810 55.880 ;
        RECT 58.290 53.240 58.640 55.400 ;
        RECT 58.290 50.540 58.640 52.700 ;
        RECT 59.120 50.060 59.290 55.880 ;
        RECT 59.770 53.240 60.120 55.400 ;
        RECT 59.770 50.540 60.120 52.700 ;
        RECT 60.600 50.060 60.770 55.880 ;
        RECT 61.250 53.240 61.600 55.400 ;
        RECT 61.250 50.540 61.600 52.700 ;
        RECT 62.080 50.060 62.250 55.880 ;
        RECT 62.730 53.240 63.080 55.400 ;
        RECT 62.730 50.540 63.080 52.700 ;
        RECT 63.560 50.060 63.730 55.880 ;
        RECT 64.210 53.240 64.560 55.400 ;
        RECT 64.210 50.540 64.560 52.700 ;
        RECT 65.040 50.060 65.210 55.880 ;
        RECT 54.680 49.890 65.210 50.060 ;
        RECT 71.590 52.370 71.760 58.190 ;
        RECT 72.240 55.550 72.590 57.710 ;
        RECT 72.240 52.850 72.590 55.010 ;
        RECT 73.070 52.370 73.240 58.190 ;
        RECT 74.550 58.030 146.400 58.190 ;
        RECT 73.720 55.550 74.070 57.710 ;
        RECT 73.720 52.850 74.070 55.010 ;
        RECT 74.550 52.370 74.720 58.030 ;
        RECT 84.490 58.020 146.400 58.030 ;
        RECT 86.120 58.010 146.400 58.020 ;
        RECT 86.120 58.000 90.950 58.010 ;
        RECT 99.470 58.000 105.920 58.010 ;
        RECT 114.480 58.000 120.280 58.010 ;
        RECT 129.490 58.000 135.620 58.010 ;
        RECT 144.480 58.000 146.400 58.010 ;
        RECT 101.090 57.980 105.920 58.000 ;
        RECT 115.450 57.950 120.280 58.000 ;
        RECT 130.790 57.990 135.620 58.000 ;
        RECT 132.390 57.490 135.520 57.510 ;
        RECT 75.120 57.430 87.920 57.470 ;
        RECT 102.260 57.460 105.390 57.470 ;
        RECT 117.240 57.460 120.370 57.490 ;
        RECT 132.390 57.460 147.930 57.490 ;
        RECT 90.100 57.430 147.930 57.460 ;
        RECT 75.120 57.380 147.930 57.430 ;
        RECT 75.120 56.670 147.940 57.380 ;
        RECT 71.590 52.200 74.720 52.370 ;
        RECT 54.760 48.350 67.560 48.460 ;
        RECT 54.760 47.660 67.570 48.350 ;
        RECT 54.720 47.490 67.570 47.660 ;
        RECT 54.720 38.000 54.890 47.490 ;
        RECT 55.520 46.980 56.520 47.150 ;
        RECT 55.290 38.725 55.460 46.765 ;
        RECT 56.580 38.725 56.750 46.765 ;
        RECT 55.520 38.340 56.520 38.510 ;
        RECT 57.150 38.000 57.320 47.490 ;
        RECT 57.950 46.980 59.950 47.150 ;
        RECT 57.720 38.725 57.890 46.765 ;
        RECT 60.010 38.725 60.180 46.765 ;
        RECT 57.950 38.340 59.950 38.510 ;
        RECT 60.580 38.000 60.750 47.490 ;
        RECT 61.380 46.980 63.380 47.150 ;
        RECT 61.150 38.725 61.320 46.765 ;
        RECT 63.440 38.725 63.610 46.765 ;
        RECT 61.380 38.340 63.380 38.510 ;
        RECT 64.010 38.000 64.180 47.490 ;
        RECT 64.810 46.980 65.810 47.150 ;
        RECT 64.580 38.725 64.750 46.765 ;
        RECT 65.870 38.725 66.040 46.765 ;
        RECT 66.440 41.890 67.570 47.490 ;
        RECT 71.590 46.380 71.760 52.200 ;
        RECT 72.240 49.560 72.590 51.720 ;
        RECT 72.240 46.860 72.590 49.020 ;
        RECT 73.070 46.380 73.240 52.200 ;
        RECT 73.720 49.560 74.070 51.720 ;
        RECT 73.720 46.860 74.070 49.020 ;
        RECT 74.550 46.380 74.720 52.200 ;
        RECT 75.080 56.560 147.940 56.670 ;
        RECT 75.080 56.540 132.930 56.560 ;
        RECT 75.080 56.520 117.950 56.540 ;
        RECT 75.080 56.500 102.910 56.520 ;
        RECT 75.080 47.010 75.250 56.500 ;
        RECT 75.880 55.990 76.880 56.160 ;
        RECT 75.650 47.735 75.820 55.775 ;
        RECT 76.940 47.735 77.110 55.775 ;
        RECT 75.880 47.350 76.880 47.520 ;
        RECT 77.510 47.010 77.680 56.500 ;
        RECT 78.310 55.990 80.310 56.160 ;
        RECT 78.080 47.735 78.250 55.775 ;
        RECT 80.370 47.735 80.540 55.775 ;
        RECT 78.310 47.350 80.310 47.520 ;
        RECT 80.940 47.010 81.110 56.500 ;
        RECT 81.740 55.990 83.740 56.160 ;
        RECT 81.510 47.735 81.680 55.775 ;
        RECT 83.800 47.735 83.970 55.775 ;
        RECT 81.740 47.350 83.740 47.520 ;
        RECT 84.370 47.010 84.540 56.500 ;
        RECT 86.800 56.490 102.910 56.500 ;
        RECT 86.800 56.480 90.490 56.490 ;
        RECT 85.170 55.990 86.170 56.160 ;
        RECT 84.940 47.735 85.110 55.775 ;
        RECT 86.230 47.735 86.400 55.775 ;
        RECT 86.800 50.900 87.930 56.480 ;
        RECT 85.170 47.350 86.170 47.520 ;
        RECT 86.800 47.010 87.950 50.900 ;
        RECT 75.080 46.840 87.950 47.010 ;
        RECT 86.830 46.810 87.950 46.840 ;
        RECT 90.060 47.000 90.230 56.480 ;
        RECT 90.860 55.980 91.860 56.150 ;
        RECT 90.630 47.725 90.800 55.765 ;
        RECT 91.920 47.725 92.090 55.765 ;
        RECT 90.860 47.340 91.860 47.510 ;
        RECT 92.490 47.000 92.660 56.490 ;
        RECT 93.290 55.980 95.290 56.150 ;
        RECT 93.060 47.725 93.230 55.765 ;
        RECT 95.350 47.725 95.520 55.765 ;
        RECT 93.290 47.340 95.290 47.510 ;
        RECT 95.920 47.000 96.090 56.490 ;
        RECT 96.720 55.980 98.720 56.150 ;
        RECT 96.490 47.725 96.660 55.765 ;
        RECT 98.780 47.725 98.950 55.765 ;
        RECT 96.720 47.340 98.720 47.510 ;
        RECT 99.350 47.000 99.520 56.490 ;
        RECT 100.150 55.980 101.150 56.150 ;
        RECT 99.920 47.725 100.090 55.765 ;
        RECT 101.210 47.725 101.380 55.765 ;
        RECT 101.780 50.890 102.910 56.490 ;
        RECT 105.100 56.490 117.950 56.520 ;
        RECT 100.150 47.340 101.150 47.510 ;
        RECT 101.780 47.000 102.930 50.890 ;
        RECT 90.060 46.830 102.930 47.000 ;
        RECT 105.100 47.000 105.270 56.490 ;
        RECT 105.900 55.980 106.900 56.150 ;
        RECT 105.670 47.725 105.840 55.765 ;
        RECT 106.960 47.725 107.130 55.765 ;
        RECT 105.900 47.340 106.900 47.510 ;
        RECT 107.530 47.000 107.700 56.490 ;
        RECT 108.330 55.980 110.330 56.150 ;
        RECT 108.100 47.725 108.270 55.765 ;
        RECT 110.390 47.725 110.560 55.765 ;
        RECT 108.330 47.340 110.330 47.510 ;
        RECT 110.960 47.000 111.130 56.490 ;
        RECT 111.760 55.980 113.760 56.150 ;
        RECT 111.530 47.725 111.700 55.765 ;
        RECT 113.820 47.725 113.990 55.765 ;
        RECT 111.760 47.340 113.760 47.510 ;
        RECT 114.390 47.000 114.560 56.490 ;
        RECT 115.190 55.980 116.190 56.150 ;
        RECT 114.960 47.725 115.130 55.765 ;
        RECT 116.250 47.725 116.420 55.765 ;
        RECT 116.820 50.890 117.950 56.490 ;
        RECT 120.080 56.490 132.930 56.540 ;
        RECT 115.190 47.340 116.190 47.510 ;
        RECT 116.820 47.000 117.970 50.890 ;
        RECT 105.100 46.830 117.970 47.000 ;
        RECT 120.080 47.000 120.250 56.490 ;
        RECT 120.880 55.980 121.880 56.150 ;
        RECT 120.650 47.725 120.820 55.765 ;
        RECT 121.940 47.725 122.110 55.765 ;
        RECT 120.880 47.340 121.880 47.510 ;
        RECT 122.510 47.000 122.680 56.490 ;
        RECT 123.310 55.980 125.310 56.150 ;
        RECT 123.080 47.725 123.250 55.765 ;
        RECT 125.370 47.725 125.540 55.765 ;
        RECT 123.310 47.340 125.310 47.510 ;
        RECT 125.940 47.000 126.110 56.490 ;
        RECT 126.740 55.980 128.740 56.150 ;
        RECT 126.510 47.725 126.680 55.765 ;
        RECT 128.800 47.725 128.970 55.765 ;
        RECT 126.740 47.340 128.740 47.510 ;
        RECT 129.370 47.000 129.540 56.490 ;
        RECT 130.170 55.980 131.170 56.150 ;
        RECT 129.940 47.725 130.110 55.765 ;
        RECT 131.230 47.725 131.400 55.765 ;
        RECT 131.800 50.890 132.930 56.490 ;
        RECT 135.090 56.520 147.940 56.560 ;
        RECT 130.170 47.340 131.170 47.510 ;
        RECT 131.800 47.000 132.950 50.890 ;
        RECT 120.080 46.830 132.950 47.000 ;
        RECT 135.090 47.030 135.260 56.520 ;
        RECT 135.890 56.010 136.890 56.180 ;
        RECT 135.660 47.755 135.830 55.795 ;
        RECT 136.950 47.755 137.120 55.795 ;
        RECT 135.890 47.370 136.890 47.540 ;
        RECT 137.520 47.030 137.690 56.520 ;
        RECT 138.320 56.010 140.320 56.180 ;
        RECT 138.090 47.755 138.260 55.795 ;
        RECT 140.380 47.755 140.550 55.795 ;
        RECT 138.320 47.370 140.320 47.540 ;
        RECT 140.950 47.030 141.120 56.520 ;
        RECT 141.750 56.010 143.750 56.180 ;
        RECT 141.520 47.755 141.690 55.795 ;
        RECT 143.810 47.755 143.980 55.795 ;
        RECT 141.750 47.370 143.750 47.540 ;
        RECT 144.380 47.030 144.550 56.520 ;
        RECT 145.180 56.010 146.180 56.180 ;
        RECT 144.950 47.755 145.120 55.795 ;
        RECT 146.240 47.755 146.410 55.795 ;
        RECT 146.810 50.920 147.940 56.520 ;
        RECT 145.180 47.370 146.180 47.540 ;
        RECT 146.810 47.030 147.960 50.920 ;
        RECT 135.090 46.860 147.960 47.030 ;
        RECT 146.840 46.830 147.960 46.860 ;
        RECT 71.590 46.210 74.720 46.380 ;
        RECT 64.810 38.340 65.810 38.510 ;
        RECT 66.440 38.000 67.590 41.890 ;
        RECT 54.720 37.830 67.590 38.000 ;
        RECT 66.470 37.800 67.590 37.830 ;
        RECT 71.590 40.390 71.760 46.210 ;
        RECT 72.240 43.570 72.590 45.730 ;
        RECT 72.240 40.870 72.590 43.030 ;
        RECT 73.070 40.390 73.240 46.210 ;
        RECT 73.720 43.570 74.070 45.730 ;
        RECT 73.720 40.870 74.070 43.030 ;
        RECT 74.550 40.390 74.720 46.210 ;
        RECT 86.940 45.590 87.940 46.810 ;
        RECT 101.810 46.800 102.930 46.830 ;
        RECT 116.850 46.800 117.970 46.830 ;
        RECT 131.830 46.800 132.950 46.830 ;
        RECT 86.940 45.520 87.960 45.590 ;
        RECT 101.920 45.580 102.920 46.800 ;
        RECT 116.960 45.580 117.960 46.800 ;
        RECT 131.940 45.580 132.940 46.800 ;
        RECT 146.950 45.610 147.950 46.830 ;
        RECT 84.390 45.250 86.630 45.260 ;
        RECT 71.590 40.220 74.720 40.390 ;
        RECT 66.580 36.580 67.580 37.800 ;
        RECT 64.030 36.240 66.270 36.250 ;
        RECT 54.730 36.080 66.270 36.240 ;
        RECT 54.730 36.070 64.690 36.080 ;
        RECT 54.730 30.680 54.900 36.070 ;
        RECT 55.530 35.560 56.530 35.730 ;
        RECT 55.300 31.350 55.470 35.390 ;
        RECT 56.590 31.350 56.760 35.390 ;
        RECT 55.530 31.010 56.530 31.180 ;
        RECT 57.160 30.680 57.330 36.070 ;
        RECT 57.960 35.560 59.960 35.730 ;
        RECT 57.730 31.350 57.900 35.390 ;
        RECT 60.020 31.350 60.190 35.390 ;
        RECT 57.960 31.010 59.960 31.180 ;
        RECT 60.590 30.680 60.760 36.070 ;
        RECT 61.390 35.560 63.390 35.730 ;
        RECT 61.160 31.350 61.330 35.390 ;
        RECT 63.450 31.350 63.620 35.390 ;
        RECT 64.020 35.170 64.690 36.070 ;
        RECT 65.230 35.570 65.560 35.740 ;
        RECT 64.020 33.990 64.710 35.170 ;
        RECT 65.090 34.360 65.260 35.400 ;
        RECT 65.530 34.360 65.700 35.400 ;
        RECT 66.100 33.990 66.270 36.080 ;
        RECT 66.580 36.190 67.600 36.580 ;
        RECT 66.580 36.050 68.380 36.190 ;
        RECT 64.020 33.820 66.270 33.990 ;
        RECT 66.630 36.020 68.380 36.050 ;
        RECT 66.630 36.010 67.600 36.020 ;
        RECT 64.020 33.660 65.880 33.820 ;
        RECT 64.020 33.430 64.790 33.660 ;
        RECT 64.020 31.920 64.780 33.430 ;
        RECT 61.390 31.010 63.390 31.180 ;
        RECT 64.020 30.680 66.050 31.920 ;
        RECT 66.630 31.880 66.800 36.010 ;
        RECT 67.340 35.505 67.670 35.675 ;
        RECT 67.200 32.250 67.370 35.290 ;
        RECT 67.640 32.250 67.810 35.290 ;
        RECT 68.210 31.880 68.380 36.020 ;
        RECT 66.630 31.710 68.380 31.880 ;
        RECT 71.590 34.400 71.760 40.220 ;
        RECT 72.240 37.580 72.590 39.740 ;
        RECT 72.240 34.880 72.590 37.040 ;
        RECT 73.070 34.400 73.240 40.220 ;
        RECT 73.720 37.580 74.070 39.740 ;
        RECT 73.720 34.880 74.070 37.040 ;
        RECT 74.550 34.400 74.720 40.220 ;
        RECT 75.090 45.090 86.630 45.250 ;
        RECT 75.090 45.080 85.050 45.090 ;
        RECT 75.090 39.690 75.260 45.080 ;
        RECT 75.890 44.570 76.890 44.740 ;
        RECT 75.660 40.360 75.830 44.400 ;
        RECT 76.950 40.360 77.120 44.400 ;
        RECT 75.890 40.020 76.890 40.190 ;
        RECT 77.520 39.690 77.690 45.080 ;
        RECT 78.320 44.570 80.320 44.740 ;
        RECT 78.090 40.360 78.260 44.400 ;
        RECT 80.380 40.360 80.550 44.400 ;
        RECT 78.320 40.020 80.320 40.190 ;
        RECT 80.950 39.690 81.120 45.080 ;
        RECT 81.750 44.570 83.750 44.740 ;
        RECT 81.520 40.360 81.690 44.400 ;
        RECT 83.810 40.360 83.980 44.400 ;
        RECT 84.380 44.180 85.050 45.080 ;
        RECT 85.590 44.580 85.920 44.750 ;
        RECT 84.380 43.000 85.070 44.180 ;
        RECT 85.450 43.370 85.620 44.410 ;
        RECT 85.890 43.370 86.060 44.410 ;
        RECT 86.460 43.000 86.630 45.090 ;
        RECT 86.940 45.060 88.740 45.520 ;
        RECT 101.920 45.510 102.940 45.580 ;
        RECT 116.960 45.510 117.980 45.580 ;
        RECT 131.940 45.510 132.960 45.580 ;
        RECT 146.950 45.540 147.970 45.610 ;
        RECT 99.370 45.240 101.610 45.250 ;
        RECT 84.380 42.830 86.630 43.000 ;
        RECT 86.990 45.020 88.740 45.060 ;
        RECT 84.380 42.670 86.240 42.830 ;
        RECT 84.380 42.440 85.150 42.670 ;
        RECT 84.380 40.930 85.140 42.440 ;
        RECT 81.750 40.020 83.750 40.190 ;
        RECT 84.380 39.710 86.410 40.930 ;
        RECT 86.990 40.890 87.160 45.020 ;
        RECT 87.700 44.515 88.030 44.685 ;
        RECT 88.370 44.310 88.740 45.020 ;
        RECT 87.560 41.260 87.730 44.300 ;
        RECT 88.000 41.260 88.170 44.300 ;
        RECT 88.430 41.340 88.740 44.310 ;
        RECT 88.570 40.890 88.740 41.340 ;
        RECT 86.990 40.720 88.740 40.890 ;
        RECT 90.070 45.080 101.610 45.240 ;
        RECT 90.070 45.070 100.030 45.080 ;
        RECT 90.070 39.710 90.240 45.070 ;
        RECT 90.870 44.560 91.870 44.730 ;
        RECT 90.640 40.350 90.810 44.390 ;
        RECT 91.930 40.350 92.100 44.390 ;
        RECT 90.870 40.010 91.870 40.180 ;
        RECT 84.380 39.690 90.750 39.710 ;
        RECT 75.090 39.680 90.750 39.690 ;
        RECT 92.500 39.680 92.670 45.070 ;
        RECT 93.300 44.560 95.300 44.730 ;
        RECT 93.070 40.350 93.240 44.390 ;
        RECT 95.360 40.350 95.530 44.390 ;
        RECT 93.300 40.010 95.300 40.180 ;
        RECT 95.930 39.680 96.100 45.070 ;
        RECT 96.730 44.560 98.730 44.730 ;
        RECT 96.500 40.350 96.670 44.390 ;
        RECT 98.790 40.350 98.960 44.390 ;
        RECT 99.360 44.170 100.030 45.070 ;
        RECT 100.570 44.570 100.900 44.740 ;
        RECT 99.360 42.990 100.050 44.170 ;
        RECT 100.430 43.360 100.600 44.400 ;
        RECT 100.870 43.360 101.040 44.400 ;
        RECT 101.440 42.990 101.610 45.080 ;
        RECT 101.920 45.050 103.720 45.510 ;
        RECT 114.410 45.240 116.650 45.250 ;
        RECT 99.360 42.820 101.610 42.990 ;
        RECT 101.970 45.010 103.720 45.050 ;
        RECT 99.360 42.660 101.220 42.820 ;
        RECT 99.360 42.430 100.130 42.660 ;
        RECT 99.360 40.920 100.120 42.430 ;
        RECT 96.730 40.010 98.730 40.180 ;
        RECT 99.360 39.730 101.390 40.920 ;
        RECT 101.970 40.880 102.140 45.010 ;
        RECT 102.680 44.505 103.010 44.675 ;
        RECT 103.350 44.300 103.720 45.010 ;
        RECT 102.540 41.250 102.710 44.290 ;
        RECT 102.980 41.250 103.150 44.290 ;
        RECT 103.410 41.330 103.720 44.300 ;
        RECT 103.550 40.880 103.720 41.330 ;
        RECT 101.970 40.710 103.720 40.880 ;
        RECT 105.110 45.080 116.650 45.240 ;
        RECT 105.110 45.070 115.070 45.080 ;
        RECT 105.110 39.730 105.280 45.070 ;
        RECT 105.910 44.560 106.910 44.730 ;
        RECT 105.680 40.350 105.850 44.390 ;
        RECT 106.970 40.350 107.140 44.390 ;
        RECT 105.910 40.010 106.910 40.180 ;
        RECT 99.360 39.680 105.750 39.730 ;
        RECT 107.540 39.680 107.710 45.070 ;
        RECT 108.340 44.560 110.340 44.730 ;
        RECT 108.110 40.350 108.280 44.390 ;
        RECT 110.400 40.350 110.570 44.390 ;
        RECT 108.340 40.010 110.340 40.180 ;
        RECT 110.970 39.680 111.140 45.070 ;
        RECT 111.770 44.560 113.770 44.730 ;
        RECT 111.540 40.350 111.710 44.390 ;
        RECT 113.830 40.350 114.000 44.390 ;
        RECT 114.400 44.170 115.070 45.070 ;
        RECT 115.610 44.570 115.940 44.740 ;
        RECT 114.400 42.990 115.090 44.170 ;
        RECT 115.470 43.360 115.640 44.400 ;
        RECT 115.910 43.360 116.080 44.400 ;
        RECT 116.480 42.990 116.650 45.080 ;
        RECT 116.960 45.050 118.760 45.510 ;
        RECT 129.390 45.240 131.630 45.250 ;
        RECT 114.400 42.820 116.650 42.990 ;
        RECT 117.010 45.010 118.760 45.050 ;
        RECT 114.400 42.660 116.260 42.820 ;
        RECT 114.400 42.430 115.170 42.660 ;
        RECT 114.400 40.920 115.160 42.430 ;
        RECT 111.770 40.010 113.770 40.180 ;
        RECT 114.400 39.690 116.430 40.920 ;
        RECT 117.010 40.880 117.180 45.010 ;
        RECT 117.720 44.505 118.050 44.675 ;
        RECT 118.390 44.300 118.760 45.010 ;
        RECT 117.580 41.250 117.750 44.290 ;
        RECT 118.020 41.250 118.190 44.290 ;
        RECT 118.450 41.330 118.760 44.300 ;
        RECT 118.590 40.880 118.760 41.330 ;
        RECT 117.010 40.710 118.760 40.880 ;
        RECT 120.090 45.080 131.630 45.240 ;
        RECT 120.090 45.070 130.050 45.080 ;
        RECT 120.090 39.690 120.260 45.070 ;
        RECT 120.890 44.560 121.890 44.730 ;
        RECT 120.660 40.350 120.830 44.390 ;
        RECT 121.950 40.350 122.120 44.390 ;
        RECT 120.890 40.010 121.890 40.180 ;
        RECT 114.400 39.680 121.040 39.690 ;
        RECT 122.520 39.680 122.690 45.070 ;
        RECT 123.320 44.560 125.320 44.730 ;
        RECT 123.090 40.350 123.260 44.390 ;
        RECT 125.380 40.350 125.550 44.390 ;
        RECT 123.320 40.010 125.320 40.180 ;
        RECT 125.950 39.680 126.120 45.070 ;
        RECT 126.750 44.560 128.750 44.730 ;
        RECT 126.520 40.350 126.690 44.390 ;
        RECT 128.810 40.350 128.980 44.390 ;
        RECT 129.380 44.170 130.050 45.070 ;
        RECT 130.590 44.570 130.920 44.740 ;
        RECT 129.380 42.990 130.070 44.170 ;
        RECT 130.450 43.360 130.620 44.400 ;
        RECT 130.890 43.360 131.060 44.400 ;
        RECT 131.460 42.990 131.630 45.080 ;
        RECT 131.940 45.050 133.740 45.510 ;
        RECT 144.400 45.270 146.640 45.280 ;
        RECT 129.380 42.820 131.630 42.990 ;
        RECT 131.990 45.010 133.740 45.050 ;
        RECT 129.380 42.660 131.240 42.820 ;
        RECT 129.380 42.430 130.150 42.660 ;
        RECT 129.380 40.920 130.140 42.430 ;
        RECT 126.750 40.010 128.750 40.180 ;
        RECT 129.380 39.680 131.410 40.920 ;
        RECT 131.990 40.880 132.160 45.010 ;
        RECT 132.700 44.505 133.030 44.675 ;
        RECT 133.370 44.300 133.740 45.010 ;
        RECT 132.560 41.250 132.730 44.290 ;
        RECT 133.000 41.250 133.170 44.290 ;
        RECT 133.430 41.330 133.740 44.300 ;
        RECT 133.570 40.880 133.740 41.330 ;
        RECT 131.990 40.710 133.740 40.880 ;
        RECT 135.100 45.110 146.640 45.270 ;
        RECT 135.100 45.100 145.060 45.110 ;
        RECT 135.100 39.710 135.270 45.100 ;
        RECT 135.900 44.590 136.900 44.760 ;
        RECT 135.670 40.380 135.840 44.420 ;
        RECT 136.960 40.380 137.130 44.420 ;
        RECT 135.900 40.040 136.900 40.210 ;
        RECT 137.530 39.710 137.700 45.100 ;
        RECT 138.330 44.590 140.330 44.760 ;
        RECT 138.100 40.380 138.270 44.420 ;
        RECT 140.390 40.380 140.560 44.420 ;
        RECT 138.330 40.040 140.330 40.210 ;
        RECT 140.960 39.710 141.130 45.100 ;
        RECT 141.760 44.590 143.760 44.760 ;
        RECT 141.530 40.380 141.700 44.420 ;
        RECT 143.820 40.380 143.990 44.420 ;
        RECT 144.390 44.200 145.060 45.100 ;
        RECT 145.600 44.600 145.930 44.770 ;
        RECT 144.390 43.020 145.080 44.200 ;
        RECT 145.460 43.390 145.630 44.430 ;
        RECT 145.900 43.390 146.070 44.430 ;
        RECT 146.470 43.020 146.640 45.110 ;
        RECT 146.950 45.080 148.750 45.540 ;
        RECT 144.390 42.850 146.640 43.020 ;
        RECT 147.000 45.040 148.750 45.080 ;
        RECT 144.390 42.690 146.250 42.850 ;
        RECT 144.390 42.460 145.160 42.690 ;
        RECT 144.390 40.950 145.150 42.460 ;
        RECT 141.760 40.040 143.760 40.210 ;
        RECT 144.390 39.710 146.420 40.950 ;
        RECT 147.000 40.910 147.170 45.040 ;
        RECT 147.710 44.535 148.040 44.705 ;
        RECT 148.380 44.330 148.750 45.040 ;
        RECT 147.570 41.280 147.740 44.320 ;
        RECT 148.010 41.280 148.180 44.320 ;
        RECT 148.440 41.360 148.750 44.330 ;
        RECT 148.580 40.910 148.750 41.360 ;
        RECT 147.000 40.740 148.750 40.910 ;
        RECT 135.100 39.680 146.420 39.710 ;
        RECT 75.090 39.510 146.420 39.680 ;
        RECT 75.100 39.040 146.420 39.510 ;
        RECT 75.100 39.020 136.020 39.040 ;
        RECT 144.500 39.030 146.420 39.040 ;
        RECT 84.490 39.010 136.020 39.020 ;
        RECT 85.920 38.980 90.750 39.010 ;
        RECT 99.470 39.000 105.750 39.010 ;
        RECT 114.510 39.000 121.040 39.010 ;
        RECT 129.490 39.000 136.020 39.010 ;
        RECT 116.210 38.960 121.040 39.000 ;
        RECT 131.190 38.950 136.020 39.000 ;
        RECT 117.460 38.460 120.590 38.490 ;
        RECT 75.160 38.440 87.960 38.460 ;
        RECT 90.100 38.440 102.900 38.460 ;
        RECT 75.160 38.430 102.900 38.440 ;
        RECT 105.110 38.430 132.950 38.460 ;
        RECT 135.110 38.430 147.910 38.460 ;
        RECT 75.160 38.350 147.910 38.430 ;
        RECT 75.160 37.660 147.920 38.350 ;
        RECT 71.590 34.230 74.720 34.400 ;
        RECT 54.730 30.500 66.050 30.680 ;
        RECT 54.740 30.010 66.050 30.500 ;
        RECT 64.130 30.000 66.050 30.010 ;
        RECT 61.490 28.260 66.810 29.180 ;
        RECT 71.590 28.410 71.760 34.230 ;
        RECT 72.240 31.590 72.590 33.750 ;
        RECT 72.240 28.890 72.590 31.050 ;
        RECT 73.070 28.410 73.240 34.230 ;
        RECT 73.720 31.590 74.070 33.750 ;
        RECT 73.720 28.890 74.070 31.050 ;
        RECT 74.550 28.410 74.720 34.230 ;
        RECT 61.490 28.160 63.250 28.260 ;
        RECT 61.500 22.770 61.670 28.160 ;
        RECT 62.210 27.750 62.540 27.920 ;
        RECT 62.070 23.495 62.240 27.535 ;
        RECT 62.510 23.495 62.680 27.535 ;
        RECT 62.210 23.110 62.540 23.280 ;
        RECT 63.080 22.770 63.250 28.160 ;
        RECT 66.620 28.160 66.810 28.260 ;
        RECT 70.110 28.240 74.720 28.410 ;
        RECT 64.290 27.750 64.620 27.920 ;
        RECT 65.250 27.750 65.580 27.920 ;
        RECT 63.650 23.495 63.820 27.535 ;
        RECT 64.130 23.495 64.300 27.535 ;
        RECT 64.610 23.495 64.780 27.535 ;
        RECT 65.090 23.495 65.260 27.535 ;
        RECT 65.570 23.495 65.740 27.535 ;
        RECT 66.050 23.495 66.220 27.535 ;
        RECT 63.810 23.110 64.140 23.280 ;
        RECT 64.770 23.110 65.100 23.280 ;
        RECT 65.730 23.110 66.060 23.280 ;
        RECT 66.620 22.770 66.790 28.160 ;
        RECT 61.500 22.600 66.790 22.770 ;
        RECT 70.110 22.420 70.280 28.240 ;
        RECT 70.760 25.600 71.110 27.760 ;
        RECT 70.760 22.900 71.110 25.060 ;
        RECT 71.590 22.420 71.760 28.240 ;
        RECT 72.240 25.600 72.590 27.760 ;
        RECT 72.240 22.900 72.590 25.060 ;
        RECT 73.070 22.420 73.240 28.240 ;
        RECT 73.720 25.600 74.070 27.760 ;
        RECT 73.720 22.900 74.070 25.060 ;
        RECT 74.550 22.420 74.720 28.240 ;
        RECT 75.120 37.540 147.920 37.660 ;
        RECT 75.120 37.490 117.920 37.540 ;
        RECT 75.120 28.000 75.290 37.490 ;
        RECT 75.920 36.980 76.920 37.150 ;
        RECT 75.690 28.725 75.860 36.765 ;
        RECT 76.980 28.725 77.150 36.765 ;
        RECT 75.920 28.340 76.920 28.510 ;
        RECT 77.550 28.000 77.720 37.490 ;
        RECT 78.350 36.980 80.350 37.150 ;
        RECT 78.120 28.725 78.290 36.765 ;
        RECT 80.410 28.725 80.580 36.765 ;
        RECT 78.350 28.340 80.350 28.510 ;
        RECT 80.980 28.000 81.150 37.490 ;
        RECT 81.780 36.980 83.780 37.150 ;
        RECT 81.550 28.725 81.720 36.765 ;
        RECT 83.840 28.725 84.010 36.765 ;
        RECT 81.780 28.340 83.780 28.510 ;
        RECT 84.410 28.000 84.580 37.490 ;
        RECT 85.210 36.980 86.210 37.150 ;
        RECT 84.980 28.725 85.150 36.765 ;
        RECT 86.270 28.725 86.440 36.765 ;
        RECT 86.840 31.890 87.970 37.490 ;
        RECT 85.210 28.340 86.210 28.510 ;
        RECT 86.840 28.000 87.990 31.890 ;
        RECT 75.120 27.830 87.990 28.000 ;
        RECT 90.060 28.000 90.230 37.490 ;
        RECT 90.860 36.980 91.860 37.150 ;
        RECT 90.630 28.725 90.800 36.765 ;
        RECT 91.920 28.725 92.090 36.765 ;
        RECT 90.860 28.340 91.860 28.510 ;
        RECT 92.490 28.000 92.660 37.490 ;
        RECT 93.290 36.980 95.290 37.150 ;
        RECT 93.060 28.725 93.230 36.765 ;
        RECT 95.350 28.725 95.520 36.765 ;
        RECT 93.290 28.340 95.290 28.510 ;
        RECT 95.920 28.000 96.090 37.490 ;
        RECT 96.720 36.980 98.720 37.150 ;
        RECT 96.490 28.725 96.660 36.765 ;
        RECT 98.780 28.725 98.950 36.765 ;
        RECT 96.720 28.340 98.720 28.510 ;
        RECT 99.350 28.000 99.520 37.490 ;
        RECT 101.780 37.480 105.800 37.490 ;
        RECT 100.150 36.980 101.150 37.150 ;
        RECT 99.920 28.725 100.090 36.765 ;
        RECT 101.210 28.725 101.380 36.765 ;
        RECT 101.780 31.890 102.910 37.480 ;
        RECT 100.150 28.340 101.150 28.510 ;
        RECT 101.780 28.000 102.930 31.890 ;
        RECT 90.060 27.830 102.930 28.000 ;
        RECT 105.070 28.000 105.240 37.480 ;
        RECT 105.870 36.980 106.870 37.150 ;
        RECT 105.640 28.725 105.810 36.765 ;
        RECT 106.930 28.725 107.100 36.765 ;
        RECT 105.870 28.340 106.870 28.510 ;
        RECT 107.500 28.000 107.670 37.490 ;
        RECT 108.300 36.980 110.300 37.150 ;
        RECT 108.070 28.725 108.240 36.765 ;
        RECT 110.360 28.725 110.530 36.765 ;
        RECT 108.300 28.340 110.300 28.510 ;
        RECT 110.930 28.000 111.100 37.490 ;
        RECT 111.730 36.980 113.730 37.150 ;
        RECT 111.500 28.725 111.670 36.765 ;
        RECT 113.790 28.725 113.960 36.765 ;
        RECT 111.730 28.340 113.730 28.510 ;
        RECT 114.360 28.000 114.530 37.490 ;
        RECT 115.160 36.980 116.160 37.150 ;
        RECT 114.930 28.725 115.100 36.765 ;
        RECT 116.220 28.725 116.390 36.765 ;
        RECT 116.790 31.890 117.920 37.490 ;
        RECT 120.110 37.490 147.920 37.540 ;
        RECT 115.160 28.340 116.160 28.510 ;
        RECT 116.790 28.000 117.940 31.890 ;
        RECT 105.070 27.830 117.940 28.000 ;
        RECT 120.110 28.000 120.280 37.490 ;
        RECT 120.910 36.980 121.910 37.150 ;
        RECT 120.680 28.725 120.850 36.765 ;
        RECT 121.970 28.725 122.140 36.765 ;
        RECT 120.910 28.340 121.910 28.510 ;
        RECT 122.540 28.000 122.710 37.490 ;
        RECT 123.340 36.980 125.340 37.150 ;
        RECT 123.110 28.725 123.280 36.765 ;
        RECT 125.400 28.725 125.570 36.765 ;
        RECT 123.340 28.340 125.340 28.510 ;
        RECT 125.970 28.000 126.140 37.490 ;
        RECT 126.770 36.980 128.770 37.150 ;
        RECT 126.540 28.725 126.710 36.765 ;
        RECT 128.830 28.725 129.000 36.765 ;
        RECT 126.770 28.340 128.770 28.510 ;
        RECT 129.400 28.000 129.570 37.490 ;
        RECT 131.830 37.480 135.350 37.490 ;
        RECT 130.200 36.980 131.200 37.150 ;
        RECT 129.970 28.725 130.140 36.765 ;
        RECT 131.260 28.725 131.430 36.765 ;
        RECT 131.830 31.890 132.960 37.480 ;
        RECT 130.200 28.340 131.200 28.510 ;
        RECT 131.830 28.000 132.980 31.890 ;
        RECT 120.110 27.830 132.980 28.000 ;
        RECT 135.070 28.000 135.240 37.480 ;
        RECT 135.870 36.980 136.870 37.150 ;
        RECT 135.640 28.725 135.810 36.765 ;
        RECT 136.930 28.725 137.100 36.765 ;
        RECT 135.870 28.340 136.870 28.510 ;
        RECT 137.500 28.000 137.670 37.490 ;
        RECT 138.300 36.980 140.300 37.150 ;
        RECT 138.070 28.725 138.240 36.765 ;
        RECT 140.360 28.725 140.530 36.765 ;
        RECT 138.300 28.340 140.300 28.510 ;
        RECT 140.930 28.000 141.100 37.490 ;
        RECT 141.730 36.980 143.730 37.150 ;
        RECT 141.500 28.725 141.670 36.765 ;
        RECT 143.790 28.725 143.960 36.765 ;
        RECT 141.730 28.340 143.730 28.510 ;
        RECT 144.360 28.000 144.530 37.490 ;
        RECT 145.160 36.980 146.160 37.150 ;
        RECT 144.930 28.725 145.100 36.765 ;
        RECT 146.220 28.725 146.390 36.765 ;
        RECT 146.790 31.890 147.920 37.490 ;
        RECT 145.160 28.340 146.160 28.510 ;
        RECT 146.790 28.000 147.940 31.890 ;
        RECT 135.070 27.830 147.940 28.000 ;
        RECT 86.870 27.800 87.990 27.830 ;
        RECT 101.810 27.800 102.930 27.830 ;
        RECT 116.820 27.800 117.940 27.830 ;
        RECT 131.860 27.800 132.980 27.830 ;
        RECT 146.820 27.800 147.940 27.830 ;
        RECT 86.980 26.580 87.980 27.800 ;
        RECT 101.920 26.580 102.920 27.800 ;
        RECT 116.930 26.580 117.930 27.800 ;
        RECT 131.970 26.580 132.970 27.800 ;
        RECT 146.930 26.580 147.930 27.800 ;
        RECT 86.980 26.510 88.000 26.580 ;
        RECT 101.920 26.510 102.940 26.580 ;
        RECT 116.930 26.510 117.950 26.580 ;
        RECT 131.970 26.510 132.990 26.580 ;
        RECT 146.930 26.510 147.950 26.580 ;
        RECT 84.430 26.240 86.670 26.250 ;
        RECT 70.110 22.250 74.720 22.420 ;
        RECT 75.130 26.080 86.670 26.240 ;
        RECT 75.130 26.070 85.090 26.080 ;
        RECT 61.490 21.710 66.780 21.880 ;
        RECT 61.490 19.310 61.660 21.710 ;
        RECT 62.200 21.200 62.530 21.370 ;
        RECT 62.060 19.990 62.230 21.030 ;
        RECT 62.500 19.990 62.670 21.030 ;
        RECT 62.200 19.650 62.530 19.820 ;
        RECT 63.070 19.310 63.240 21.710 ;
        RECT 64.280 21.200 64.610 21.370 ;
        RECT 65.240 21.200 65.570 21.370 ;
        RECT 63.640 19.990 63.810 21.030 ;
        RECT 64.120 19.990 64.290 21.030 ;
        RECT 64.600 19.990 64.770 21.030 ;
        RECT 65.080 19.990 65.250 21.030 ;
        RECT 65.560 19.990 65.730 21.030 ;
        RECT 66.040 19.990 66.210 21.030 ;
        RECT 63.800 19.650 64.130 19.820 ;
        RECT 64.760 19.650 65.090 19.820 ;
        RECT 65.720 19.650 66.050 19.820 ;
        RECT 66.610 19.310 66.780 21.710 ;
        RECT 75.130 20.680 75.300 26.070 ;
        RECT 75.930 25.560 76.930 25.730 ;
        RECT 75.700 21.350 75.870 25.390 ;
        RECT 76.990 21.350 77.160 25.390 ;
        RECT 75.930 21.010 76.930 21.180 ;
        RECT 77.560 20.680 77.730 26.070 ;
        RECT 78.360 25.560 80.360 25.730 ;
        RECT 78.130 21.350 78.300 25.390 ;
        RECT 80.420 21.350 80.590 25.390 ;
        RECT 78.360 21.010 80.360 21.180 ;
        RECT 80.990 20.680 81.160 26.070 ;
        RECT 81.790 25.560 83.790 25.730 ;
        RECT 81.560 21.350 81.730 25.390 ;
        RECT 83.850 21.350 84.020 25.390 ;
        RECT 84.420 25.170 85.090 26.070 ;
        RECT 85.630 25.570 85.960 25.740 ;
        RECT 84.420 23.990 85.110 25.170 ;
        RECT 85.490 24.360 85.660 25.400 ;
        RECT 85.930 24.360 86.100 25.400 ;
        RECT 86.500 23.990 86.670 26.080 ;
        RECT 86.980 26.050 88.780 26.510 ;
        RECT 99.370 26.240 101.610 26.250 ;
        RECT 84.420 23.820 86.670 23.990 ;
        RECT 87.030 26.010 88.780 26.050 ;
        RECT 84.420 23.660 86.280 23.820 ;
        RECT 84.420 23.430 85.190 23.660 ;
        RECT 84.420 21.920 85.180 23.430 ;
        RECT 81.790 21.010 83.790 21.180 ;
        RECT 84.420 20.720 86.450 21.920 ;
        RECT 87.030 21.880 87.200 26.010 ;
        RECT 87.740 25.505 88.070 25.675 ;
        RECT 88.410 25.300 88.780 26.010 ;
        RECT 87.600 22.250 87.770 25.290 ;
        RECT 88.040 22.250 88.210 25.290 ;
        RECT 88.470 22.330 88.780 25.300 ;
        RECT 88.610 21.880 88.780 22.330 ;
        RECT 87.030 21.710 88.780 21.880 ;
        RECT 90.070 26.080 101.610 26.240 ;
        RECT 90.070 26.070 100.030 26.080 ;
        RECT 90.070 20.720 90.240 26.070 ;
        RECT 90.870 25.560 91.870 25.730 ;
        RECT 90.640 21.350 90.810 25.390 ;
        RECT 91.930 21.350 92.100 25.390 ;
        RECT 90.870 21.010 91.870 21.180 ;
        RECT 84.420 20.680 90.730 20.720 ;
        RECT 92.500 20.680 92.670 26.070 ;
        RECT 93.300 25.560 95.300 25.730 ;
        RECT 93.070 21.350 93.240 25.390 ;
        RECT 95.360 21.350 95.530 25.390 ;
        RECT 93.300 21.010 95.300 21.180 ;
        RECT 95.930 20.680 96.100 26.070 ;
        RECT 96.730 25.560 98.730 25.730 ;
        RECT 96.500 21.350 96.670 25.390 ;
        RECT 98.790 21.350 98.960 25.390 ;
        RECT 99.360 25.170 100.030 26.070 ;
        RECT 100.570 25.570 100.900 25.740 ;
        RECT 99.360 23.990 100.050 25.170 ;
        RECT 100.430 24.360 100.600 25.400 ;
        RECT 100.870 24.360 101.040 25.400 ;
        RECT 101.440 23.990 101.610 26.080 ;
        RECT 101.920 26.050 103.720 26.510 ;
        RECT 114.380 26.240 116.620 26.250 ;
        RECT 99.360 23.820 101.610 23.990 ;
        RECT 101.970 26.010 103.720 26.050 ;
        RECT 99.360 23.660 101.220 23.820 ;
        RECT 99.360 23.430 100.130 23.660 ;
        RECT 99.360 21.920 100.120 23.430 ;
        RECT 96.730 21.010 98.730 21.180 ;
        RECT 99.360 20.730 101.390 21.920 ;
        RECT 101.970 21.880 102.140 26.010 ;
        RECT 102.680 25.505 103.010 25.675 ;
        RECT 103.350 25.300 103.720 26.010 ;
        RECT 102.540 22.250 102.710 25.290 ;
        RECT 102.980 22.250 103.150 25.290 ;
        RECT 103.410 22.330 103.720 25.300 ;
        RECT 103.550 21.880 103.720 22.330 ;
        RECT 101.970 21.710 103.720 21.880 ;
        RECT 105.080 26.080 116.620 26.240 ;
        RECT 105.080 26.070 115.040 26.080 ;
        RECT 105.080 20.730 105.250 26.070 ;
        RECT 105.880 25.560 106.880 25.730 ;
        RECT 105.650 21.350 105.820 25.390 ;
        RECT 106.940 21.350 107.110 25.390 ;
        RECT 105.880 21.010 106.880 21.180 ;
        RECT 99.360 20.680 105.860 20.730 ;
        RECT 107.510 20.680 107.680 26.070 ;
        RECT 108.310 25.560 110.310 25.730 ;
        RECT 108.080 21.350 108.250 25.390 ;
        RECT 110.370 21.350 110.540 25.390 ;
        RECT 108.310 21.010 110.310 21.180 ;
        RECT 110.940 20.680 111.110 26.070 ;
        RECT 111.740 25.560 113.740 25.730 ;
        RECT 111.510 21.350 111.680 25.390 ;
        RECT 113.800 21.350 113.970 25.390 ;
        RECT 114.370 25.170 115.040 26.070 ;
        RECT 115.580 25.570 115.910 25.740 ;
        RECT 114.370 23.990 115.060 25.170 ;
        RECT 115.440 24.360 115.610 25.400 ;
        RECT 115.880 24.360 116.050 25.400 ;
        RECT 116.450 23.990 116.620 26.080 ;
        RECT 116.930 26.050 118.730 26.510 ;
        RECT 129.420 26.240 131.660 26.250 ;
        RECT 114.370 23.820 116.620 23.990 ;
        RECT 116.980 26.010 118.730 26.050 ;
        RECT 114.370 23.660 116.230 23.820 ;
        RECT 114.370 23.430 115.140 23.660 ;
        RECT 114.370 21.920 115.130 23.430 ;
        RECT 111.740 21.010 113.740 21.180 ;
        RECT 114.370 20.730 116.400 21.920 ;
        RECT 116.980 21.880 117.150 26.010 ;
        RECT 117.690 25.505 118.020 25.675 ;
        RECT 118.360 25.300 118.730 26.010 ;
        RECT 117.550 22.250 117.720 25.290 ;
        RECT 117.990 22.250 118.160 25.290 ;
        RECT 118.420 22.330 118.730 25.300 ;
        RECT 118.560 21.880 118.730 22.330 ;
        RECT 116.980 21.710 118.730 21.880 ;
        RECT 120.120 26.080 131.660 26.240 ;
        RECT 120.120 26.070 130.080 26.080 ;
        RECT 120.120 20.730 120.290 26.070 ;
        RECT 120.920 25.560 121.920 25.730 ;
        RECT 120.690 21.350 120.860 25.390 ;
        RECT 121.980 21.350 122.150 25.390 ;
        RECT 120.920 21.010 121.920 21.180 ;
        RECT 114.370 20.680 120.760 20.730 ;
        RECT 122.550 20.680 122.720 26.070 ;
        RECT 123.350 25.560 125.350 25.730 ;
        RECT 123.120 21.350 123.290 25.390 ;
        RECT 125.410 21.350 125.580 25.390 ;
        RECT 123.350 21.010 125.350 21.180 ;
        RECT 125.980 20.680 126.150 26.070 ;
        RECT 126.780 25.560 128.780 25.730 ;
        RECT 126.550 21.350 126.720 25.390 ;
        RECT 128.840 21.350 129.010 25.390 ;
        RECT 129.410 25.170 130.080 26.070 ;
        RECT 130.620 25.570 130.950 25.740 ;
        RECT 129.410 23.990 130.100 25.170 ;
        RECT 130.480 24.360 130.650 25.400 ;
        RECT 130.920 24.360 131.090 25.400 ;
        RECT 131.490 23.990 131.660 26.080 ;
        RECT 131.970 26.050 133.770 26.510 ;
        RECT 144.380 26.240 146.620 26.250 ;
        RECT 129.410 23.820 131.660 23.990 ;
        RECT 132.020 26.010 133.770 26.050 ;
        RECT 129.410 23.660 131.270 23.820 ;
        RECT 129.410 23.430 130.180 23.660 ;
        RECT 129.410 21.920 130.170 23.430 ;
        RECT 126.780 21.010 128.780 21.180 ;
        RECT 129.410 20.680 131.440 21.920 ;
        RECT 132.020 21.880 132.190 26.010 ;
        RECT 132.730 25.505 133.060 25.675 ;
        RECT 133.400 25.300 133.770 26.010 ;
        RECT 132.590 22.250 132.760 25.290 ;
        RECT 133.030 22.250 133.200 25.290 ;
        RECT 133.460 22.330 133.770 25.300 ;
        RECT 133.600 21.880 133.770 22.330 ;
        RECT 132.020 21.710 133.770 21.880 ;
        RECT 135.080 26.080 146.620 26.240 ;
        RECT 135.080 26.070 145.040 26.080 ;
        RECT 75.130 20.670 131.440 20.680 ;
        RECT 135.080 20.680 135.250 26.070 ;
        RECT 135.880 25.560 136.880 25.730 ;
        RECT 135.650 21.350 135.820 25.390 ;
        RECT 136.940 21.350 137.110 25.390 ;
        RECT 135.880 21.010 136.880 21.180 ;
        RECT 137.510 20.680 137.680 26.070 ;
        RECT 138.310 25.560 140.310 25.730 ;
        RECT 138.080 21.350 138.250 25.390 ;
        RECT 140.370 21.350 140.540 25.390 ;
        RECT 138.310 21.010 140.310 21.180 ;
        RECT 140.940 20.680 141.110 26.070 ;
        RECT 141.740 25.560 143.740 25.730 ;
        RECT 141.510 21.350 141.680 25.390 ;
        RECT 143.800 21.350 143.970 25.390 ;
        RECT 144.370 25.170 145.040 26.070 ;
        RECT 145.580 25.570 145.910 25.740 ;
        RECT 144.370 23.990 145.060 25.170 ;
        RECT 145.440 24.360 145.610 25.400 ;
        RECT 145.880 24.360 146.050 25.400 ;
        RECT 146.450 23.990 146.620 26.080 ;
        RECT 146.930 26.050 148.730 26.510 ;
        RECT 144.370 23.820 146.620 23.990 ;
        RECT 146.980 26.010 148.730 26.050 ;
        RECT 144.370 23.660 146.230 23.820 ;
        RECT 144.370 23.430 145.140 23.660 ;
        RECT 144.370 21.920 145.130 23.430 ;
        RECT 141.740 21.010 143.740 21.180 ;
        RECT 144.370 20.680 146.400 21.920 ;
        RECT 146.980 21.880 147.150 26.010 ;
        RECT 147.690 25.505 148.020 25.675 ;
        RECT 148.360 25.300 148.730 26.010 ;
        RECT 147.550 22.250 147.720 25.290 ;
        RECT 147.990 22.250 148.160 25.290 ;
        RECT 148.420 22.330 148.730 25.300 ;
        RECT 148.560 21.880 148.730 22.330 ;
        RECT 146.980 21.710 148.730 21.880 ;
        RECT 135.080 20.670 146.400 20.680 ;
        RECT 75.130 20.500 146.400 20.670 ;
        RECT 75.140 20.010 146.400 20.500 ;
        RECT 84.530 20.000 90.730 20.010 ;
        RECT 99.470 20.000 105.860 20.010 ;
        RECT 114.480 20.000 120.760 20.010 ;
        RECT 129.520 20.000 135.840 20.010 ;
        RECT 144.480 20.000 146.400 20.010 ;
        RECT 85.900 19.990 90.730 20.000 ;
        RECT 131.010 19.940 135.840 20.000 ;
        RECT 61.490 19.140 66.780 19.310 ;
        RECT 61.500 18.310 66.780 19.140 ;
      LAYER met1 ;
        RECT 33.300 224.810 33.870 225.380 ;
        RECT 74.640 224.940 75.350 225.590 ;
        RECT 12.330 223.740 12.470 223.910 ;
        RECT 74.910 223.740 75.050 224.940 ;
        RECT 77.450 224.860 78.030 225.470 ;
        RECT 80.190 224.880 80.730 225.500 ;
        RECT 88.520 225.060 89.040 225.620 ;
        RECT 12.330 223.600 75.050 223.740 ;
        RECT 12.330 128.470 12.470 223.600 ;
        RECT 77.615 223.370 77.840 224.860 ;
        RECT 13.830 223.245 14.090 223.260 ;
        RECT 16.825 223.245 77.840 223.370 ;
        RECT 13.830 223.145 77.840 223.245 ;
        RECT 13.830 223.070 17.050 223.145 ;
        RECT 13.830 145.050 14.090 223.070 ;
        RECT 80.380 222.895 80.535 224.880 ;
        RECT 14.435 222.740 80.535 222.895 ;
        RECT 14.435 149.220 14.590 222.740 ;
        RECT 88.690 222.585 88.895 225.060 ;
        RECT 91.220 224.940 91.850 225.620 ;
        RECT 15.035 222.380 88.895 222.585 ;
        RECT 15.035 203.870 15.190 222.380 ;
        RECT 91.440 222.240 91.580 224.940 ;
        RECT 93.980 224.910 94.550 225.440 ;
        RECT 137.980 224.970 138.430 225.420 ;
        RECT 15.400 222.100 91.580 222.240 ;
        RECT 94.225 222.250 94.375 224.910 ;
        RECT 125.800 224.280 126.280 224.400 ;
        RECT 136.550 224.280 137.150 224.410 ;
        RECT 125.800 224.085 137.150 224.280 ;
        RECT 125.800 223.980 126.280 224.085 ;
        RECT 136.550 223.930 137.150 224.085 ;
        RECT 95.960 222.250 96.290 222.270 ;
        RECT 94.225 222.100 96.290 222.250 ;
        RECT 14.990 177.720 15.230 203.870 ;
        RECT 12.940 144.895 14.120 145.050 ;
        RECT 12.935 144.730 14.120 144.895 ;
        RECT 12.935 141.070 13.270 144.730 ;
        RECT 13.500 144.405 14.200 144.420 ;
        RECT 14.350 144.405 14.670 149.220 ;
        RECT 13.500 143.930 14.670 144.405 ;
        RECT 13.500 143.775 14.465 143.930 ;
        RECT 13.500 143.750 14.200 143.775 ;
        RECT 12.935 140.525 14.220 141.070 ;
        RECT 13.150 140.350 14.220 140.525 ;
        RECT 12.330 128.330 14.790 128.470 ;
        RECT 14.650 122.610 14.790 128.330 ;
        RECT 14.970 124.320 15.250 177.720 ;
        RECT 15.400 128.010 15.540 222.100 ;
        RECT 95.960 221.950 96.290 222.100 ;
        RECT 138.140 221.790 138.280 224.970 ;
        RECT 16.840 221.650 138.280 221.790 ;
        RECT 15.960 163.030 16.280 163.090 ;
        RECT 16.840 163.030 16.980 221.650 ;
        RECT 17.270 221.030 146.990 221.510 ;
        RECT 79.440 220.490 79.760 220.550 ;
        RECT 80.375 220.490 80.665 220.535 ;
        RECT 79.440 220.350 80.665 220.490 ;
        RECT 79.440 220.290 79.760 220.350 ;
        RECT 80.375 220.305 80.665 220.350 ;
        RECT 84.055 220.490 84.345 220.535 ;
        RECT 87.720 220.490 88.040 220.550 ;
        RECT 84.055 220.350 88.040 220.490 ;
        RECT 84.055 220.305 84.345 220.350 ;
        RECT 87.720 220.290 88.040 220.350 ;
        RECT 95.540 220.490 95.860 220.550 ;
        RECT 96.475 220.490 96.765 220.535 ;
        RECT 95.540 220.350 96.765 220.490 ;
        RECT 95.540 220.290 95.860 220.350 ;
        RECT 96.475 220.305 96.765 220.350 ;
        RECT 85.880 220.150 86.200 220.210 ;
        RECT 85.880 220.010 87.950 220.150 ;
        RECT 85.880 219.950 86.200 220.010 ;
        RECT 60.120 219.810 60.440 219.870 ;
        RECT 60.595 219.810 60.885 219.855 ;
        RECT 60.120 219.670 60.885 219.810 ;
        RECT 60.120 219.610 60.440 219.670 ;
        RECT 60.595 219.625 60.885 219.670 ;
        RECT 81.295 219.625 81.585 219.855 ;
        RECT 82.660 219.810 82.980 219.870 ;
        RECT 83.135 219.810 83.425 219.855 ;
        RECT 82.660 219.670 83.425 219.810 ;
        RECT 51.840 219.470 52.160 219.530 ;
        RECT 61.975 219.470 62.265 219.515 ;
        RECT 51.840 219.330 62.265 219.470 ;
        RECT 81.370 219.470 81.510 219.625 ;
        RECT 82.660 219.610 82.980 219.670 ;
        RECT 83.135 219.625 83.425 219.670 ;
        RECT 86.355 219.625 86.645 219.855 ;
        RECT 84.500 219.470 84.820 219.530 ;
        RECT 81.370 219.330 84.820 219.470 ;
        RECT 86.430 219.470 86.570 219.625 ;
        RECT 87.260 219.610 87.580 219.870 ;
        RECT 87.810 219.855 87.950 220.010 ;
        RECT 87.735 219.625 88.025 219.855 ;
        RECT 89.100 219.810 89.420 219.870 ;
        RECT 90.495 219.810 90.785 219.855 ;
        RECT 89.100 219.670 90.785 219.810 ;
        RECT 89.100 219.610 89.420 219.670 ;
        RECT 90.495 219.625 90.785 219.670 ;
        RECT 97.395 219.810 97.685 219.855 ;
        RECT 103.360 219.810 103.680 219.870 ;
        RECT 97.395 219.670 103.680 219.810 ;
        RECT 97.395 219.625 97.685 219.670 ;
        RECT 103.360 219.610 103.680 219.670 ;
        RECT 89.560 219.470 89.880 219.530 ;
        RECT 86.430 219.330 89.880 219.470 ;
        RECT 51.840 219.270 52.160 219.330 ;
        RECT 61.975 219.285 62.265 219.330 ;
        RECT 84.500 219.270 84.820 219.330 ;
        RECT 89.560 219.270 89.880 219.330 ;
        RECT 85.420 218.930 85.740 219.190 ;
        RECT 88.180 219.130 88.500 219.190 ;
        RECT 88.655 219.130 88.945 219.175 ;
        RECT 88.180 218.990 88.945 219.130 ;
        RECT 88.180 218.930 88.500 218.990 ;
        RECT 88.655 218.945 88.945 218.990 ;
        RECT 90.940 218.930 91.260 219.190 ;
        RECT 17.270 218.310 146.990 218.790 ;
        RECT 55.060 218.110 55.380 218.170 ;
        RECT 55.060 217.970 70.470 218.110 ;
        RECT 55.060 217.910 55.380 217.970 ;
        RECT 60.135 217.770 60.425 217.815 ;
        RECT 64.260 217.770 64.580 217.830 ;
        RECT 67.495 217.770 67.785 217.815 ;
        RECT 53.310 217.630 58.510 217.770 ;
        RECT 53.310 217.475 53.450 217.630 ;
        RECT 53.235 217.245 53.525 217.475 ;
        RECT 53.680 217.230 54.000 217.490 ;
        RECT 54.155 217.430 54.445 217.475 ;
        RECT 55.060 217.430 55.380 217.490 ;
        RECT 54.155 217.290 55.380 217.430 ;
        RECT 54.155 217.245 54.445 217.290 ;
        RECT 55.060 217.230 55.380 217.290 ;
        RECT 55.535 217.430 55.825 217.475 ;
        RECT 58.370 217.430 58.510 217.630 ;
        RECT 60.135 217.630 61.730 217.770 ;
        RECT 60.135 217.585 60.425 217.630 ;
        RECT 60.580 217.430 60.900 217.490 ;
        RECT 61.590 217.475 61.730 217.630 ;
        RECT 64.260 217.630 67.785 217.770 ;
        RECT 64.260 217.570 64.580 217.630 ;
        RECT 67.495 217.585 67.785 217.630 ;
        RECT 55.535 217.290 58.050 217.430 ;
        RECT 58.370 217.290 60.900 217.430 ;
        RECT 55.535 217.245 55.825 217.290 ;
        RECT 52.300 216.890 52.620 217.150 ;
        RECT 56.900 216.890 57.220 217.150 ;
        RECT 57.910 217.090 58.050 217.290 ;
        RECT 60.580 217.230 60.900 217.290 ;
        RECT 61.515 217.245 61.805 217.475 ;
        RECT 67.035 217.245 67.325 217.475 ;
        RECT 61.055 217.090 61.345 217.135 ;
        RECT 57.910 216.950 61.345 217.090 ;
        RECT 61.055 216.905 61.345 216.950 ;
        RECT 55.075 216.750 55.365 216.795 ;
        RECT 60.120 216.750 60.440 216.810 ;
        RECT 67.110 216.750 67.250 217.245 ;
        RECT 68.400 217.230 68.720 217.490 ;
        RECT 68.860 217.430 69.180 217.490 ;
        RECT 70.330 217.475 70.470 217.970 ;
        RECT 89.100 217.910 89.420 218.170 ;
        RECT 89.560 217.910 89.880 218.170 ;
        RECT 93.240 218.110 93.560 218.170 ;
        RECT 90.110 217.970 93.560 218.110 ;
        RECT 69.335 217.430 69.625 217.475 ;
        RECT 68.860 217.290 69.625 217.430 ;
        RECT 68.860 217.230 69.180 217.290 ;
        RECT 69.335 217.245 69.625 217.290 ;
        RECT 70.255 217.430 70.545 217.475 ;
        RECT 70.700 217.430 71.020 217.490 ;
        RECT 70.255 217.290 71.020 217.430 ;
        RECT 70.255 217.245 70.545 217.290 ;
        RECT 70.700 217.230 71.020 217.290 ;
        RECT 81.295 217.090 81.585 217.135 ;
        RECT 82.660 217.090 82.980 217.150 ;
        RECT 81.295 216.950 82.980 217.090 ;
        RECT 81.295 216.905 81.585 216.950 ;
        RECT 82.660 216.890 82.980 216.950 ;
        RECT 85.880 217.090 86.200 217.150 ;
        RECT 90.110 217.090 90.250 217.970 ;
        RECT 93.240 217.910 93.560 217.970 ;
        RECT 97.855 217.925 98.145 218.155 ;
        RECT 90.480 217.770 90.800 217.830 ;
        RECT 95.540 217.770 95.860 217.830 ;
        RECT 96.935 217.770 97.225 217.815 ;
        RECT 90.480 217.630 91.195 217.770 ;
        RECT 90.480 217.570 90.800 217.630 ;
        RECT 91.055 217.475 91.195 217.630 ;
        RECT 91.950 217.630 97.225 217.770 ;
        RECT 90.955 217.245 91.245 217.475 ;
        RECT 91.950 217.420 92.090 217.630 ;
        RECT 95.540 217.570 95.860 217.630 ;
        RECT 96.935 217.585 97.225 217.630 ;
        RECT 97.380 217.770 97.700 217.830 ;
        RECT 97.930 217.770 98.070 217.925 ;
        RECT 102.455 217.770 102.745 217.815 ;
        RECT 97.380 217.630 102.745 217.770 ;
        RECT 91.490 217.280 92.090 217.420 ;
        RECT 91.490 217.135 91.630 217.280 ;
        RECT 93.240 217.230 93.560 217.490 ;
        RECT 94.175 217.430 94.465 217.475 ;
        RECT 96.460 217.430 96.780 217.490 ;
        RECT 94.175 217.290 96.780 217.430 ;
        RECT 97.010 217.430 97.150 217.585 ;
        RECT 97.380 217.570 97.700 217.630 ;
        RECT 102.455 217.585 102.745 217.630 ;
        RECT 103.360 217.570 103.680 217.830 ;
        RECT 100.155 217.430 100.445 217.475 ;
        RECT 97.010 217.290 100.445 217.430 ;
        RECT 94.175 217.245 94.465 217.290 ;
        RECT 96.460 217.230 96.780 217.290 ;
        RECT 100.155 217.245 100.445 217.290 ;
        RECT 90.495 217.090 90.785 217.135 ;
        RECT 85.880 216.950 90.785 217.090 ;
        RECT 85.880 216.890 86.200 216.950 ;
        RECT 90.495 216.905 90.785 216.950 ;
        RECT 91.415 216.905 91.705 217.135 ;
        RECT 91.875 216.905 92.165 217.135 ;
        RECT 93.715 217.090 94.005 217.135 ;
        RECT 98.760 217.090 99.080 217.150 ;
        RECT 99.695 217.090 99.985 217.135 ;
        RECT 93.715 216.950 99.985 217.090 ;
        RECT 93.715 216.905 94.005 216.950 ;
        RECT 91.950 216.750 92.090 216.905 ;
        RECT 98.760 216.890 99.080 216.950 ;
        RECT 99.695 216.905 99.985 216.950 ;
        RECT 55.075 216.610 67.250 216.750 ;
        RECT 91.030 216.610 92.090 216.750 ;
        RECT 95.095 216.750 95.385 216.795 ;
        RECT 96.460 216.750 96.780 216.810 ;
        RECT 95.095 216.610 96.780 216.750 ;
        RECT 55.075 216.565 55.365 216.610 ;
        RECT 60.120 216.550 60.440 216.610 ;
        RECT 53.695 216.410 53.985 216.455 ;
        RECT 54.140 216.410 54.460 216.470 ;
        RECT 53.695 216.270 54.460 216.410 ;
        RECT 53.695 216.225 53.985 216.270 ;
        RECT 54.140 216.210 54.460 216.270 ;
        RECT 55.520 216.210 55.840 216.470 ;
        RECT 65.180 216.410 65.500 216.470 ;
        RECT 68.415 216.410 68.705 216.455 ;
        RECT 65.180 216.270 68.705 216.410 ;
        RECT 65.180 216.210 65.500 216.270 ;
        RECT 68.415 216.225 68.705 216.270 ;
        RECT 69.320 216.210 69.640 216.470 ;
        RECT 71.620 216.410 71.940 216.470 ;
        RECT 84.055 216.410 84.345 216.455 ;
        RECT 91.030 216.410 91.170 216.610 ;
        RECT 95.095 216.565 95.385 216.610 ;
        RECT 96.460 216.550 96.780 216.610 ;
        RECT 101.995 216.750 102.285 216.795 ;
        RECT 106.580 216.750 106.900 216.810 ;
        RECT 101.995 216.610 106.900 216.750 ;
        RECT 101.995 216.565 102.285 216.610 ;
        RECT 106.580 216.550 106.900 216.610 ;
        RECT 71.620 216.270 91.170 216.410 ;
        RECT 93.240 216.410 93.560 216.470 ;
        RECT 96.935 216.410 97.225 216.455 ;
        RECT 93.240 216.270 97.225 216.410 ;
        RECT 71.620 216.210 71.940 216.270 ;
        RECT 84.055 216.225 84.345 216.270 ;
        RECT 93.240 216.210 93.560 216.270 ;
        RECT 96.935 216.225 97.225 216.270 ;
        RECT 104.280 216.210 104.600 216.470 ;
        RECT 17.270 215.590 146.990 216.070 ;
        RECT 56.455 215.390 56.745 215.435 ;
        RECT 56.900 215.390 57.220 215.450 ;
        RECT 56.455 215.250 57.220 215.390 ;
        RECT 56.455 215.205 56.745 215.250 ;
        RECT 56.900 215.190 57.220 215.250 ;
        RECT 89.560 215.390 89.880 215.450 ;
        RECT 97.380 215.390 97.700 215.450 ;
        RECT 89.560 215.250 97.700 215.390 ;
        RECT 89.560 215.190 89.880 215.250 ;
        RECT 97.380 215.190 97.700 215.250 ;
        RECT 103.360 215.390 103.680 215.450 ;
        RECT 104.295 215.390 104.585 215.435 ;
        RECT 103.360 215.250 104.585 215.390 ;
        RECT 103.360 215.190 103.680 215.250 ;
        RECT 104.295 215.205 104.585 215.250 ;
        RECT 50.920 215.050 51.240 215.110 ;
        RECT 52.775 215.050 53.065 215.095 ;
        RECT 50.920 214.910 53.065 215.050 ;
        RECT 50.920 214.850 51.240 214.910 ;
        RECT 52.775 214.865 53.065 214.910 ;
        RECT 59.200 215.050 59.490 215.095 ;
        RECT 60.770 215.050 61.060 215.095 ;
        RECT 62.870 215.050 63.160 215.095 ;
        RECT 59.200 214.910 63.160 215.050 ;
        RECT 59.200 214.865 59.490 214.910 ;
        RECT 60.770 214.865 61.060 214.910 ;
        RECT 62.870 214.865 63.160 214.910 ;
        RECT 67.020 215.050 67.310 215.095 ;
        RECT 68.590 215.050 68.880 215.095 ;
        RECT 70.690 215.050 70.980 215.095 ;
        RECT 67.020 214.910 70.980 215.050 ;
        RECT 67.020 214.865 67.310 214.910 ;
        RECT 68.590 214.865 68.880 214.910 ;
        RECT 70.690 214.865 70.980 214.910 ;
        RECT 85.420 215.050 85.710 215.095 ;
        RECT 86.990 215.050 87.280 215.095 ;
        RECT 89.090 215.050 89.380 215.095 ;
        RECT 85.420 214.910 89.380 215.050 ;
        RECT 85.420 214.865 85.710 214.910 ;
        RECT 86.990 214.865 87.280 214.910 ;
        RECT 89.090 214.865 89.380 214.910 ;
        RECT 90.520 215.050 90.810 215.095 ;
        RECT 92.620 215.050 92.910 215.095 ;
        RECT 94.190 215.050 94.480 215.095 ;
        RECT 90.520 214.910 94.480 215.050 ;
        RECT 90.520 214.865 90.810 214.910 ;
        RECT 92.620 214.865 92.910 214.910 ;
        RECT 94.190 214.865 94.480 214.910 ;
        RECT 97.880 215.050 98.170 215.095 ;
        RECT 99.980 215.050 100.270 215.095 ;
        RECT 101.550 215.050 101.840 215.095 ;
        RECT 97.880 214.910 101.840 215.050 ;
        RECT 97.880 214.865 98.170 214.910 ;
        RECT 99.980 214.865 100.270 214.910 ;
        RECT 101.550 214.865 101.840 214.910 ;
        RECT 53.220 214.710 53.540 214.770 ;
        RECT 54.155 214.710 54.445 214.755 ;
        RECT 53.220 214.570 54.445 214.710 ;
        RECT 53.220 214.510 53.540 214.570 ;
        RECT 54.155 214.525 54.445 214.570 ;
        RECT 58.765 214.710 59.055 214.755 ;
        RECT 61.285 214.710 61.575 214.755 ;
        RECT 62.475 214.710 62.765 214.755 ;
        RECT 58.765 214.570 62.765 214.710 ;
        RECT 58.765 214.525 59.055 214.570 ;
        RECT 61.285 214.525 61.575 214.570 ;
        RECT 62.475 214.525 62.765 214.570 ;
        RECT 66.585 214.710 66.875 214.755 ;
        RECT 69.105 214.710 69.395 214.755 ;
        RECT 70.295 214.710 70.585 214.755 ;
        RECT 66.585 214.570 70.585 214.710 ;
        RECT 66.585 214.525 66.875 214.570 ;
        RECT 69.105 214.525 69.395 214.570 ;
        RECT 70.295 214.525 70.585 214.570 ;
        RECT 84.985 214.710 85.275 214.755 ;
        RECT 87.505 214.710 87.795 214.755 ;
        RECT 88.695 214.710 88.985 214.755 ;
        RECT 84.985 214.570 88.985 214.710 ;
        RECT 84.985 214.525 85.275 214.570 ;
        RECT 87.505 214.525 87.795 214.570 ;
        RECT 88.695 214.525 88.985 214.570 ;
        RECT 90.915 214.710 91.205 214.755 ;
        RECT 92.105 214.710 92.395 214.755 ;
        RECT 94.625 214.710 94.915 214.755 ;
        RECT 90.915 214.570 94.915 214.710 ;
        RECT 90.915 214.525 91.205 214.570 ;
        RECT 92.105 214.525 92.395 214.570 ;
        RECT 94.625 214.525 94.915 214.570 ;
        RECT 98.275 214.710 98.565 214.755 ;
        RECT 99.465 214.710 99.755 214.755 ;
        RECT 101.985 214.710 102.275 214.755 ;
        RECT 98.275 214.570 102.275 214.710 ;
        RECT 98.275 214.525 98.565 214.570 ;
        RECT 99.465 214.525 99.755 214.570 ;
        RECT 101.985 214.525 102.275 214.570 ;
        RECT 52.315 214.370 52.605 214.415 ;
        RECT 54.600 214.370 54.920 214.430 ;
        RECT 52.315 214.230 54.920 214.370 ;
        RECT 52.315 214.185 52.605 214.230 ;
        RECT 54.600 214.170 54.920 214.230 ;
        RECT 55.520 214.370 55.840 214.430 ;
        RECT 62.020 214.370 62.310 214.415 ;
        RECT 55.520 214.230 62.310 214.370 ;
        RECT 55.520 214.170 55.840 214.230 ;
        RECT 62.020 214.185 62.310 214.230 ;
        RECT 63.355 214.370 63.645 214.415 ;
        RECT 65.640 214.370 65.960 214.430 ;
        RECT 71.175 214.370 71.465 214.415 ;
        RECT 89.575 214.370 89.865 214.415 ;
        RECT 90.035 214.370 90.325 214.415 ;
        RECT 63.355 214.230 71.465 214.370 ;
        RECT 63.355 214.185 63.645 214.230 ;
        RECT 65.640 214.170 65.960 214.230 ;
        RECT 71.175 214.185 71.465 214.230 ;
        RECT 80.450 214.230 90.325 214.370 ;
        RECT 69.320 214.030 69.640 214.090 ;
        RECT 69.840 214.030 70.130 214.075 ;
        RECT 69.320 213.890 70.130 214.030 ;
        RECT 69.320 213.830 69.640 213.890 ;
        RECT 69.840 213.845 70.130 213.890 ;
        RECT 80.450 213.750 80.590 214.230 ;
        RECT 89.575 214.185 89.865 214.230 ;
        RECT 90.035 214.185 90.325 214.230 ;
        RECT 96.460 214.370 96.780 214.430 ;
        RECT 97.395 214.370 97.685 214.415 ;
        RECT 96.460 214.230 97.685 214.370 ;
        RECT 96.460 214.170 96.780 214.230 ;
        RECT 97.395 214.185 97.685 214.230 ;
        RECT 85.420 214.030 85.740 214.090 ;
        RECT 88.240 214.030 88.530 214.075 ;
        RECT 85.420 213.890 88.530 214.030 ;
        RECT 85.420 213.830 85.740 213.890 ;
        RECT 88.240 213.845 88.530 213.890 ;
        RECT 91.370 214.030 91.660 214.075 ;
        RECT 91.860 214.030 92.180 214.090 ;
        RECT 91.370 213.890 92.180 214.030 ;
        RECT 91.370 213.845 91.660 213.890 ;
        RECT 91.860 213.830 92.180 213.890 ;
        RECT 98.730 214.030 99.020 214.075 ;
        RECT 100.600 214.030 100.920 214.090 ;
        RECT 98.730 213.890 100.920 214.030 ;
        RECT 98.730 213.845 99.020 213.890 ;
        RECT 100.600 213.830 100.920 213.890 ;
        RECT 103.360 214.030 103.680 214.090 ;
        RECT 104.755 214.030 105.045 214.075 ;
        RECT 103.360 213.890 105.045 214.030 ;
        RECT 103.360 213.830 103.680 213.890 ;
        RECT 104.755 213.845 105.045 213.890 ;
        RECT 106.595 214.030 106.885 214.075 ;
        RECT 107.040 214.030 107.360 214.090 ;
        RECT 106.595 213.890 107.360 214.030 ;
        RECT 106.595 213.845 106.885 213.890 ;
        RECT 107.040 213.830 107.360 213.890 ;
        RECT 49.080 213.490 49.400 213.750 ;
        RECT 64.260 213.490 64.580 213.750 ;
        RECT 80.360 213.490 80.680 213.750 ;
        RECT 82.660 213.490 82.980 213.750 ;
        RECT 96.920 213.490 97.240 213.750 ;
        RECT 17.270 212.870 146.990 213.350 ;
        RECT 49.080 212.670 49.400 212.730 ;
        RECT 45.030 212.530 49.400 212.670 ;
        RECT 45.030 212.035 45.170 212.530 ;
        RECT 49.080 212.470 49.400 212.530 ;
        RECT 68.400 212.470 68.720 212.730 ;
        RECT 79.915 212.670 80.205 212.715 ;
        RECT 85.880 212.670 86.200 212.730 ;
        RECT 79.915 212.530 86.200 212.670 ;
        RECT 79.915 212.485 80.205 212.530 ;
        RECT 85.880 212.470 86.200 212.530 ;
        RECT 87.260 212.670 87.580 212.730 ;
        RECT 87.260 212.530 90.710 212.670 ;
        RECT 87.260 212.470 87.580 212.530 ;
        RECT 45.400 212.330 45.720 212.390 ;
        RECT 86.340 212.330 86.660 212.390 ;
        RECT 90.035 212.330 90.325 212.375 ;
        RECT 45.400 212.190 53.910 212.330 ;
        RECT 45.400 212.130 45.720 212.190 ;
        RECT 46.410 212.035 46.550 212.190 ;
        RECT 44.955 211.805 45.245 212.035 ;
        RECT 45.875 211.805 46.165 212.035 ;
        RECT 46.335 211.805 46.625 212.035 ;
        RECT 47.670 211.990 47.960 212.035 ;
        RECT 50.460 211.990 50.780 212.050 ;
        RECT 53.770 212.035 53.910 212.190 ;
        RECT 72.170 212.190 80.590 212.330 ;
        RECT 47.670 211.850 50.780 211.990 ;
        RECT 47.670 211.805 47.960 211.850 ;
        RECT 45.950 211.310 46.090 211.805 ;
        RECT 50.460 211.790 50.780 211.850 ;
        RECT 53.695 211.805 53.985 212.035 ;
        RECT 54.140 211.990 54.460 212.050 ;
        RECT 54.975 211.990 55.265 212.035 ;
        RECT 54.140 211.850 55.265 211.990 ;
        RECT 54.140 211.790 54.460 211.850 ;
        RECT 54.975 211.805 55.265 211.850 ;
        RECT 65.195 211.990 65.485 212.035 ;
        RECT 66.100 211.990 66.420 212.050 ;
        RECT 65.195 211.850 66.420 211.990 ;
        RECT 65.195 211.805 65.485 211.850 ;
        RECT 66.100 211.790 66.420 211.850 ;
        RECT 69.320 211.790 69.640 212.050 ;
        RECT 70.255 211.990 70.545 212.035 ;
        RECT 71.160 211.990 71.480 212.050 ;
        RECT 70.255 211.850 71.480 211.990 ;
        RECT 70.255 211.805 70.545 211.850 ;
        RECT 71.160 211.790 71.480 211.850 ;
        RECT 71.620 211.790 71.940 212.050 ;
        RECT 47.215 211.650 47.505 211.695 ;
        RECT 48.405 211.650 48.695 211.695 ;
        RECT 50.925 211.650 51.215 211.695 ;
        RECT 47.215 211.510 51.215 211.650 ;
        RECT 47.215 211.465 47.505 211.510 ;
        RECT 48.405 211.465 48.695 211.510 ;
        RECT 50.925 211.465 51.215 211.510 ;
        RECT 54.575 211.650 54.865 211.695 ;
        RECT 55.765 211.650 56.055 211.695 ;
        RECT 58.285 211.650 58.575 211.695 ;
        RECT 63.815 211.650 64.105 211.695 ;
        RECT 54.575 211.510 58.575 211.650 ;
        RECT 54.575 211.465 54.865 211.510 ;
        RECT 55.765 211.465 56.055 211.510 ;
        RECT 58.285 211.465 58.575 211.510 ;
        RECT 60.670 211.510 64.105 211.650 ;
        RECT 46.820 211.310 47.110 211.355 ;
        RECT 48.920 211.310 49.210 211.355 ;
        RECT 50.490 211.310 50.780 211.355 ;
        RECT 54.180 211.310 54.470 211.355 ;
        RECT 56.280 211.310 56.570 211.355 ;
        RECT 57.850 211.310 58.140 211.355 ;
        RECT 45.950 211.170 46.550 211.310 ;
        RECT 45.860 210.770 46.180 211.030 ;
        RECT 46.410 210.970 46.550 211.170 ;
        RECT 46.820 211.170 50.780 211.310 ;
        RECT 46.820 211.125 47.110 211.170 ;
        RECT 48.920 211.125 49.210 211.170 ;
        RECT 50.490 211.125 50.780 211.170 ;
        RECT 52.850 211.170 53.910 211.310 ;
        RECT 52.850 210.970 52.990 211.170 ;
        RECT 46.410 210.830 52.990 210.970 ;
        RECT 53.220 210.770 53.540 211.030 ;
        RECT 53.770 210.970 53.910 211.170 ;
        RECT 54.180 211.170 58.140 211.310 ;
        RECT 54.180 211.125 54.470 211.170 ;
        RECT 56.280 211.125 56.570 211.170 ;
        RECT 57.850 211.125 58.140 211.170 ;
        RECT 59.660 211.310 59.980 211.370 ;
        RECT 60.670 211.355 60.810 211.510 ;
        RECT 63.815 211.465 64.105 211.510 ;
        RECT 65.640 211.650 65.960 211.710 ;
        RECT 72.170 211.650 72.310 212.190 ;
        RECT 80.450 212.050 80.590 212.190 ;
        RECT 86.340 212.190 90.325 212.330 ;
        RECT 90.570 212.330 90.710 212.530 ;
        RECT 91.860 212.470 92.180 212.730 ;
        RECT 96.935 212.670 97.225 212.715 ;
        RECT 107.040 212.670 107.360 212.730 ;
        RECT 96.935 212.530 107.360 212.670 ;
        RECT 96.935 212.485 97.225 212.530 ;
        RECT 107.040 212.470 107.360 212.530 ;
        RECT 96.460 212.330 96.780 212.390 ;
        RECT 90.570 212.190 92.550 212.330 ;
        RECT 86.340 212.130 86.660 212.190 ;
        RECT 90.035 212.145 90.325 212.190 ;
        RECT 92.410 212.050 92.550 212.190 ;
        RECT 96.460 212.190 108.190 212.330 ;
        RECT 96.460 212.130 96.780 212.190 ;
        RECT 72.555 212.020 72.845 212.035 ;
        RECT 72.555 211.990 73.690 212.020 ;
        RECT 74.295 211.990 74.585 212.035 ;
        RECT 72.555 211.880 74.585 211.990 ;
        RECT 72.555 211.805 72.845 211.880 ;
        RECT 73.550 211.850 74.585 211.880 ;
        RECT 74.295 211.805 74.585 211.850 ;
        RECT 80.360 211.790 80.680 212.050 ;
        RECT 81.740 212.035 82.060 212.050 ;
        RECT 89.560 212.035 89.880 212.050 ;
        RECT 81.710 211.805 82.060 212.035 ;
        RECT 88.655 211.805 88.945 212.035 ;
        RECT 89.395 211.805 89.880 212.035 ;
        RECT 81.740 211.790 82.060 211.805 ;
        RECT 73.015 211.650 73.305 211.695 ;
        RECT 65.640 211.510 73.305 211.650 ;
        RECT 65.640 211.450 65.960 211.510 ;
        RECT 73.015 211.465 73.305 211.510 ;
        RECT 73.895 211.650 74.185 211.695 ;
        RECT 75.085 211.650 75.375 211.695 ;
        RECT 77.605 211.650 77.895 211.695 ;
        RECT 73.895 211.510 77.895 211.650 ;
        RECT 73.895 211.465 74.185 211.510 ;
        RECT 75.085 211.465 75.375 211.510 ;
        RECT 77.605 211.465 77.895 211.510 ;
        RECT 81.255 211.650 81.545 211.695 ;
        RECT 82.445 211.650 82.735 211.695 ;
        RECT 84.965 211.650 85.255 211.695 ;
        RECT 81.255 211.510 85.255 211.650 ;
        RECT 88.730 211.650 88.870 211.805 ;
        RECT 89.560 211.790 89.880 211.805 ;
        RECT 90.480 211.790 90.800 212.050 ;
        RECT 90.940 212.035 91.260 212.050 ;
        RECT 90.940 211.990 91.270 212.035 ;
        RECT 92.320 211.990 92.640 212.050 ;
        RECT 93.255 211.990 93.545 212.035 ;
        RECT 90.940 211.850 91.455 211.990 ;
        RECT 92.320 211.850 93.545 211.990 ;
        RECT 90.940 211.805 91.270 211.850 ;
        RECT 90.940 211.790 91.260 211.805 ;
        RECT 92.320 211.790 92.640 211.850 ;
        RECT 93.255 211.805 93.545 211.850 ;
        RECT 95.095 211.990 95.385 212.035 ;
        RECT 97.380 211.990 97.700 212.050 ;
        RECT 95.095 211.850 97.700 211.990 ;
        RECT 95.095 211.805 95.385 211.850 ;
        RECT 97.380 211.790 97.700 211.850 ;
        RECT 98.760 211.790 99.080 212.050 ;
        RECT 100.615 211.990 100.905 212.035 ;
        RECT 104.280 211.990 104.600 212.050 ;
        RECT 100.615 211.850 104.600 211.990 ;
        RECT 100.615 211.805 100.905 211.850 ;
        RECT 104.280 211.790 104.600 211.850 ;
        RECT 106.580 212.035 106.900 212.050 ;
        RECT 108.050 212.035 108.190 212.190 ;
        RECT 106.580 211.990 106.930 212.035 ;
        RECT 106.580 211.850 107.095 211.990 ;
        RECT 106.580 211.805 106.930 211.850 ;
        RECT 107.975 211.805 108.265 212.035 ;
        RECT 106.580 211.790 106.900 211.805 ;
        RECT 92.795 211.650 93.085 211.695 ;
        RECT 88.730 211.510 93.085 211.650 ;
        RECT 81.255 211.465 81.545 211.510 ;
        RECT 82.445 211.465 82.735 211.510 ;
        RECT 84.965 211.465 85.255 211.510 ;
        RECT 92.795 211.465 93.085 211.510 ;
        RECT 95.540 211.650 95.860 211.710 ;
        RECT 98.315 211.650 98.605 211.695 ;
        RECT 95.540 211.510 98.605 211.650 ;
        RECT 95.540 211.450 95.860 211.510 ;
        RECT 98.315 211.465 98.605 211.510 ;
        RECT 100.155 211.650 100.445 211.695 ;
        RECT 102.900 211.650 103.220 211.710 ;
        RECT 100.155 211.510 103.220 211.650 ;
        RECT 100.155 211.465 100.445 211.510 ;
        RECT 60.595 211.310 60.885 211.355 ;
        RECT 59.660 211.170 60.885 211.310 ;
        RECT 59.660 211.110 59.980 211.170 ;
        RECT 60.595 211.125 60.885 211.170 ;
        RECT 73.500 211.310 73.790 211.355 ;
        RECT 75.600 211.310 75.890 211.355 ;
        RECT 77.170 211.310 77.460 211.355 ;
        RECT 73.500 211.170 77.460 211.310 ;
        RECT 73.500 211.125 73.790 211.170 ;
        RECT 75.600 211.125 75.890 211.170 ;
        RECT 77.170 211.125 77.460 211.170 ;
        RECT 80.860 211.310 81.150 211.355 ;
        RECT 82.960 211.310 83.250 211.355 ;
        RECT 84.530 211.310 84.820 211.355 ;
        RECT 80.860 211.170 84.820 211.310 ;
        RECT 80.860 211.125 81.150 211.170 ;
        RECT 82.960 211.125 83.250 211.170 ;
        RECT 84.530 211.125 84.820 211.170 ;
        RECT 93.240 211.310 93.560 211.370 ;
        RECT 95.630 211.310 95.770 211.450 ;
        RECT 93.240 211.170 95.770 211.310 ;
        RECT 98.390 211.310 98.530 211.465 ;
        RECT 102.900 211.450 103.220 211.510 ;
        RECT 103.385 211.650 103.675 211.695 ;
        RECT 105.905 211.650 106.195 211.695 ;
        RECT 107.095 211.650 107.385 211.695 ;
        RECT 103.385 211.510 107.385 211.650 ;
        RECT 103.385 211.465 103.675 211.510 ;
        RECT 105.905 211.465 106.195 211.510 ;
        RECT 107.095 211.465 107.385 211.510 ;
        RECT 99.680 211.310 100.000 211.370 ;
        RECT 101.075 211.310 101.365 211.355 ;
        RECT 98.390 211.170 101.365 211.310 ;
        RECT 93.240 211.110 93.560 211.170 ;
        RECT 99.680 211.110 100.000 211.170 ;
        RECT 101.075 211.125 101.365 211.170 ;
        RECT 103.820 211.310 104.110 211.355 ;
        RECT 105.390 211.310 105.680 211.355 ;
        RECT 107.490 211.310 107.780 211.355 ;
        RECT 103.820 211.170 107.780 211.310 ;
        RECT 103.820 211.125 104.110 211.170 ;
        RECT 105.390 211.125 105.680 211.170 ;
        RECT 107.490 211.125 107.780 211.170 ;
        RECT 55.060 210.970 55.380 211.030 ;
        RECT 53.770 210.830 55.380 210.970 ;
        RECT 55.060 210.770 55.380 210.830 ;
        RECT 61.040 210.770 61.360 211.030 ;
        RECT 87.275 210.970 87.565 211.015 ;
        RECT 89.100 210.970 89.420 211.030 ;
        RECT 87.275 210.830 89.420 210.970 ;
        RECT 87.275 210.785 87.565 210.830 ;
        RECT 89.100 210.770 89.420 210.830 ;
        RECT 90.480 210.970 90.800 211.030 ;
        RECT 95.095 210.970 95.385 211.015 ;
        RECT 96.920 210.970 97.240 211.030 ;
        RECT 90.480 210.830 97.240 210.970 ;
        RECT 90.480 210.770 90.800 210.830 ;
        RECT 95.095 210.785 95.385 210.830 ;
        RECT 96.920 210.770 97.240 210.830 ;
        RECT 97.395 210.970 97.685 211.015 ;
        RECT 98.300 210.970 98.620 211.030 ;
        RECT 97.395 210.830 98.620 210.970 ;
        RECT 97.395 210.785 97.685 210.830 ;
        RECT 98.300 210.770 98.620 210.830 ;
        RECT 17.270 210.150 146.990 210.630 ;
        RECT 53.680 209.950 54.000 210.010 ;
        RECT 55.535 209.950 55.825 209.995 ;
        RECT 53.680 209.810 55.825 209.950 ;
        RECT 53.680 209.750 54.000 209.810 ;
        RECT 55.535 209.765 55.825 209.810 ;
        RECT 60.135 209.950 60.425 209.995 ;
        RECT 60.580 209.950 60.900 210.010 ;
        RECT 60.135 209.810 60.900 209.950 ;
        RECT 60.135 209.765 60.425 209.810 ;
        RECT 60.580 209.750 60.900 209.810 ;
        RECT 61.055 209.765 61.345 209.995 ;
        RECT 64.735 209.950 65.025 209.995 ;
        RECT 68.860 209.950 69.180 210.010 ;
        RECT 64.735 209.810 69.180 209.950 ;
        RECT 64.735 209.765 65.025 209.810 ;
        RECT 46.360 209.610 46.650 209.655 ;
        RECT 48.460 209.610 48.750 209.655 ;
        RECT 50.030 209.610 50.320 209.655 ;
        RECT 46.360 209.470 50.320 209.610 ;
        RECT 46.360 209.425 46.650 209.470 ;
        RECT 48.460 209.425 48.750 209.470 ;
        RECT 50.030 209.425 50.320 209.470 ;
        RECT 59.660 209.610 59.980 209.670 ;
        RECT 61.130 209.610 61.270 209.765 ;
        RECT 68.860 209.750 69.180 209.810 ;
        RECT 69.320 209.950 69.640 210.010 ;
        RECT 73.015 209.950 73.305 209.995 ;
        RECT 69.320 209.810 73.305 209.950 ;
        RECT 69.320 209.750 69.640 209.810 ;
        RECT 73.015 209.765 73.305 209.810 ;
        RECT 81.740 209.950 82.060 210.010 ;
        RECT 82.675 209.950 82.965 209.995 ;
        RECT 81.740 209.810 82.965 209.950 ;
        RECT 81.740 209.750 82.060 209.810 ;
        RECT 82.675 209.765 82.965 209.810 ;
        RECT 86.340 209.750 86.660 210.010 ;
        RECT 90.940 209.750 91.260 210.010 ;
        RECT 100.600 209.750 100.920 210.010 ;
        RECT 59.660 209.470 61.270 209.610 ;
        RECT 66.140 209.610 66.430 209.655 ;
        RECT 68.240 209.610 68.530 209.655 ;
        RECT 69.810 209.610 70.100 209.655 ;
        RECT 66.140 209.470 70.100 209.610 ;
        RECT 59.660 209.410 59.980 209.470 ;
        RECT 66.140 209.425 66.430 209.470 ;
        RECT 68.240 209.425 68.530 209.470 ;
        RECT 69.810 209.425 70.100 209.470 ;
        RECT 70.700 209.610 71.020 209.670 ;
        RECT 74.855 209.610 75.145 209.655 ;
        RECT 70.700 209.470 75.145 209.610 ;
        RECT 70.700 209.410 71.020 209.470 ;
        RECT 74.855 209.425 75.145 209.470 ;
        RECT 90.035 209.425 90.325 209.655 ;
        RECT 92.320 209.610 92.640 209.670 ;
        RECT 92.320 209.470 97.610 209.610 ;
        RECT 43.560 209.270 43.880 209.330 ;
        RECT 45.400 209.270 45.720 209.330 ;
        RECT 45.875 209.270 46.165 209.315 ;
        RECT 43.560 209.130 46.165 209.270 ;
        RECT 43.560 209.070 43.880 209.130 ;
        RECT 45.400 209.070 45.720 209.130 ;
        RECT 45.875 209.085 46.165 209.130 ;
        RECT 46.755 209.270 47.045 209.315 ;
        RECT 47.945 209.270 48.235 209.315 ;
        RECT 50.465 209.270 50.755 209.315 ;
        RECT 46.755 209.130 50.755 209.270 ;
        RECT 46.755 209.085 47.045 209.130 ;
        RECT 47.945 209.085 48.235 209.130 ;
        RECT 50.465 209.085 50.755 209.130 ;
        RECT 59.215 209.270 59.505 209.315 ;
        RECT 60.120 209.270 60.440 209.330 ;
        RECT 62.880 209.270 63.200 209.330 ;
        RECT 59.215 209.130 63.200 209.270 ;
        RECT 59.215 209.085 59.505 209.130 ;
        RECT 60.120 209.070 60.440 209.130 ;
        RECT 62.880 209.070 63.200 209.130 ;
        RECT 65.640 209.070 65.960 209.330 ;
        RECT 66.535 209.270 66.825 209.315 ;
        RECT 67.725 209.270 68.015 209.315 ;
        RECT 70.245 209.270 70.535 209.315 ;
        RECT 66.535 209.130 70.535 209.270 ;
        RECT 66.535 209.085 66.825 209.130 ;
        RECT 67.725 209.085 68.015 209.130 ;
        RECT 70.245 209.085 70.535 209.130 ;
        RECT 83.595 209.270 83.885 209.315 ;
        RECT 90.110 209.270 90.250 209.425 ;
        RECT 92.320 209.410 92.640 209.470 ;
        RECT 83.595 209.130 93.470 209.270 ;
        RECT 83.595 209.085 83.885 209.130 ;
        RECT 53.220 208.930 53.540 208.990 ;
        RECT 54.140 208.930 54.460 208.990 ;
        RECT 53.220 208.790 54.460 208.930 ;
        RECT 53.220 208.730 53.540 208.790 ;
        RECT 54.140 208.730 54.460 208.790 ;
        RECT 55.535 208.930 55.825 208.975 ;
        RECT 61.040 208.930 61.360 208.990 ;
        RECT 55.535 208.790 61.360 208.930 ;
        RECT 55.535 208.745 55.825 208.790 ;
        RECT 61.040 208.730 61.360 208.790 ;
        RECT 61.500 208.930 61.820 208.990 ;
        RECT 63.355 208.930 63.645 208.975 ;
        RECT 64.260 208.930 64.580 208.990 ;
        RECT 61.500 208.790 64.580 208.930 ;
        RECT 61.500 208.730 61.820 208.790 ;
        RECT 63.355 208.745 63.645 208.790 ;
        RECT 64.260 208.730 64.580 208.790 ;
        RECT 71.620 208.930 71.940 208.990 ;
        RECT 73.015 208.930 73.305 208.975 ;
        RECT 71.620 208.790 73.305 208.930 ;
        RECT 71.620 208.730 71.940 208.790 ;
        RECT 73.015 208.745 73.305 208.790 ;
        RECT 73.935 208.930 74.225 208.975 ;
        RECT 82.660 208.930 82.980 208.990 ;
        RECT 73.935 208.790 82.980 208.930 ;
        RECT 73.935 208.745 74.225 208.790 ;
        RECT 82.660 208.730 82.980 208.790 ;
        RECT 84.055 208.930 84.345 208.975 ;
        RECT 86.340 208.930 86.660 208.990 ;
        RECT 84.055 208.790 86.660 208.930 ;
        RECT 84.055 208.745 84.345 208.790 ;
        RECT 86.340 208.730 86.660 208.790 ;
        RECT 89.100 208.730 89.420 208.990 ;
        RECT 90.480 208.930 90.800 208.990 ;
        RECT 90.955 208.930 91.245 208.975 ;
        RECT 90.480 208.790 91.245 208.930 ;
        RECT 90.480 208.730 90.800 208.790 ;
        RECT 90.955 208.745 91.245 208.790 ;
        RECT 92.780 208.730 93.100 208.990 ;
        RECT 93.330 208.975 93.470 209.130 ;
        RECT 97.470 208.975 97.610 209.470 ;
        RECT 98.760 209.410 99.080 209.670 ;
        RECT 99.235 209.270 99.525 209.315 ;
        RECT 107.960 209.270 108.280 209.330 ;
        RECT 99.235 209.130 108.280 209.270 ;
        RECT 99.235 209.085 99.525 209.130 ;
        RECT 107.960 209.070 108.280 209.130 ;
        RECT 93.255 208.745 93.545 208.975 ;
        RECT 97.395 208.745 97.685 208.975 ;
        RECT 45.860 208.590 46.180 208.650 ;
        RECT 47.100 208.590 47.390 208.635 ;
        RECT 54.600 208.590 54.920 208.650 ;
        RECT 56.440 208.590 56.760 208.650 ;
        RECT 45.860 208.450 47.390 208.590 ;
        RECT 45.860 208.390 46.180 208.450 ;
        RECT 47.100 208.405 47.390 208.450 ;
        RECT 52.850 208.450 56.760 208.590 ;
        RECT 52.850 208.295 52.990 208.450 ;
        RECT 54.600 208.390 54.920 208.450 ;
        RECT 56.440 208.390 56.760 208.450 ;
        RECT 56.900 208.590 57.220 208.650 ;
        RECT 57.375 208.590 57.665 208.635 ;
        RECT 56.900 208.450 57.665 208.590 ;
        RECT 56.900 208.390 57.220 208.450 ;
        RECT 57.375 208.405 57.665 208.450 ;
        RECT 57.835 208.590 58.125 208.635 ;
        RECT 59.200 208.590 59.520 208.650 ;
        RECT 57.835 208.450 59.520 208.590 ;
        RECT 57.835 208.405 58.125 208.450 ;
        RECT 59.200 208.390 59.520 208.450 ;
        RECT 59.660 208.590 59.980 208.650 ;
        RECT 67.020 208.635 67.340 208.650 ;
        RECT 61.975 208.590 62.265 208.635 ;
        RECT 59.660 208.450 62.265 208.590 ;
        RECT 59.660 208.390 59.980 208.450 ;
        RECT 61.975 208.405 62.265 208.450 ;
        RECT 66.990 208.405 67.340 208.635 ;
        RECT 89.190 208.590 89.330 208.730 ;
        RECT 94.175 208.590 94.465 208.635 ;
        RECT 89.190 208.450 94.465 208.590 ;
        RECT 97.470 208.590 97.610 208.745 ;
        RECT 98.300 208.730 98.620 208.990 ;
        RECT 99.680 208.730 100.000 208.990 ;
        RECT 103.360 208.590 103.680 208.650 ;
        RECT 97.470 208.450 103.680 208.590 ;
        RECT 94.175 208.405 94.465 208.450 ;
        RECT 67.020 208.390 67.340 208.405 ;
        RECT 103.360 208.390 103.680 208.450 ;
        RECT 52.775 208.065 53.065 208.295 ;
        RECT 58.280 208.250 58.600 208.310 ;
        RECT 60.925 208.250 61.215 208.295 ;
        RECT 58.280 208.110 61.215 208.250 ;
        RECT 58.280 208.050 58.600 208.110 ;
        RECT 60.925 208.065 61.215 208.110 ;
        RECT 66.100 208.250 66.420 208.310 ;
        RECT 68.400 208.250 68.720 208.310 ;
        RECT 72.555 208.250 72.845 208.295 ;
        RECT 66.100 208.110 72.845 208.250 ;
        RECT 66.100 208.050 66.420 208.110 ;
        RECT 68.400 208.050 68.720 208.110 ;
        RECT 72.555 208.065 72.845 208.110 ;
        RECT 85.880 208.050 86.200 208.310 ;
        RECT 95.095 208.250 95.385 208.295 ;
        RECT 95.540 208.250 95.860 208.310 ;
        RECT 95.095 208.110 95.860 208.250 ;
        RECT 95.095 208.065 95.385 208.110 ;
        RECT 95.540 208.050 95.860 208.110 ;
        RECT 17.270 207.430 146.990 207.910 ;
        RECT 50.460 207.230 50.780 207.290 ;
        RECT 50.935 207.230 51.225 207.275 ;
        RECT 50.460 207.090 51.225 207.230 ;
        RECT 50.460 207.030 50.780 207.090 ;
        RECT 50.935 207.045 51.225 207.090 ;
        RECT 62.880 207.230 63.200 207.290 ;
        RECT 67.365 207.230 67.655 207.275 ;
        RECT 62.880 207.090 67.655 207.230 ;
        RECT 62.880 207.030 63.200 207.090 ;
        RECT 67.365 207.045 67.655 207.090 ;
        RECT 64.810 206.750 65.870 206.890 ;
        RECT 50.475 206.550 50.765 206.595 ;
        RECT 50.920 206.550 51.240 206.610 ;
        RECT 50.475 206.410 51.240 206.550 ;
        RECT 50.475 206.365 50.765 206.410 ;
        RECT 50.920 206.350 51.240 206.410 ;
        RECT 51.395 206.550 51.685 206.595 ;
        RECT 52.300 206.550 52.620 206.610 ;
        RECT 51.395 206.410 52.620 206.550 ;
        RECT 51.395 206.365 51.685 206.410 ;
        RECT 52.300 206.350 52.620 206.410 ;
        RECT 55.995 206.550 56.285 206.595 ;
        RECT 56.440 206.550 56.760 206.610 ;
        RECT 59.660 206.550 59.980 206.610 ;
        RECT 64.810 206.550 64.950 206.750 ;
        RECT 55.995 206.410 59.980 206.550 ;
        RECT 55.995 206.365 56.285 206.410 ;
        RECT 56.440 206.350 56.760 206.410 ;
        RECT 59.660 206.350 59.980 206.410 ;
        RECT 63.890 206.410 64.950 206.550 ;
        RECT 52.390 206.210 52.530 206.350 ;
        RECT 63.890 206.255 64.030 206.410 ;
        RECT 65.180 206.350 65.500 206.610 ;
        RECT 65.730 206.550 65.870 206.750 ;
        RECT 68.400 206.690 68.720 206.950 ;
        RECT 89.560 206.890 89.880 206.950 ;
        RECT 86.430 206.750 89.880 206.890 ;
        RECT 65.730 206.410 69.550 206.550 ;
        RECT 63.815 206.210 64.105 206.255 ;
        RECT 68.860 206.210 69.180 206.270 ;
        RECT 52.390 206.070 64.105 206.210 ;
        RECT 63.815 206.025 64.105 206.070 ;
        RECT 64.810 206.070 69.180 206.210 ;
        RECT 50.460 205.870 50.780 205.930 ;
        RECT 59.200 205.870 59.520 205.930 ;
        RECT 64.810 205.915 64.950 206.070 ;
        RECT 68.860 206.010 69.180 206.070 ;
        RECT 50.460 205.730 59.520 205.870 ;
        RECT 50.460 205.670 50.780 205.730 ;
        RECT 59.200 205.670 59.520 205.730 ;
        RECT 64.735 205.685 65.025 205.915 ;
        RECT 65.195 205.870 65.485 205.915 ;
        RECT 67.020 205.870 67.340 205.930 ;
        RECT 65.195 205.730 67.340 205.870 ;
        RECT 69.410 205.870 69.550 206.410 ;
        RECT 70.700 206.350 71.020 206.610 ;
        RECT 86.430 206.595 86.570 206.750 ;
        RECT 89.560 206.690 89.880 206.750 ;
        RECT 86.355 206.365 86.645 206.595 ;
        RECT 87.735 206.550 88.025 206.595 ;
        RECT 89.100 206.550 89.420 206.610 ;
        RECT 87.735 206.410 89.420 206.550 ;
        RECT 87.735 206.365 88.025 206.410 ;
        RECT 89.100 206.350 89.420 206.410 ;
        RECT 94.160 206.550 94.480 206.610 ;
        RECT 95.095 206.550 95.385 206.595 ;
        RECT 94.160 206.410 95.385 206.550 ;
        RECT 94.160 206.350 94.480 206.410 ;
        RECT 95.095 206.365 95.385 206.410 ;
        RECT 96.000 206.350 96.320 206.610 ;
        RECT 107.960 206.550 108.280 206.610 ;
        RECT 113.955 206.550 114.245 206.595 ;
        RECT 107.960 206.410 114.245 206.550 ;
        RECT 107.960 206.350 108.280 206.410 ;
        RECT 113.955 206.365 114.245 206.410 ;
        RECT 108.420 206.210 108.740 206.270 ;
        RECT 110.735 206.210 111.025 206.255 ;
        RECT 108.420 206.070 111.025 206.210 ;
        RECT 108.420 206.010 108.740 206.070 ;
        RECT 110.735 206.025 111.025 206.070 ;
        RECT 69.795 205.870 70.085 205.915 ;
        RECT 72.540 205.870 72.860 205.930 ;
        RECT 69.410 205.730 72.860 205.870 ;
        RECT 65.195 205.685 65.485 205.730 ;
        RECT 51.380 205.530 51.700 205.590 ;
        RECT 55.535 205.530 55.825 205.575 ;
        RECT 51.380 205.390 55.825 205.530 ;
        RECT 64.810 205.530 64.950 205.685 ;
        RECT 67.020 205.670 67.340 205.730 ;
        RECT 69.795 205.685 70.085 205.730 ;
        RECT 72.540 205.670 72.860 205.730 ;
        RECT 66.575 205.530 66.865 205.575 ;
        RECT 64.810 205.390 66.865 205.530 ;
        RECT 51.380 205.330 51.700 205.390 ;
        RECT 55.535 205.345 55.825 205.390 ;
        RECT 66.575 205.345 66.865 205.390 ;
        RECT 67.480 205.330 67.800 205.590 ;
        RECT 80.820 205.530 81.140 205.590 ;
        RECT 84.960 205.530 85.280 205.590 ;
        RECT 85.435 205.530 85.725 205.575 ;
        RECT 80.820 205.390 85.725 205.530 ;
        RECT 80.820 205.330 81.140 205.390 ;
        RECT 84.960 205.330 85.280 205.390 ;
        RECT 85.435 205.345 85.725 205.390 ;
        RECT 87.275 205.530 87.565 205.575 ;
        RECT 91.400 205.530 91.720 205.590 ;
        RECT 87.275 205.390 91.720 205.530 ;
        RECT 87.275 205.345 87.565 205.390 ;
        RECT 91.400 205.330 91.720 205.390 ;
        RECT 94.620 205.530 94.940 205.590 ;
        RECT 95.095 205.530 95.385 205.575 ;
        RECT 94.620 205.390 95.385 205.530 ;
        RECT 94.620 205.330 94.940 205.390 ;
        RECT 95.095 205.345 95.385 205.390 ;
        RECT 17.270 204.710 146.990 205.190 ;
        RECT 61.500 204.510 61.820 204.570 ;
        RECT 67.480 204.510 67.800 204.570 ;
        RECT 61.500 204.370 67.800 204.510 ;
        RECT 61.500 204.310 61.820 204.370 ;
        RECT 67.480 204.310 67.800 204.370 ;
        RECT 81.280 204.510 81.600 204.570 ;
        RECT 85.880 204.510 86.200 204.570 ;
        RECT 93.255 204.510 93.545 204.555 ;
        RECT 81.280 204.370 93.545 204.510 ;
        RECT 81.280 204.310 81.600 204.370 ;
        RECT 85.880 204.310 86.200 204.370 ;
        RECT 93.255 204.325 93.545 204.370 ;
        RECT 95.540 204.310 95.860 204.570 ;
        RECT 96.000 204.510 96.320 204.570 ;
        RECT 97.840 204.510 98.160 204.570 ;
        RECT 103.375 204.510 103.665 204.555 ;
        RECT 96.000 204.370 103.665 204.510 ;
        RECT 96.000 204.310 96.320 204.370 ;
        RECT 97.840 204.310 98.160 204.370 ;
        RECT 103.375 204.325 103.665 204.370 ;
        RECT 42.640 204.170 42.960 204.230 ;
        RECT 59.215 204.170 59.505 204.215 ;
        RECT 60.580 204.170 60.900 204.230 ;
        RECT 42.640 204.030 58.510 204.170 ;
        RECT 42.640 203.970 42.960 204.030 ;
        RECT 52.760 203.830 53.080 203.890 ;
        RECT 56.915 203.830 57.205 203.875 ;
        RECT 52.760 203.690 57.205 203.830 ;
        RECT 52.760 203.630 53.080 203.690 ;
        RECT 56.915 203.645 57.205 203.690 ;
        RECT 21.480 203.490 21.800 203.550 ;
        RECT 26.080 203.490 26.400 203.550 ;
        RECT 21.480 203.350 26.400 203.490 ;
        RECT 21.480 203.290 21.800 203.350 ;
        RECT 26.080 203.290 26.400 203.350 ;
        RECT 26.555 203.490 26.845 203.535 ;
        RECT 32.060 203.490 32.380 203.550 ;
        RECT 26.555 203.350 32.380 203.490 ;
        RECT 26.555 203.305 26.845 203.350 ;
        RECT 32.060 203.290 32.380 203.350 ;
        RECT 54.140 203.490 54.460 203.550 ;
        RECT 56.455 203.490 56.745 203.535 ;
        RECT 54.140 203.350 56.745 203.490 ;
        RECT 54.140 203.290 54.460 203.350 ;
        RECT 56.455 203.305 56.745 203.350 ;
        RECT 27.475 203.150 27.765 203.195 ;
        RECT 28.840 203.150 29.160 203.210 ;
        RECT 27.475 203.010 29.160 203.150 ;
        RECT 27.475 202.965 27.765 203.010 ;
        RECT 28.840 202.950 29.160 203.010 ;
        RECT 39.420 202.950 39.740 203.210 ;
        RECT 53.680 202.950 54.000 203.210 ;
        RECT 54.615 203.150 54.905 203.195 ;
        RECT 55.980 203.150 56.300 203.210 ;
        RECT 54.615 203.010 56.300 203.150 ;
        RECT 54.615 202.965 54.905 203.010 ;
        RECT 55.980 202.950 56.300 203.010 ;
        RECT 27.000 202.610 27.320 202.870 ;
        RECT 39.880 202.610 40.200 202.870 ;
        RECT 55.060 202.810 55.380 202.870 ;
        RECT 55.535 202.810 55.825 202.855 ;
        RECT 55.060 202.670 55.825 202.810 ;
        RECT 56.530 202.810 56.670 203.305 ;
        RECT 56.990 203.150 57.130 203.645 ;
        RECT 57.835 203.490 58.125 203.535 ;
        RECT 58.370 203.490 58.510 204.030 ;
        RECT 59.215 204.030 60.900 204.170 ;
        RECT 59.215 203.985 59.505 204.030 ;
        RECT 60.580 203.970 60.900 204.030 ;
        RECT 80.360 204.170 80.680 204.230 ;
        RECT 82.700 204.170 82.990 204.215 ;
        RECT 84.800 204.170 85.090 204.215 ;
        RECT 86.370 204.170 86.660 204.215 ;
        RECT 80.360 204.030 82.430 204.170 ;
        RECT 80.360 203.970 80.680 204.030 ;
        RECT 58.740 203.630 59.060 203.890 ;
        RECT 81.280 203.630 81.600 203.890 ;
        RECT 82.290 203.875 82.430 204.030 ;
        RECT 82.700 204.030 86.660 204.170 ;
        RECT 82.700 203.985 82.990 204.030 ;
        RECT 84.800 203.985 85.090 204.030 ;
        RECT 86.370 203.985 86.660 204.030 ;
        RECT 89.115 204.170 89.405 204.215 ;
        RECT 96.960 204.170 97.250 204.215 ;
        RECT 99.060 204.170 99.350 204.215 ;
        RECT 100.630 204.170 100.920 204.215 ;
        RECT 89.115 204.030 92.550 204.170 ;
        RECT 89.115 203.985 89.405 204.030 ;
        RECT 92.410 203.875 92.550 204.030 ;
        RECT 96.960 204.030 100.920 204.170 ;
        RECT 96.960 203.985 97.250 204.030 ;
        RECT 99.060 203.985 99.350 204.030 ;
        RECT 100.630 203.985 100.920 204.030 ;
        RECT 82.215 203.645 82.505 203.875 ;
        RECT 83.095 203.830 83.385 203.875 ;
        RECT 84.285 203.830 84.575 203.875 ;
        RECT 86.805 203.830 87.095 203.875 ;
        RECT 83.095 203.690 87.095 203.830 ;
        RECT 83.095 203.645 83.385 203.690 ;
        RECT 84.285 203.645 84.575 203.690 ;
        RECT 86.805 203.645 87.095 203.690 ;
        RECT 92.335 203.830 92.625 203.875 ;
        RECT 94.635 203.830 94.925 203.875 ;
        RECT 92.335 203.690 94.925 203.830 ;
        RECT 92.335 203.645 92.625 203.690 ;
        RECT 94.635 203.645 94.925 203.690 ;
        RECT 96.460 203.630 96.780 203.890 ;
        RECT 97.355 203.830 97.645 203.875 ;
        RECT 98.545 203.830 98.835 203.875 ;
        RECT 101.065 203.830 101.355 203.875 ;
        RECT 97.355 203.690 101.355 203.830 ;
        RECT 103.450 203.830 103.590 204.325 ;
        RECT 111.180 204.170 111.470 204.215 ;
        RECT 112.750 204.170 113.040 204.215 ;
        RECT 114.850 204.170 115.140 204.215 ;
        RECT 111.180 204.030 115.140 204.170 ;
        RECT 111.180 203.985 111.470 204.030 ;
        RECT 112.750 203.985 113.040 204.030 ;
        RECT 114.850 203.985 115.140 204.030 ;
        RECT 106.595 203.830 106.885 203.875 ;
        RECT 103.450 203.690 106.885 203.830 ;
        RECT 97.355 203.645 97.645 203.690 ;
        RECT 98.545 203.645 98.835 203.690 ;
        RECT 101.065 203.645 101.355 203.690 ;
        RECT 106.595 203.645 106.885 203.690 ;
        RECT 110.745 203.830 111.035 203.875 ;
        RECT 113.265 203.830 113.555 203.875 ;
        RECT 114.455 203.830 114.745 203.875 ;
        RECT 110.745 203.690 114.745 203.830 ;
        RECT 110.745 203.645 111.035 203.690 ;
        RECT 113.265 203.645 113.555 203.690 ;
        RECT 114.455 203.645 114.745 203.690 ;
        RECT 60.595 203.490 60.885 203.535 ;
        RECT 62.420 203.490 62.740 203.550 ;
        RECT 57.835 203.350 62.740 203.490 ;
        RECT 57.835 203.305 58.125 203.350 ;
        RECT 60.595 203.305 60.885 203.350 ;
        RECT 62.420 203.290 62.740 203.350 ;
        RECT 79.900 203.290 80.220 203.550 ;
        RECT 80.375 203.490 80.665 203.535 ;
        RECT 80.820 203.490 81.140 203.550 ;
        RECT 89.575 203.490 89.865 203.535 ;
        RECT 80.375 203.350 81.140 203.490 ;
        RECT 80.375 203.305 80.665 203.350 ;
        RECT 80.820 203.290 81.140 203.350 ;
        RECT 82.750 203.350 89.865 203.490 ;
        RECT 59.215 203.150 59.505 203.195 ;
        RECT 56.990 203.010 59.505 203.150 ;
        RECT 59.215 202.965 59.505 203.010 ;
        RECT 82.200 203.150 82.520 203.210 ;
        RECT 82.750 203.150 82.890 203.350 ;
        RECT 89.575 203.305 89.865 203.350 ;
        RECT 91.400 203.490 91.720 203.550 ;
        RECT 96.015 203.490 96.305 203.535 ;
        RECT 91.400 203.350 96.305 203.490 ;
        RECT 91.400 203.290 91.720 203.350 ;
        RECT 96.015 203.305 96.305 203.350 ;
        RECT 107.960 203.490 108.280 203.550 ;
        RECT 115.335 203.490 115.625 203.535 ;
        RECT 107.960 203.350 115.625 203.490 ;
        RECT 107.960 203.290 108.280 203.350 ;
        RECT 115.335 203.305 115.625 203.350 ;
        RECT 82.200 203.010 82.890 203.150 ;
        RECT 83.550 203.150 83.840 203.195 ;
        RECT 85.880 203.150 86.200 203.210 ;
        RECT 83.550 203.010 86.200 203.150 ;
        RECT 82.200 202.950 82.520 203.010 ;
        RECT 83.550 202.965 83.840 203.010 ;
        RECT 85.880 202.950 86.200 203.010 ;
        RECT 97.810 203.150 98.100 203.195 ;
        RECT 99.220 203.150 99.540 203.210 ;
        RECT 106.120 203.150 106.440 203.210 ;
        RECT 97.810 203.010 99.540 203.150 ;
        RECT 97.810 202.965 98.100 203.010 ;
        RECT 99.220 202.950 99.540 203.010 ;
        RECT 101.610 203.010 106.440 203.150 ;
        RECT 101.610 202.870 101.750 203.010 ;
        RECT 106.120 202.950 106.440 203.010 ;
        RECT 114.110 203.150 114.400 203.195 ;
        RECT 114.860 203.150 115.180 203.210 ;
        RECT 114.110 203.010 115.180 203.150 ;
        RECT 114.110 202.965 114.400 203.010 ;
        RECT 114.860 202.950 115.180 203.010 ;
        RECT 58.280 202.810 58.600 202.870 ;
        RECT 60.135 202.810 60.425 202.855 ;
        RECT 56.530 202.670 60.425 202.810 ;
        RECT 55.060 202.610 55.380 202.670 ;
        RECT 55.535 202.625 55.825 202.670 ;
        RECT 58.280 202.610 58.600 202.670 ;
        RECT 60.135 202.625 60.425 202.670 ;
        RECT 81.295 202.810 81.585 202.855 ;
        RECT 82.660 202.810 82.980 202.870 ;
        RECT 81.295 202.670 82.980 202.810 ;
        RECT 81.295 202.625 81.585 202.670 ;
        RECT 82.660 202.610 82.980 202.670 ;
        RECT 94.160 202.810 94.480 202.870 ;
        RECT 101.520 202.810 101.840 202.870 ;
        RECT 94.160 202.670 101.840 202.810 ;
        RECT 94.160 202.610 94.480 202.670 ;
        RECT 101.520 202.610 101.840 202.670 ;
        RECT 103.820 202.610 104.140 202.870 ;
        RECT 108.420 202.610 108.740 202.870 ;
        RECT 17.270 201.990 146.990 202.470 ;
        RECT 19.655 201.790 19.945 201.835 ;
        RECT 39.420 201.790 39.740 201.850 ;
        RECT 19.655 201.650 39.740 201.790 ;
        RECT 19.655 201.605 19.945 201.650 ;
        RECT 39.420 201.590 39.740 201.650 ;
        RECT 51.380 201.590 51.700 201.850 ;
        RECT 52.760 201.790 53.080 201.850 ;
        RECT 54.615 201.790 54.905 201.835 ;
        RECT 55.060 201.790 55.380 201.850 ;
        RECT 52.760 201.650 53.450 201.790 ;
        RECT 52.760 201.590 53.080 201.650 ;
        RECT 21.480 201.250 21.800 201.510 ;
        RECT 43.560 201.450 43.880 201.510 ;
        RECT 25.250 201.310 43.880 201.450 ;
        RECT 25.250 201.170 25.390 201.310 ;
        RECT 18.720 200.910 19.040 201.170 ;
        RECT 25.160 200.910 25.480 201.170 ;
        RECT 25.620 201.110 25.940 201.170 ;
        RECT 32.610 201.155 32.750 201.310 ;
        RECT 43.560 201.250 43.880 201.310 ;
        RECT 46.320 201.450 46.640 201.510 ;
        RECT 50.935 201.450 51.225 201.495 ;
        RECT 51.840 201.450 52.160 201.510 ;
        RECT 53.310 201.495 53.450 201.650 ;
        RECT 54.615 201.650 55.380 201.790 ;
        RECT 54.615 201.605 54.905 201.650 ;
        RECT 55.060 201.590 55.380 201.650 ;
        RECT 55.535 201.790 55.825 201.835 ;
        RECT 79.900 201.790 80.220 201.850 ;
        RECT 81.755 201.790 82.045 201.835 ;
        RECT 55.535 201.650 56.210 201.790 ;
        RECT 55.535 201.605 55.825 201.650 ;
        RECT 46.320 201.310 52.160 201.450 ;
        RECT 46.320 201.250 46.640 201.310 ;
        RECT 26.455 201.110 26.745 201.155 ;
        RECT 25.620 200.970 26.745 201.110 ;
        RECT 25.620 200.910 25.940 200.970 ;
        RECT 26.455 200.925 26.745 200.970 ;
        RECT 32.535 200.925 32.825 201.155 ;
        RECT 33.870 201.110 34.160 201.155 ;
        RECT 35.740 201.110 36.060 201.170 ;
        RECT 33.870 200.970 36.060 201.110 ;
        RECT 33.870 200.925 34.160 200.970 ;
        RECT 35.740 200.910 36.060 200.970 ;
        RECT 39.895 200.925 40.185 201.155 ;
        RECT 26.055 200.770 26.345 200.815 ;
        RECT 27.245 200.770 27.535 200.815 ;
        RECT 29.765 200.770 30.055 200.815 ;
        RECT 26.055 200.630 30.055 200.770 ;
        RECT 26.055 200.585 26.345 200.630 ;
        RECT 27.245 200.585 27.535 200.630 ;
        RECT 29.765 200.585 30.055 200.630 ;
        RECT 33.415 200.770 33.705 200.815 ;
        RECT 34.605 200.770 34.895 200.815 ;
        RECT 37.125 200.770 37.415 200.815 ;
        RECT 33.415 200.630 37.415 200.770 ;
        RECT 33.415 200.585 33.705 200.630 ;
        RECT 34.605 200.585 34.895 200.630 ;
        RECT 37.125 200.585 37.415 200.630 ;
        RECT 23.335 200.430 23.625 200.475 ;
        RECT 24.700 200.430 25.020 200.490 ;
        RECT 23.335 200.290 25.020 200.430 ;
        RECT 23.335 200.245 23.625 200.290 ;
        RECT 24.700 200.230 25.020 200.290 ;
        RECT 25.660 200.430 25.950 200.475 ;
        RECT 27.760 200.430 28.050 200.475 ;
        RECT 29.330 200.430 29.620 200.475 ;
        RECT 25.660 200.290 29.620 200.430 ;
        RECT 25.660 200.245 25.950 200.290 ;
        RECT 27.760 200.245 28.050 200.290 ;
        RECT 29.330 200.245 29.620 200.290 ;
        RECT 32.060 200.230 32.380 200.490 ;
        RECT 33.020 200.430 33.310 200.475 ;
        RECT 35.120 200.430 35.410 200.475 ;
        RECT 36.690 200.430 36.980 200.475 ;
        RECT 33.020 200.290 36.980 200.430 ;
        RECT 33.020 200.245 33.310 200.290 ;
        RECT 35.120 200.245 35.410 200.290 ;
        RECT 36.690 200.245 36.980 200.290 ;
        RECT 39.435 200.430 39.725 200.475 ;
        RECT 39.970 200.430 40.110 200.925 ;
        RECT 40.800 200.910 41.120 201.170 ;
        RECT 42.655 201.110 42.945 201.155 ;
        RECT 44.940 201.110 45.260 201.170 ;
        RECT 45.430 201.155 45.690 201.200 ;
        RECT 48.710 201.155 48.850 201.310 ;
        RECT 50.935 201.265 51.225 201.310 ;
        RECT 51.840 201.250 52.160 201.310 ;
        RECT 53.235 201.265 53.525 201.495 ;
        RECT 56.070 201.450 56.210 201.650 ;
        RECT 79.900 201.650 82.045 201.790 ;
        RECT 79.900 201.590 80.220 201.650 ;
        RECT 81.755 201.605 82.045 201.650 ;
        RECT 85.880 201.590 86.200 201.850 ;
        RECT 94.160 201.590 94.480 201.850 ;
        RECT 95.540 201.790 95.860 201.850 ;
        RECT 97.395 201.790 97.685 201.835 ;
        RECT 95.540 201.650 97.685 201.790 ;
        RECT 95.540 201.590 95.860 201.650 ;
        RECT 97.395 201.605 97.685 201.650 ;
        RECT 77.155 201.450 77.445 201.495 ;
        RECT 78.520 201.450 78.840 201.510 ;
        RECT 80.360 201.450 80.680 201.510 ;
        RECT 89.560 201.450 89.880 201.510 ;
        RECT 96.920 201.450 97.240 201.510 ;
        RECT 54.690 201.310 56.210 201.450 ;
        RECT 56.530 201.310 64.490 201.450 ;
        RECT 42.655 200.970 45.260 201.110 ;
        RECT 42.655 200.925 42.945 200.970 ;
        RECT 44.940 200.910 45.260 200.970 ;
        RECT 45.415 201.110 45.705 201.155 ;
        RECT 48.175 201.110 48.465 201.155 ;
        RECT 45.415 200.970 48.465 201.110 ;
        RECT 45.415 200.925 45.705 200.970 ;
        RECT 48.175 200.925 48.465 200.970 ;
        RECT 48.635 200.925 48.925 201.155 ;
        RECT 52.775 201.110 53.065 201.155 ;
        RECT 54.140 201.110 54.460 201.170 ;
        RECT 52.775 200.970 54.460 201.110 ;
        RECT 52.775 200.925 53.065 200.970 ;
        RECT 45.430 200.880 45.690 200.925 ;
        RECT 54.140 200.910 54.460 200.970 ;
        RECT 43.100 200.770 43.420 200.830 ;
        RECT 43.575 200.770 43.865 200.815 ;
        RECT 43.100 200.630 43.865 200.770 ;
        RECT 43.100 200.570 43.420 200.630 ;
        RECT 43.575 200.585 43.865 200.630 ;
        RECT 51.840 200.770 52.160 200.830 ;
        RECT 54.690 200.770 54.830 201.310 ;
        RECT 55.075 201.110 55.365 201.155 ;
        RECT 56.530 201.110 56.670 201.310 ;
        RECT 55.075 200.970 56.670 201.110 ;
        RECT 55.075 200.925 55.365 200.970 ;
        RECT 56.915 200.925 57.205 201.155 ;
        RECT 51.840 200.630 54.830 200.770 ;
        RECT 51.840 200.570 52.160 200.630 ;
        RECT 40.340 200.430 40.660 200.490 ;
        RECT 39.435 200.290 40.660 200.430 ;
        RECT 39.435 200.245 39.725 200.290 ;
        RECT 40.340 200.230 40.660 200.290 ;
        RECT 53.695 200.430 53.985 200.475 ;
        RECT 54.600 200.430 54.920 200.490 ;
        RECT 53.695 200.290 54.920 200.430 ;
        RECT 53.695 200.245 53.985 200.290 ;
        RECT 54.600 200.230 54.920 200.290 ;
        RECT 56.455 200.430 56.745 200.475 ;
        RECT 56.990 200.430 57.130 200.925 ;
        RECT 58.740 200.910 59.060 201.170 ;
        RECT 59.200 200.910 59.520 201.170 ;
        RECT 61.500 200.910 61.820 201.170 ;
        RECT 64.350 201.155 64.490 201.310 ;
        RECT 77.155 201.310 87.490 201.450 ;
        RECT 77.155 201.265 77.445 201.310 ;
        RECT 78.520 201.250 78.840 201.310 ;
        RECT 80.360 201.250 80.680 201.310 ;
        RECT 62.435 201.110 62.725 201.155 ;
        RECT 64.275 201.110 64.565 201.155 ;
        RECT 66.560 201.110 66.880 201.170 ;
        RECT 62.435 200.970 64.030 201.110 ;
        RECT 62.435 200.925 62.725 200.970 ;
        RECT 57.360 200.770 57.680 200.830 ;
        RECT 59.290 200.770 59.430 200.910 ;
        RECT 57.360 200.630 59.430 200.770 ;
        RECT 57.360 200.570 57.680 200.630 ;
        RECT 62.880 200.570 63.200 200.830 ;
        RECT 63.890 200.770 64.030 200.970 ;
        RECT 64.275 200.970 66.880 201.110 ;
        RECT 64.275 200.925 64.565 200.970 ;
        RECT 66.560 200.910 66.880 200.970 ;
        RECT 68.860 201.110 69.180 201.170 ;
        RECT 74.395 201.110 74.685 201.155 ;
        RECT 68.860 200.970 74.685 201.110 ;
        RECT 68.860 200.910 69.180 200.970 ;
        RECT 74.395 200.925 74.685 200.970 ;
        RECT 80.820 200.910 81.140 201.170 ;
        RECT 82.200 200.910 82.520 201.170 ;
        RECT 82.660 200.910 82.980 201.170 ;
        RECT 87.350 201.155 87.490 201.310 ;
        RECT 89.560 201.310 97.240 201.450 ;
        RECT 97.470 201.450 97.610 201.605 ;
        RECT 99.220 201.590 99.540 201.850 ;
        RECT 102.900 201.590 103.220 201.850 ;
        RECT 107.500 201.790 107.820 201.850 ;
        RECT 112.575 201.790 112.865 201.835 ;
        RECT 107.500 201.650 112.865 201.790 ;
        RECT 107.500 201.590 107.820 201.650 ;
        RECT 112.575 201.605 112.865 201.650 ;
        RECT 114.860 201.590 115.180 201.850 ;
        RECT 103.820 201.450 104.140 201.510 ;
        RECT 97.470 201.310 101.290 201.450 ;
        RECT 89.560 201.250 89.880 201.310 ;
        RECT 96.920 201.250 97.240 201.310 ;
        RECT 87.275 200.925 87.565 201.155 ;
        RECT 88.610 201.110 88.900 201.155 ;
        RECT 92.320 201.110 92.640 201.170 ;
        RECT 88.610 200.970 92.640 201.110 ;
        RECT 88.610 200.925 88.900 200.970 ;
        RECT 92.320 200.910 92.640 200.970 ;
        RECT 94.620 201.110 94.940 201.170 ;
        RECT 99.220 201.110 99.540 201.170 ;
        RECT 101.150 201.155 101.290 201.310 ;
        RECT 101.610 201.310 104.140 201.450 ;
        RECT 101.610 201.155 101.750 201.310 ;
        RECT 103.820 201.250 104.140 201.310 ;
        RECT 100.155 201.110 100.445 201.155 ;
        RECT 94.620 200.970 98.990 201.110 ;
        RECT 94.620 200.910 94.940 200.970 ;
        RECT 66.100 200.770 66.420 200.830 ;
        RECT 63.890 200.630 66.420 200.770 ;
        RECT 66.100 200.570 66.420 200.630 ;
        RECT 67.020 200.770 67.340 200.830 ;
        RECT 72.555 200.770 72.845 200.815 ;
        RECT 75.300 200.770 75.620 200.830 ;
        RECT 67.020 200.630 75.620 200.770 ;
        RECT 67.020 200.570 67.340 200.630 ;
        RECT 72.555 200.585 72.845 200.630 ;
        RECT 75.300 200.570 75.620 200.630 ;
        RECT 88.155 200.770 88.445 200.815 ;
        RECT 89.345 200.770 89.635 200.815 ;
        RECT 91.865 200.770 92.155 200.815 ;
        RECT 88.155 200.630 92.155 200.770 ;
        RECT 88.155 200.585 88.445 200.630 ;
        RECT 89.345 200.585 89.635 200.630 ;
        RECT 91.865 200.585 92.155 200.630 ;
        RECT 98.315 200.585 98.605 200.815 ;
        RECT 65.180 200.430 65.500 200.490 ;
        RECT 56.455 200.290 65.500 200.430 ;
        RECT 56.455 200.245 56.745 200.290 ;
        RECT 65.180 200.230 65.500 200.290 ;
        RECT 87.760 200.430 88.050 200.475 ;
        RECT 89.860 200.430 90.150 200.475 ;
        RECT 91.430 200.430 91.720 200.475 ;
        RECT 87.760 200.290 91.720 200.430 ;
        RECT 87.760 200.245 88.050 200.290 ;
        RECT 89.860 200.245 90.150 200.290 ;
        RECT 91.430 200.245 91.720 200.290 ;
        RECT 98.390 200.150 98.530 200.585 ;
        RECT 98.850 200.430 98.990 200.970 ;
        RECT 99.220 200.970 100.445 201.110 ;
        RECT 99.220 200.910 99.540 200.970 ;
        RECT 100.155 200.925 100.445 200.970 ;
        RECT 101.075 200.925 101.365 201.155 ;
        RECT 101.535 200.925 101.825 201.155 ;
        RECT 102.440 200.910 102.760 201.170 ;
        RECT 104.295 201.110 104.585 201.155 ;
        RECT 102.990 200.970 104.585 201.110 ;
        RECT 99.680 200.770 100.000 200.830 ;
        RECT 102.990 200.770 103.130 200.970 ;
        RECT 104.295 200.925 104.585 200.970 ;
        RECT 106.120 200.910 106.440 201.170 ;
        RECT 113.035 201.110 113.325 201.155 ;
        RECT 120.840 201.110 121.160 201.170 ;
        RECT 113.035 200.970 121.160 201.110 ;
        RECT 113.035 200.925 113.325 200.970 ;
        RECT 120.840 200.910 121.160 200.970 ;
        RECT 99.680 200.630 103.130 200.770 ;
        RECT 99.680 200.570 100.000 200.630 ;
        RECT 103.820 200.570 104.140 200.830 ;
        RECT 104.740 200.570 105.060 200.830 ;
        RECT 105.200 200.570 105.520 200.830 ;
        RECT 107.040 200.770 107.360 200.830 ;
        RECT 111.655 200.770 111.945 200.815 ;
        RECT 107.040 200.630 111.945 200.770 ;
        RECT 107.040 200.570 107.360 200.630 ;
        RECT 111.655 200.585 111.945 200.630 ;
        RECT 100.615 200.430 100.905 200.475 ;
        RECT 98.850 200.290 100.905 200.430 ;
        RECT 100.615 200.245 100.905 200.290 ;
        RECT 23.780 199.890 24.100 200.150 ;
        RECT 39.880 199.890 40.200 200.150 ;
        RECT 41.735 200.090 42.025 200.135 ;
        RECT 42.640 200.090 42.960 200.150 ;
        RECT 41.735 199.950 42.960 200.090 ;
        RECT 41.735 199.905 42.025 199.950 ;
        RECT 42.640 199.890 42.960 199.950 ;
        RECT 48.175 200.090 48.465 200.135 ;
        RECT 49.095 200.090 49.385 200.135 ;
        RECT 48.175 199.950 49.385 200.090 ;
        RECT 48.175 199.905 48.465 199.950 ;
        RECT 49.095 199.905 49.385 199.950 ;
        RECT 52.300 199.890 52.620 200.150 ;
        RECT 53.220 200.090 53.540 200.150 ;
        RECT 56.900 200.090 57.220 200.150 ;
        RECT 53.220 199.950 57.220 200.090 ;
        RECT 53.220 199.890 53.540 199.950 ;
        RECT 56.900 199.890 57.220 199.950 ;
        RECT 57.360 199.890 57.680 200.150 ;
        RECT 60.120 199.890 60.440 200.150 ;
        RECT 60.595 200.090 60.885 200.135 ;
        RECT 61.040 200.090 61.360 200.150 ;
        RECT 60.595 199.950 61.360 200.090 ;
        RECT 60.595 199.905 60.885 199.950 ;
        RECT 61.040 199.890 61.360 199.950 ;
        RECT 63.800 199.890 64.120 200.150 ;
        RECT 69.780 199.890 70.100 200.150 ;
        RECT 73.460 199.890 73.780 200.150 ;
        RECT 94.620 200.090 94.940 200.150 ;
        RECT 95.095 200.090 95.385 200.135 ;
        RECT 94.620 199.950 95.385 200.090 ;
        RECT 94.620 199.890 94.940 199.950 ;
        RECT 95.095 199.905 95.385 199.950 ;
        RECT 98.300 200.090 98.620 200.150 ;
        RECT 106.580 200.090 106.900 200.150 ;
        RECT 98.300 199.950 106.900 200.090 ;
        RECT 98.300 199.890 98.620 199.950 ;
        RECT 106.580 199.890 106.900 199.950 ;
        RECT 17.270 199.270 146.990 199.750 ;
        RECT 35.740 198.870 36.060 199.130 ;
        RECT 36.675 198.885 36.965 199.115 ;
        RECT 48.635 199.070 48.925 199.115 ;
        RECT 57.360 199.070 57.680 199.130 ;
        RECT 63.355 199.070 63.645 199.115 ;
        RECT 48.635 198.930 63.645 199.070 ;
        RECT 48.635 198.885 48.925 198.930 ;
        RECT 21.980 198.730 22.270 198.775 ;
        RECT 24.080 198.730 24.370 198.775 ;
        RECT 25.650 198.730 25.940 198.775 ;
        RECT 21.980 198.590 25.940 198.730 ;
        RECT 21.980 198.545 22.270 198.590 ;
        RECT 24.080 198.545 24.370 198.590 ;
        RECT 25.650 198.545 25.940 198.590 ;
        RECT 29.315 198.730 29.605 198.775 ;
        RECT 36.750 198.730 36.890 198.885 ;
        RECT 57.360 198.870 57.680 198.930 ;
        RECT 63.355 198.885 63.645 198.930 ;
        RECT 66.100 198.870 66.420 199.130 ;
        RECT 66.560 198.870 66.880 199.130 ;
        RECT 75.300 199.070 75.620 199.130 ;
        RECT 77.155 199.070 77.445 199.115 ;
        RECT 75.300 198.930 77.445 199.070 ;
        RECT 75.300 198.870 75.620 198.930 ;
        RECT 77.155 198.885 77.445 198.930 ;
        RECT 91.400 198.870 91.720 199.130 ;
        RECT 92.320 198.870 92.640 199.130 ;
        RECT 96.015 199.070 96.305 199.115 ;
        RECT 104.740 199.070 105.060 199.130 ;
        RECT 107.975 199.070 108.265 199.115 ;
        RECT 92.870 198.930 95.770 199.070 ;
        RECT 29.315 198.590 36.890 198.730 ;
        RECT 29.315 198.545 29.605 198.590 ;
        RECT 40.340 198.530 40.660 198.790 ;
        RECT 46.320 198.730 46.640 198.790 ;
        RECT 57.820 198.730 58.140 198.790 ;
        RECT 58.295 198.730 58.585 198.775 ;
        RECT 63.800 198.730 64.120 198.790 ;
        RECT 69.320 198.730 69.640 198.790 ;
        RECT 44.110 198.590 46.640 198.730 ;
        RECT 22.375 198.390 22.665 198.435 ;
        RECT 23.565 198.390 23.855 198.435 ;
        RECT 26.085 198.390 26.375 198.435 ;
        RECT 40.430 198.390 40.570 198.530 ;
        RECT 44.110 198.435 44.250 198.590 ;
        RECT 46.320 198.530 46.640 198.590 ;
        RECT 49.630 198.590 52.990 198.730 ;
        RECT 22.375 198.250 26.375 198.390 ;
        RECT 22.375 198.205 22.665 198.250 ;
        RECT 23.565 198.205 23.855 198.250 ;
        RECT 26.085 198.205 26.375 198.250 ;
        RECT 28.930 198.250 40.570 198.390 ;
        RECT 28.930 198.110 29.070 198.250 ;
        RECT 21.495 198.050 21.785 198.095 ;
        RECT 25.160 198.050 25.480 198.110 ;
        RECT 21.495 197.910 25.480 198.050 ;
        RECT 21.495 197.865 21.785 197.910 ;
        RECT 25.160 197.850 25.480 197.910 ;
        RECT 28.840 197.850 29.160 198.110 ;
        RECT 29.775 198.050 30.065 198.095 ;
        RECT 29.775 197.910 31.370 198.050 ;
        RECT 29.775 197.865 30.065 197.910 ;
        RECT 22.860 197.755 23.180 197.770 ;
        RECT 22.830 197.525 23.180 197.755 ;
        RECT 22.860 197.510 23.180 197.525 ;
        RECT 26.080 197.710 26.400 197.770 ;
        RECT 29.850 197.710 29.990 197.865 ;
        RECT 26.080 197.570 29.990 197.710 ;
        RECT 26.080 197.510 26.400 197.570 ;
        RECT 28.380 197.170 28.700 197.430 ;
        RECT 30.680 197.170 31.000 197.430 ;
        RECT 31.230 197.370 31.370 197.910 ;
        RECT 31.600 197.850 31.920 198.110 ;
        RECT 32.520 197.850 32.840 198.110 ;
        RECT 33.070 198.095 33.210 198.250 ;
        RECT 44.035 198.205 44.325 198.435 ;
        RECT 44.495 198.390 44.785 198.435 ;
        RECT 45.860 198.390 46.180 198.450 ;
        RECT 44.495 198.250 46.180 198.390 ;
        RECT 44.495 198.205 44.785 198.250 ;
        RECT 45.860 198.190 46.180 198.250 ;
        RECT 32.995 198.050 33.285 198.095 ;
        RECT 33.455 198.050 33.745 198.095 ;
        RECT 32.995 197.910 33.745 198.050 ;
        RECT 32.995 197.865 33.285 197.910 ;
        RECT 33.455 197.865 33.745 197.910 ;
        RECT 33.900 198.050 34.220 198.110 ;
        RECT 34.375 198.050 34.665 198.095 ;
        RECT 33.900 197.910 38.270 198.050 ;
        RECT 33.900 197.850 34.220 197.910 ;
        RECT 34.375 197.865 34.665 197.910 ;
        RECT 32.060 197.710 32.380 197.770 ;
        RECT 35.295 197.710 35.585 197.755 ;
        RECT 36.515 197.710 36.805 197.755 ;
        RECT 32.060 197.570 33.210 197.710 ;
        RECT 32.060 197.510 32.380 197.570 ;
        RECT 32.520 197.370 32.840 197.430 ;
        RECT 31.230 197.230 32.840 197.370 ;
        RECT 33.070 197.370 33.210 197.570 ;
        RECT 35.295 197.570 36.805 197.710 ;
        RECT 35.295 197.525 35.585 197.570 ;
        RECT 36.515 197.525 36.805 197.570 ;
        RECT 37.595 197.525 37.885 197.755 ;
        RECT 38.130 197.710 38.270 197.910 ;
        RECT 38.960 197.850 39.280 198.110 ;
        RECT 40.355 198.050 40.645 198.095 ;
        RECT 40.800 198.050 41.120 198.110 ;
        RECT 42.655 198.050 42.945 198.095 ;
        RECT 40.355 197.910 42.945 198.050 ;
        RECT 40.355 197.865 40.645 197.910 ;
        RECT 40.800 197.850 41.120 197.910 ;
        RECT 42.655 197.865 42.945 197.910 ;
        RECT 43.100 198.050 43.420 198.110 ;
        RECT 49.630 198.095 49.770 198.590 ;
        RECT 50.460 198.190 50.780 198.450 ;
        RECT 48.635 198.050 48.925 198.095 ;
        RECT 43.100 197.910 48.925 198.050 ;
        RECT 41.260 197.710 41.580 197.770 ;
        RECT 38.130 197.570 41.580 197.710 ;
        RECT 37.670 197.370 37.810 197.525 ;
        RECT 41.260 197.510 41.580 197.570 ;
        RECT 33.070 197.230 37.810 197.370 ;
        RECT 42.730 197.370 42.870 197.865 ;
        RECT 43.100 197.850 43.420 197.910 ;
        RECT 48.635 197.865 48.925 197.910 ;
        RECT 49.555 197.865 49.845 198.095 ;
        RECT 50.015 198.050 50.305 198.095 ;
        RECT 50.550 198.050 50.690 198.190 ;
        RECT 51.395 198.050 51.685 198.095 ;
        RECT 52.300 198.050 52.620 198.110 ;
        RECT 50.015 197.910 50.690 198.050 ;
        RECT 51.010 197.910 52.620 198.050 ;
        RECT 52.850 198.050 52.990 198.590 ;
        RECT 53.310 198.590 56.210 198.730 ;
        RECT 53.310 198.435 53.450 198.590 ;
        RECT 53.235 198.205 53.525 198.435 ;
        RECT 53.695 198.390 53.985 198.435 ;
        RECT 55.520 198.390 55.840 198.450 ;
        RECT 53.695 198.250 55.840 198.390 ;
        RECT 56.070 198.390 56.210 198.590 ;
        RECT 57.820 198.590 58.585 198.730 ;
        RECT 57.820 198.530 58.140 198.590 ;
        RECT 58.295 198.545 58.585 198.590 ;
        RECT 58.830 198.590 64.120 198.730 ;
        RECT 58.830 198.390 58.970 198.590 ;
        RECT 63.800 198.530 64.120 198.590 ;
        RECT 66.650 198.590 69.640 198.730 ;
        RECT 56.070 198.250 58.970 198.390 ;
        RECT 53.695 198.205 53.985 198.250 ;
        RECT 55.520 198.190 55.840 198.250 ;
        RECT 60.580 198.190 60.900 198.450 ;
        RECT 61.975 198.390 62.265 198.435 ;
        RECT 66.650 198.390 66.790 198.590 ;
        RECT 69.320 198.530 69.640 198.590 ;
        RECT 70.740 198.730 71.030 198.775 ;
        RECT 72.840 198.730 73.130 198.775 ;
        RECT 74.410 198.730 74.700 198.775 ;
        RECT 92.870 198.730 93.010 198.930 ;
        RECT 70.740 198.590 74.700 198.730 ;
        RECT 70.740 198.545 71.030 198.590 ;
        RECT 72.840 198.545 73.130 198.590 ;
        RECT 74.410 198.545 74.700 198.590 ;
        RECT 91.490 198.590 93.010 198.730 ;
        RECT 61.975 198.250 66.790 198.390 ;
        RECT 61.975 198.205 62.265 198.250 ;
        RECT 67.020 198.190 67.340 198.450 ;
        RECT 71.135 198.390 71.425 198.435 ;
        RECT 72.325 198.390 72.615 198.435 ;
        RECT 74.845 198.390 75.135 198.435 ;
        RECT 71.135 198.250 75.135 198.390 ;
        RECT 71.135 198.205 71.425 198.250 ;
        RECT 72.325 198.205 72.615 198.250 ;
        RECT 74.845 198.205 75.135 198.250 ;
        RECT 52.850 197.910 53.450 198.050 ;
        RECT 50.015 197.865 50.305 197.910 ;
        RECT 45.400 197.510 45.720 197.770 ;
        RECT 46.320 197.510 46.640 197.770 ;
        RECT 48.710 197.710 48.850 197.865 ;
        RECT 51.010 197.710 51.150 197.910 ;
        RECT 51.395 197.865 51.685 197.910 ;
        RECT 52.300 197.850 52.620 197.910 ;
        RECT 48.710 197.570 51.150 197.710 ;
        RECT 53.310 197.710 53.450 197.910 ;
        RECT 54.140 197.850 54.460 198.110 ;
        RECT 54.615 198.050 54.905 198.095 ;
        RECT 55.060 198.050 55.380 198.110 ;
        RECT 54.615 197.910 55.380 198.050 ;
        RECT 54.615 197.865 54.905 197.910 ;
        RECT 55.060 197.850 55.380 197.910 ;
        RECT 57.360 197.850 57.680 198.110 ;
        RECT 59.200 198.050 59.520 198.110 ;
        RECT 63.355 198.050 63.645 198.095 ;
        RECT 59.200 197.910 63.645 198.050 ;
        RECT 59.200 197.850 59.520 197.910 ;
        RECT 63.355 197.865 63.645 197.910 ;
        RECT 65.180 197.850 65.500 198.110 ;
        RECT 65.640 197.850 65.960 198.110 ;
        RECT 68.860 197.850 69.180 198.110 ;
        RECT 69.780 197.850 70.100 198.110 ;
        RECT 70.255 197.865 70.545 198.095 ;
        RECT 71.590 197.865 71.880 198.095 ;
        RECT 78.520 198.050 78.840 198.110 ;
        RECT 73.780 197.910 78.840 198.050 ;
        RECT 56.915 197.710 57.205 197.755 ;
        RECT 53.310 197.570 57.205 197.710 ;
        RECT 56.915 197.525 57.205 197.570 ;
        RECT 58.295 197.710 58.585 197.755 ;
        RECT 58.295 197.570 62.650 197.710 ;
        RECT 58.295 197.525 58.585 197.570 ;
        RECT 45.490 197.370 45.630 197.510 ;
        RECT 42.730 197.230 45.630 197.370 ;
        RECT 46.780 197.370 47.100 197.430 ;
        RECT 47.255 197.370 47.545 197.415 ;
        RECT 46.780 197.230 47.545 197.370 ;
        RECT 32.520 197.170 32.840 197.230 ;
        RECT 46.780 197.170 47.100 197.230 ;
        RECT 47.255 197.185 47.545 197.230 ;
        RECT 52.315 197.370 52.605 197.415 ;
        RECT 53.220 197.370 53.540 197.430 ;
        RECT 52.315 197.230 53.540 197.370 ;
        RECT 52.315 197.185 52.605 197.230 ;
        RECT 53.220 197.170 53.540 197.230 ;
        RECT 55.535 197.370 55.825 197.415 ;
        RECT 56.440 197.370 56.760 197.430 ;
        RECT 55.535 197.230 56.760 197.370 ;
        RECT 55.535 197.185 55.825 197.230 ;
        RECT 56.440 197.170 56.760 197.230 ;
        RECT 61.040 197.170 61.360 197.430 ;
        RECT 62.510 197.415 62.650 197.570 ;
        RECT 62.435 197.185 62.725 197.415 ;
        RECT 69.320 197.170 69.640 197.430 ;
        RECT 70.330 197.370 70.470 197.865 ;
        RECT 71.160 197.710 71.480 197.770 ;
        RECT 71.710 197.710 71.850 197.865 ;
        RECT 71.160 197.570 71.850 197.710 ;
        RECT 71.160 197.510 71.480 197.570 ;
        RECT 73.780 197.370 73.920 197.910 ;
        RECT 78.520 197.850 78.840 197.910 ;
        RECT 84.960 197.850 85.280 198.110 ;
        RECT 86.355 197.865 86.645 198.095 ;
        RECT 86.430 197.710 86.570 197.865 ;
        RECT 89.100 197.850 89.420 198.110 ;
        RECT 90.035 197.865 90.325 198.095 ;
        RECT 89.575 197.710 89.865 197.755 ;
        RECT 86.430 197.570 89.865 197.710 ;
        RECT 90.110 197.710 90.250 197.865 ;
        RECT 90.480 197.850 90.800 198.110 ;
        RECT 91.490 198.095 91.630 198.590 ;
        RECT 94.620 198.530 94.940 198.790 ;
        RECT 95.630 198.730 95.770 198.930 ;
        RECT 96.015 198.930 105.060 199.070 ;
        RECT 96.015 198.885 96.305 198.930 ;
        RECT 104.740 198.870 105.060 198.930 ;
        RECT 105.290 198.930 108.265 199.070 ;
        RECT 99.680 198.730 100.000 198.790 ;
        RECT 105.290 198.730 105.430 198.930 ;
        RECT 107.975 198.885 108.265 198.930 ;
        RECT 108.420 198.730 108.740 198.790 ;
        RECT 95.630 198.590 100.000 198.730 ;
        RECT 99.680 198.530 100.000 198.590 ;
        RECT 103.910 198.590 105.430 198.730 ;
        RECT 107.130 198.590 108.740 198.730 ;
        RECT 94.710 198.390 94.850 198.530 ;
        RECT 96.000 198.390 96.320 198.450 ;
        RECT 92.870 198.250 94.850 198.390 ;
        RECT 95.170 198.250 96.320 198.390 ;
        RECT 92.870 198.095 93.010 198.250 ;
        RECT 91.415 197.865 91.705 198.095 ;
        RECT 92.795 197.865 93.085 198.095 ;
        RECT 93.255 197.865 93.545 198.095 ;
        RECT 93.715 198.050 94.005 198.095 ;
        RECT 94.160 198.050 94.480 198.110 ;
        RECT 93.715 197.910 94.480 198.050 ;
        RECT 93.715 197.865 94.005 197.910 ;
        RECT 93.330 197.710 93.470 197.865 ;
        RECT 94.160 197.850 94.480 197.910 ;
        RECT 94.635 198.050 94.925 198.095 ;
        RECT 95.170 198.050 95.310 198.250 ;
        RECT 96.000 198.190 96.320 198.250 ;
        RECT 100.140 198.390 100.460 198.450 ;
        RECT 103.910 198.390 104.050 198.590 ;
        RECT 107.130 198.390 107.270 198.590 ;
        RECT 108.420 198.530 108.740 198.590 ;
        RECT 100.140 198.250 104.050 198.390 ;
        RECT 100.140 198.190 100.460 198.250 ;
        RECT 94.635 197.910 95.310 198.050 ;
        RECT 95.540 198.050 95.860 198.110 ;
        RECT 96.935 198.050 97.225 198.095 ;
        RECT 95.540 197.910 97.225 198.050 ;
        RECT 94.635 197.865 94.925 197.910 ;
        RECT 95.540 197.850 95.860 197.910 ;
        RECT 96.935 197.865 97.225 197.910 ;
        RECT 97.395 198.050 97.685 198.095 ;
        RECT 98.300 198.050 98.620 198.110 ;
        RECT 97.395 197.910 98.620 198.050 ;
        RECT 97.395 197.865 97.685 197.910 ;
        RECT 98.300 197.850 98.620 197.910 ;
        RECT 98.760 197.850 99.080 198.110 ;
        RECT 99.235 198.050 99.525 198.095 ;
        RECT 101.060 198.050 101.380 198.110 ;
        RECT 102.900 198.095 103.220 198.110 ;
        RECT 103.910 198.095 104.050 198.250 ;
        RECT 104.830 198.250 107.270 198.390 ;
        RECT 107.500 198.390 107.820 198.450 ;
        RECT 113.035 198.390 113.325 198.435 ;
        RECT 107.500 198.250 113.325 198.390 ;
        RECT 104.830 198.095 104.970 198.250 ;
        RECT 107.500 198.190 107.820 198.250 ;
        RECT 113.035 198.205 113.325 198.250 ;
        RECT 99.235 197.910 101.380 198.050 ;
        RECT 99.235 197.865 99.525 197.910 ;
        RECT 101.060 197.850 101.380 197.910 ;
        RECT 102.890 197.865 103.220 198.095 ;
        RECT 103.835 197.865 104.125 198.095 ;
        RECT 104.750 197.865 105.040 198.095 ;
        RECT 105.215 197.865 105.505 198.095 ;
        RECT 102.900 197.850 103.220 197.865 ;
        RECT 97.840 197.710 98.160 197.770 ;
        RECT 100.600 197.710 100.920 197.770 ;
        RECT 90.110 197.570 90.710 197.710 ;
        RECT 93.330 197.570 94.850 197.710 ;
        RECT 89.575 197.525 89.865 197.570 ;
        RECT 70.330 197.230 73.920 197.370 ;
        RECT 84.040 197.170 84.360 197.430 ;
        RECT 85.880 197.170 86.200 197.430 ;
        RECT 90.570 197.370 90.710 197.570 ;
        RECT 94.710 197.430 94.850 197.570 ;
        RECT 97.840 197.570 100.920 197.710 ;
        RECT 97.840 197.510 98.160 197.570 ;
        RECT 100.600 197.510 100.920 197.570 ;
        RECT 94.160 197.370 94.480 197.430 ;
        RECT 90.570 197.230 94.480 197.370 ;
        RECT 94.160 197.170 94.480 197.230 ;
        RECT 94.620 197.170 94.940 197.430 ;
        RECT 95.555 197.370 95.845 197.415 ;
        RECT 96.000 197.370 96.320 197.430 ;
        RECT 95.555 197.230 96.320 197.370 ;
        RECT 95.555 197.185 95.845 197.230 ;
        RECT 96.000 197.170 96.320 197.230 ;
        RECT 100.140 197.370 100.460 197.430 ;
        RECT 101.150 197.370 101.290 197.850 ;
        RECT 101.520 197.510 101.840 197.770 ;
        RECT 103.375 197.525 103.665 197.755 ;
        RECT 105.290 197.710 105.430 197.865 ;
        RECT 105.660 197.850 105.980 198.110 ;
        RECT 106.580 198.050 106.900 198.110 ;
        RECT 107.975 198.050 108.265 198.095 ;
        RECT 106.580 197.910 108.265 198.050 ;
        RECT 106.580 197.850 106.900 197.910 ;
        RECT 107.975 197.865 108.265 197.910 ;
        RECT 108.895 197.865 109.185 198.095 ;
        RECT 106.135 197.710 106.425 197.755 ;
        RECT 108.970 197.710 109.110 197.865 ;
        RECT 117.160 197.850 117.480 198.110 ;
        RECT 123.155 198.050 123.445 198.095 ;
        RECT 124.520 198.050 124.840 198.110 ;
        RECT 123.155 197.910 124.840 198.050 ;
        RECT 123.155 197.865 123.445 197.910 ;
        RECT 124.520 197.850 124.840 197.910 ;
        RECT 124.980 197.850 125.300 198.110 ;
        RECT 105.290 197.570 106.425 197.710 ;
        RECT 106.135 197.525 106.425 197.570 ;
        RECT 106.670 197.570 109.110 197.710 ;
        RECT 112.115 197.710 112.405 197.755 ;
        RECT 118.080 197.710 118.400 197.770 ;
        RECT 112.115 197.570 118.400 197.710 ;
        RECT 100.140 197.230 101.290 197.370 ;
        RECT 100.140 197.170 100.460 197.230 ;
        RECT 101.980 197.170 102.300 197.430 ;
        RECT 102.440 197.370 102.760 197.430 ;
        RECT 103.450 197.370 103.590 197.525 ;
        RECT 105.200 197.370 105.520 197.430 ;
        RECT 106.670 197.370 106.810 197.570 ;
        RECT 112.115 197.525 112.405 197.570 ;
        RECT 118.080 197.510 118.400 197.570 ;
        RECT 123.615 197.525 123.905 197.755 ;
        RECT 124.075 197.710 124.365 197.755 ;
        RECT 126.820 197.710 127.140 197.770 ;
        RECT 124.075 197.570 127.140 197.710 ;
        RECT 124.075 197.525 124.365 197.570 ;
        RECT 102.440 197.230 106.810 197.370 ;
        RECT 102.440 197.170 102.760 197.230 ;
        RECT 105.200 197.170 105.520 197.230 ;
        RECT 110.260 197.170 110.580 197.430 ;
        RECT 112.575 197.370 112.865 197.415 ;
        RECT 114.415 197.370 114.705 197.415 ;
        RECT 112.575 197.230 114.705 197.370 ;
        RECT 112.575 197.185 112.865 197.230 ;
        RECT 114.415 197.185 114.705 197.230 ;
        RECT 122.220 197.170 122.540 197.430 ;
        RECT 123.690 197.370 123.830 197.525 ;
        RECT 126.820 197.510 127.140 197.570 ;
        RECT 131.880 197.370 132.200 197.430 ;
        RECT 123.690 197.230 132.200 197.370 ;
        RECT 131.880 197.170 132.200 197.230 ;
        RECT 17.270 196.550 146.990 197.030 ;
        RECT 19.195 196.350 19.485 196.395 ;
        RECT 21.480 196.350 21.800 196.410 ;
        RECT 19.195 196.210 21.800 196.350 ;
        RECT 19.195 196.165 19.485 196.210 ;
        RECT 21.480 196.150 21.800 196.210 ;
        RECT 25.160 196.150 25.480 196.410 ;
        RECT 27.475 196.350 27.765 196.395 ;
        RECT 28.840 196.350 29.160 196.410 ;
        RECT 43.100 196.350 43.420 196.410 ;
        RECT 27.475 196.210 29.160 196.350 ;
        RECT 27.475 196.165 27.765 196.210 ;
        RECT 28.840 196.150 29.160 196.210 ;
        RECT 37.670 196.210 43.420 196.350 ;
        RECT 23.780 196.010 24.100 196.070 ;
        RECT 24.760 196.010 25.050 196.055 ;
        RECT 23.780 195.870 25.050 196.010 ;
        RECT 23.780 195.810 24.100 195.870 ;
        RECT 24.760 195.825 25.050 195.870 ;
        RECT 25.250 195.670 25.390 196.150 ;
        RECT 27.935 196.010 28.225 196.055 ;
        RECT 31.600 196.010 31.920 196.070 ;
        RECT 37.670 196.010 37.810 196.210 ;
        RECT 43.100 196.150 43.420 196.210 ;
        RECT 51.840 196.150 52.160 196.410 ;
        RECT 54.140 196.150 54.460 196.410 ;
        RECT 54.600 196.150 54.920 196.410 ;
        RECT 55.060 196.350 55.380 196.410 ;
        RECT 60.580 196.350 60.900 196.410 ;
        RECT 55.060 196.210 60.900 196.350 ;
        RECT 55.060 196.150 55.380 196.210 ;
        RECT 27.935 195.870 31.920 196.010 ;
        RECT 27.935 195.825 28.225 195.870 ;
        RECT 31.600 195.810 31.920 195.870 ;
        RECT 33.530 195.870 37.810 196.010 ;
        RECT 26.095 195.670 26.385 195.715 ;
        RECT 25.250 195.530 26.385 195.670 ;
        RECT 26.095 195.485 26.385 195.530 ;
        RECT 28.380 195.670 28.700 195.730 ;
        RECT 33.530 195.715 33.670 195.870 ;
        RECT 28.380 195.530 32.290 195.670 ;
        RECT 28.380 195.470 28.700 195.530 ;
        RECT 21.505 195.330 21.795 195.375 ;
        RECT 24.025 195.330 24.315 195.375 ;
        RECT 25.215 195.330 25.505 195.375 ;
        RECT 21.505 195.190 25.505 195.330 ;
        RECT 21.505 195.145 21.795 195.190 ;
        RECT 24.025 195.145 24.315 195.190 ;
        RECT 25.215 195.145 25.505 195.190 ;
        RECT 28.840 195.330 29.160 195.390 ;
        RECT 30.695 195.330 30.985 195.375 ;
        RECT 28.840 195.190 30.985 195.330 ;
        RECT 28.840 195.130 29.160 195.190 ;
        RECT 30.695 195.145 30.985 195.190 ;
        RECT 31.140 195.130 31.460 195.390 ;
        RECT 32.150 195.375 32.290 195.530 ;
        RECT 33.455 195.485 33.745 195.715 ;
        RECT 34.375 195.670 34.665 195.715 ;
        RECT 35.740 195.670 36.060 195.730 ;
        RECT 34.375 195.530 36.060 195.670 ;
        RECT 34.375 195.485 34.665 195.530 ;
        RECT 31.615 195.145 31.905 195.375 ;
        RECT 32.075 195.330 32.365 195.375 ;
        RECT 34.450 195.330 34.590 195.485 ;
        RECT 35.740 195.470 36.060 195.530 ;
        RECT 37.120 195.470 37.440 195.730 ;
        RECT 37.670 195.715 37.810 195.870 ;
        RECT 39.895 196.010 40.185 196.055 ;
        RECT 45.415 196.010 45.705 196.055 ;
        RECT 39.895 195.870 45.705 196.010 ;
        RECT 39.895 195.825 40.185 195.870 ;
        RECT 45.415 195.825 45.705 195.870 ;
        RECT 46.780 195.810 47.100 196.070 ;
        RECT 53.680 196.010 54.000 196.070 ;
        RECT 51.010 195.870 54.000 196.010 ;
        RECT 51.010 195.730 51.150 195.870 ;
        RECT 53.680 195.810 54.000 195.870 ;
        RECT 37.595 195.670 37.885 195.715 ;
        RECT 38.500 195.670 38.820 195.730 ;
        RECT 37.595 195.530 38.820 195.670 ;
        RECT 37.595 195.485 37.885 195.530 ;
        RECT 38.500 195.470 38.820 195.530 ;
        RECT 38.975 195.670 39.265 195.715 ;
        RECT 39.420 195.670 39.740 195.730 ;
        RECT 38.975 195.530 39.740 195.670 ;
        RECT 38.975 195.485 39.265 195.530 ;
        RECT 39.420 195.470 39.740 195.530 ;
        RECT 40.340 195.470 40.660 195.730 ;
        RECT 40.815 195.485 41.105 195.715 ;
        RECT 41.260 195.670 41.580 195.730 ;
        RECT 43.575 195.670 43.865 195.715 ;
        RECT 41.260 195.530 43.865 195.670 ;
        RECT 39.880 195.330 40.200 195.390 ;
        RECT 32.075 195.190 34.590 195.330 ;
        RECT 35.370 195.190 40.200 195.330 ;
        RECT 40.890 195.330 41.030 195.485 ;
        RECT 41.260 195.470 41.580 195.530 ;
        RECT 43.575 195.485 43.865 195.530 ;
        RECT 44.345 195.670 44.635 195.715 ;
        RECT 44.940 195.670 45.260 195.730 ;
        RECT 45.875 195.670 46.165 195.715 ;
        RECT 44.345 195.485 44.710 195.670 ;
        RECT 43.100 195.330 43.420 195.390 ;
        RECT 40.890 195.190 43.420 195.330 ;
        RECT 44.570 195.330 44.710 195.485 ;
        RECT 44.940 195.530 46.165 195.670 ;
        RECT 44.940 195.470 45.260 195.530 ;
        RECT 45.875 195.485 46.165 195.530 ;
        RECT 50.920 195.470 51.240 195.730 ;
        RECT 51.855 195.485 52.145 195.715 ;
        RECT 46.320 195.330 46.640 195.390 ;
        RECT 44.570 195.190 46.640 195.330 ;
        RECT 51.930 195.330 52.070 195.485 ;
        RECT 52.300 195.470 52.620 195.730 ;
        RECT 55.520 195.470 55.840 195.730 ;
        RECT 55.995 195.670 56.285 195.715 ;
        RECT 56.900 195.670 57.220 195.730 ;
        RECT 55.995 195.530 57.220 195.670 ;
        RECT 55.995 195.485 56.285 195.530 ;
        RECT 56.900 195.470 57.220 195.530 ;
        RECT 57.360 195.470 57.680 195.730 ;
        RECT 58.830 195.715 58.970 196.210 ;
        RECT 60.580 196.150 60.900 196.210 ;
        RECT 61.040 196.150 61.360 196.410 ;
        RECT 71.160 196.150 71.480 196.410 ;
        RECT 78.520 196.150 78.840 196.410 ;
        RECT 85.880 196.350 86.200 196.410 ;
        RECT 87.735 196.350 88.025 196.395 ;
        RECT 90.480 196.350 90.800 196.410 ;
        RECT 85.880 196.210 90.800 196.350 ;
        RECT 85.880 196.150 86.200 196.210 ;
        RECT 87.735 196.165 88.025 196.210 ;
        RECT 90.480 196.150 90.800 196.210 ;
        RECT 98.760 196.350 99.080 196.410 ;
        RECT 100.615 196.350 100.905 196.395 ;
        RECT 98.760 196.210 100.905 196.350 ;
        RECT 98.760 196.150 99.080 196.210 ;
        RECT 100.615 196.165 100.905 196.210 ;
        RECT 101.060 196.350 101.380 196.410 ;
        RECT 103.820 196.350 104.140 196.410 ;
        RECT 104.295 196.350 104.585 196.395 ;
        RECT 101.060 196.210 103.590 196.350 ;
        RECT 101.060 196.150 101.380 196.210 ;
        RECT 60.120 196.010 60.440 196.070 ;
        RECT 61.975 196.010 62.265 196.055 ;
        RECT 60.120 195.870 62.265 196.010 ;
        RECT 60.120 195.810 60.440 195.870 ;
        RECT 61.975 195.825 62.265 195.870 ;
        RECT 72.540 195.810 72.860 196.070 ;
        RECT 78.610 196.010 78.750 196.150 ;
        RECT 82.170 196.010 82.460 196.055 ;
        RECT 84.040 196.010 84.360 196.070 ;
        RECT 78.610 195.870 80.130 196.010 ;
        RECT 57.835 195.485 58.125 195.715 ;
        RECT 58.755 195.485 59.045 195.715 ;
        RECT 52.775 195.330 53.065 195.375 ;
        RECT 57.910 195.330 58.050 195.485 ;
        RECT 59.200 195.470 59.520 195.730 ;
        RECT 59.660 195.470 59.980 195.730 ;
        RECT 61.500 195.470 61.820 195.730 ;
        RECT 62.895 195.485 63.185 195.715 ;
        RECT 69.320 195.670 69.640 195.730 ;
        RECT 71.175 195.670 71.465 195.715 ;
        RECT 69.320 195.530 71.465 195.670 ;
        RECT 61.040 195.330 61.360 195.390 ;
        RECT 51.930 195.190 56.210 195.330 ;
        RECT 57.910 195.190 61.360 195.330 ;
        RECT 32.075 195.145 32.365 195.190 ;
        RECT 21.940 194.990 22.230 195.035 ;
        RECT 23.510 194.990 23.800 195.035 ;
        RECT 25.610 194.990 25.900 195.035 ;
        RECT 21.940 194.850 25.900 194.990 ;
        RECT 21.940 194.805 22.230 194.850 ;
        RECT 23.510 194.805 23.800 194.850 ;
        RECT 25.610 194.805 25.900 194.850 ;
        RECT 29.315 194.990 29.605 195.035 ;
        RECT 31.690 194.990 31.830 195.145 ;
        RECT 32.520 194.990 32.840 195.050 ;
        RECT 34.820 194.990 35.140 195.050 ;
        RECT 35.370 195.035 35.510 195.190 ;
        RECT 39.880 195.130 40.200 195.190 ;
        RECT 43.100 195.130 43.420 195.190 ;
        RECT 46.320 195.130 46.640 195.190 ;
        RECT 52.775 195.145 53.065 195.190 ;
        RECT 56.070 195.050 56.210 195.190 ;
        RECT 61.040 195.130 61.360 195.190 ;
        RECT 29.315 194.850 35.140 194.990 ;
        RECT 29.315 194.805 29.605 194.850 ;
        RECT 32.520 194.790 32.840 194.850 ;
        RECT 34.820 194.790 35.140 194.850 ;
        RECT 35.295 194.805 35.585 195.035 ;
        RECT 36.215 194.990 36.505 195.035 ;
        RECT 40.800 194.990 41.120 195.050 ;
        RECT 36.215 194.850 41.120 194.990 ;
        RECT 36.215 194.805 36.505 194.850 ;
        RECT 40.800 194.790 41.120 194.850 ;
        RECT 55.980 194.790 56.300 195.050 ;
        RECT 57.820 194.990 58.140 195.050 ;
        RECT 62.970 194.990 63.110 195.485 ;
        RECT 69.320 195.470 69.640 195.530 ;
        RECT 71.175 195.485 71.465 195.530 ;
        RECT 71.635 195.670 71.925 195.715 ;
        RECT 73.460 195.670 73.780 195.730 ;
        RECT 79.990 195.715 80.130 195.870 ;
        RECT 82.170 195.870 84.360 196.010 ;
        RECT 82.170 195.825 82.460 195.870 ;
        RECT 84.040 195.810 84.360 195.870 ;
        RECT 99.235 196.010 99.525 196.055 ;
        RECT 102.440 196.010 102.760 196.070 ;
        RECT 99.235 195.870 102.760 196.010 ;
        RECT 103.450 196.010 103.590 196.210 ;
        RECT 103.820 196.210 104.585 196.350 ;
        RECT 103.820 196.150 104.140 196.210 ;
        RECT 104.295 196.165 104.585 196.210 ;
        RECT 105.200 196.150 105.520 196.410 ;
        RECT 120.840 196.150 121.160 196.410 ;
        RECT 123.155 196.350 123.445 196.395 ;
        RECT 125.915 196.350 126.205 196.395 ;
        RECT 127.280 196.350 127.600 196.410 ;
        RECT 123.155 196.210 127.600 196.350 ;
        RECT 123.155 196.165 123.445 196.210 ;
        RECT 125.915 196.165 126.205 196.210 ;
        RECT 127.280 196.150 127.600 196.210 ;
        RECT 108.850 196.010 109.140 196.055 ;
        RECT 110.260 196.010 110.580 196.070 ;
        RECT 103.450 195.870 104.970 196.010 ;
        RECT 99.235 195.825 99.525 195.870 ;
        RECT 102.440 195.810 102.760 195.870 ;
        RECT 71.635 195.530 73.780 195.670 ;
        RECT 71.635 195.485 71.925 195.530 ;
        RECT 73.460 195.470 73.780 195.530 ;
        RECT 78.635 195.670 78.925 195.715 ;
        RECT 79.915 195.670 80.205 195.715 ;
        RECT 80.835 195.670 81.125 195.715 ;
        RECT 78.635 195.530 79.670 195.670 ;
        RECT 78.635 195.485 78.925 195.530 ;
        RECT 75.325 195.330 75.615 195.375 ;
        RECT 77.845 195.330 78.135 195.375 ;
        RECT 79.035 195.330 79.325 195.375 ;
        RECT 75.325 195.190 79.325 195.330 ;
        RECT 79.530 195.330 79.670 195.530 ;
        RECT 79.915 195.530 81.125 195.670 ;
        RECT 79.915 195.485 80.205 195.530 ;
        RECT 80.835 195.485 81.125 195.530 ;
        RECT 97.855 195.670 98.145 195.715 ;
        RECT 98.300 195.670 98.620 195.730 ;
        RECT 97.855 195.530 98.620 195.670 ;
        RECT 97.855 195.485 98.145 195.530 ;
        RECT 98.300 195.470 98.620 195.530 ;
        RECT 98.760 195.470 99.080 195.730 ;
        RECT 99.695 195.670 99.985 195.715 ;
        RECT 101.520 195.670 101.840 195.730 ;
        RECT 99.695 195.530 101.840 195.670 ;
        RECT 99.695 195.485 99.985 195.530 ;
        RECT 101.520 195.470 101.840 195.530 ;
        RECT 101.980 195.470 102.300 195.730 ;
        RECT 104.830 195.715 104.970 195.870 ;
        RECT 108.850 195.870 110.580 196.010 ;
        RECT 108.850 195.825 109.140 195.870 ;
        RECT 110.260 195.810 110.580 195.870 ;
        RECT 123.600 196.010 123.920 196.070 ;
        RECT 123.600 195.870 133.030 196.010 ;
        RECT 123.600 195.810 123.920 195.870 ;
        RECT 102.915 195.660 103.205 195.715 ;
        RECT 103.450 195.660 104.510 195.670 ;
        RECT 102.915 195.530 104.510 195.660 ;
        RECT 102.915 195.520 103.590 195.530 ;
        RECT 102.915 195.485 103.205 195.520 ;
        RECT 81.715 195.330 82.005 195.375 ;
        RECT 82.905 195.330 83.195 195.375 ;
        RECT 85.425 195.330 85.715 195.375 ;
        RECT 79.530 195.190 81.050 195.330 ;
        RECT 75.325 195.145 75.615 195.190 ;
        RECT 77.845 195.145 78.135 195.190 ;
        RECT 79.035 195.145 79.325 195.190 ;
        RECT 67.020 194.990 67.340 195.050 ;
        RECT 57.820 194.850 63.110 194.990 ;
        RECT 63.430 194.850 67.340 194.990 ;
        RECT 57.820 194.790 58.140 194.850 ;
        RECT 26.080 194.650 26.400 194.710 ;
        RECT 26.555 194.650 26.845 194.695 ;
        RECT 26.080 194.510 26.845 194.650 ;
        RECT 26.080 194.450 26.400 194.510 ;
        RECT 26.555 194.465 26.845 194.510 ;
        RECT 27.460 194.650 27.780 194.710 ;
        RECT 29.775 194.650 30.065 194.695 ;
        RECT 27.460 194.510 30.065 194.650 ;
        RECT 27.460 194.450 27.780 194.510 ;
        RECT 29.775 194.465 30.065 194.510 ;
        RECT 31.140 194.650 31.460 194.710 ;
        RECT 33.455 194.650 33.745 194.695 ;
        RECT 37.120 194.650 37.440 194.710 ;
        RECT 31.140 194.510 37.440 194.650 ;
        RECT 31.140 194.450 31.460 194.510 ;
        RECT 33.455 194.465 33.745 194.510 ;
        RECT 37.120 194.450 37.440 194.510 ;
        RECT 38.515 194.650 38.805 194.695 ;
        RECT 40.340 194.650 40.660 194.710 ;
        RECT 38.515 194.510 40.660 194.650 ;
        RECT 38.515 194.465 38.805 194.510 ;
        RECT 40.340 194.450 40.660 194.510 ;
        RECT 41.735 194.650 42.025 194.695 ;
        RECT 42.640 194.650 42.960 194.710 ;
        RECT 41.735 194.510 42.960 194.650 ;
        RECT 41.735 194.465 42.025 194.510 ;
        RECT 42.640 194.450 42.960 194.510 ;
        RECT 50.460 194.650 50.780 194.710 ;
        RECT 52.315 194.650 52.605 194.695 ;
        RECT 50.460 194.510 52.605 194.650 ;
        RECT 50.460 194.450 50.780 194.510 ;
        RECT 52.315 194.465 52.605 194.510 ;
        RECT 56.915 194.650 57.205 194.695 ;
        RECT 63.430 194.650 63.570 194.850 ;
        RECT 67.020 194.790 67.340 194.850 ;
        RECT 75.760 194.990 76.050 195.035 ;
        RECT 77.330 194.990 77.620 195.035 ;
        RECT 79.430 194.990 79.720 195.035 ;
        RECT 75.760 194.850 79.720 194.990 ;
        RECT 75.760 194.805 76.050 194.850 ;
        RECT 77.330 194.805 77.620 194.850 ;
        RECT 79.430 194.805 79.720 194.850 ;
        RECT 56.915 194.510 63.570 194.650 ;
        RECT 56.915 194.465 57.205 194.510 ;
        RECT 63.800 194.450 64.120 194.710 ;
        RECT 69.780 194.650 70.100 194.710 ;
        RECT 73.015 194.650 73.305 194.695 ;
        RECT 69.780 194.510 73.305 194.650 ;
        RECT 80.910 194.650 81.050 195.190 ;
        RECT 81.715 195.190 85.715 195.330 ;
        RECT 81.715 195.145 82.005 195.190 ;
        RECT 82.905 195.145 83.195 195.190 ;
        RECT 85.425 195.145 85.715 195.190 ;
        RECT 100.600 195.330 100.920 195.390 ;
        RECT 102.455 195.330 102.745 195.375 ;
        RECT 103.375 195.330 103.665 195.375 ;
        RECT 100.600 195.190 102.745 195.330 ;
        RECT 100.600 195.130 100.920 195.190 ;
        RECT 102.455 195.145 102.745 195.190 ;
        RECT 102.990 195.190 103.665 195.330 ;
        RECT 104.370 195.330 104.510 195.530 ;
        RECT 104.755 195.485 105.045 195.715 ;
        RECT 107.515 195.670 107.805 195.715 ;
        RECT 107.960 195.670 108.280 195.730 ;
        RECT 107.515 195.530 108.280 195.670 ;
        RECT 107.515 195.485 107.805 195.530 ;
        RECT 107.960 195.470 108.280 195.530 ;
        RECT 122.695 195.670 122.985 195.715 ;
        RECT 125.440 195.670 125.760 195.730 ;
        RECT 122.695 195.530 125.760 195.670 ;
        RECT 122.695 195.485 122.985 195.530 ;
        RECT 125.440 195.470 125.760 195.530 ;
        RECT 131.535 195.670 131.825 195.715 ;
        RECT 132.340 195.670 132.660 195.730 ;
        RECT 132.890 195.715 133.030 195.870 ;
        RECT 131.535 195.530 132.660 195.670 ;
        RECT 131.535 195.485 131.825 195.530 ;
        RECT 132.340 195.470 132.660 195.530 ;
        RECT 132.815 195.485 133.105 195.715 ;
        RECT 134.180 195.470 134.500 195.730 ;
        RECT 106.580 195.330 106.900 195.390 ;
        RECT 104.370 195.190 106.900 195.330 ;
        RECT 81.320 194.990 81.610 195.035 ;
        RECT 83.420 194.990 83.710 195.035 ;
        RECT 84.990 194.990 85.280 195.035 ;
        RECT 81.320 194.850 85.280 194.990 ;
        RECT 81.320 194.805 81.610 194.850 ;
        RECT 83.420 194.805 83.710 194.850 ;
        RECT 84.990 194.805 85.280 194.850 ;
        RECT 82.200 194.650 82.520 194.710 ;
        RECT 80.910 194.510 82.520 194.650 ;
        RECT 102.990 194.650 103.130 195.190 ;
        RECT 103.375 195.145 103.665 195.190 ;
        RECT 106.580 195.130 106.900 195.190 ;
        RECT 108.395 195.330 108.685 195.375 ;
        RECT 109.585 195.330 109.875 195.375 ;
        RECT 112.105 195.330 112.395 195.375 ;
        RECT 108.395 195.190 112.395 195.330 ;
        RECT 108.395 195.145 108.685 195.190 ;
        RECT 109.585 195.145 109.875 195.190 ;
        RECT 112.105 195.145 112.395 195.190 ;
        RECT 120.840 195.330 121.160 195.390 ;
        RECT 123.615 195.330 123.905 195.375 ;
        RECT 120.840 195.190 123.905 195.330 ;
        RECT 120.840 195.130 121.160 195.190 ;
        RECT 123.615 195.145 123.905 195.190 ;
        RECT 128.225 195.330 128.515 195.375 ;
        RECT 130.745 195.330 131.035 195.375 ;
        RECT 131.935 195.330 132.225 195.375 ;
        RECT 128.225 195.190 132.225 195.330 ;
        RECT 128.225 195.145 128.515 195.190 ;
        RECT 130.745 195.145 131.035 195.190 ;
        RECT 131.935 195.145 132.225 195.190 ;
        RECT 108.000 194.990 108.290 195.035 ;
        RECT 110.100 194.990 110.390 195.035 ;
        RECT 111.670 194.990 111.960 195.035 ;
        RECT 108.000 194.850 111.960 194.990 ;
        RECT 108.000 194.805 108.290 194.850 ;
        RECT 110.100 194.805 110.390 194.850 ;
        RECT 111.670 194.805 111.960 194.850 ;
        RECT 128.660 194.990 128.950 195.035 ;
        RECT 130.230 194.990 130.520 195.035 ;
        RECT 132.330 194.990 132.620 195.035 ;
        RECT 128.660 194.850 132.620 194.990 ;
        RECT 128.660 194.805 128.950 194.850 ;
        RECT 130.230 194.805 130.520 194.850 ;
        RECT 132.330 194.805 132.620 194.850 ;
        RECT 132.800 194.990 133.120 195.050 ;
        RECT 133.275 194.990 133.565 195.035 ;
        RECT 132.800 194.850 133.565 194.990 ;
        RECT 132.800 194.790 133.120 194.850 ;
        RECT 133.275 194.805 133.565 194.850 ;
        RECT 114.415 194.650 114.705 194.695 ;
        RECT 117.160 194.650 117.480 194.710 ;
        RECT 102.990 194.510 117.480 194.650 ;
        RECT 69.780 194.450 70.100 194.510 ;
        RECT 73.015 194.465 73.305 194.510 ;
        RECT 82.200 194.450 82.520 194.510 ;
        RECT 114.415 194.465 114.705 194.510 ;
        RECT 117.160 194.450 117.480 194.510 ;
        RECT 17.270 193.830 146.990 194.310 ;
        RECT 22.860 193.430 23.180 193.690 ;
        RECT 23.795 193.445 24.085 193.675 ;
        RECT 23.870 193.290 24.010 193.445 ;
        RECT 27.000 193.430 27.320 193.690 ;
        RECT 35.280 193.630 35.600 193.690 ;
        RECT 38.960 193.630 39.280 193.690 ;
        RECT 35.280 193.490 39.280 193.630 ;
        RECT 35.280 193.430 35.600 193.490 ;
        RECT 38.960 193.430 39.280 193.490 ;
        RECT 59.215 193.630 59.505 193.675 ;
        RECT 61.500 193.630 61.820 193.690 ;
        RECT 96.460 193.630 96.780 193.690 ;
        RECT 99.680 193.630 100.000 193.690 ;
        RECT 59.215 193.490 61.820 193.630 ;
        RECT 59.215 193.445 59.505 193.490 ;
        RECT 61.500 193.430 61.820 193.490 ;
        RECT 95.170 193.490 100.000 193.630 ;
        RECT 43.100 193.290 43.420 193.350 ;
        RECT 23.870 193.150 29.070 193.290 ;
        RECT 26.080 192.950 26.400 193.010 ;
        RECT 28.930 192.995 29.070 193.150 ;
        RECT 41.810 193.150 43.420 193.290 ;
        RECT 28.855 192.950 29.145 192.995 ;
        RECT 38.975 192.950 39.265 192.995 ;
        RECT 41.810 192.950 41.950 193.150 ;
        RECT 43.100 193.090 43.420 193.150 ;
        RECT 45.860 193.290 46.180 193.350 ;
        RECT 50.920 193.290 51.240 193.350 ;
        RECT 45.860 193.150 51.240 193.290 ;
        RECT 45.860 193.090 46.180 193.150 ;
        RECT 50.920 193.090 51.240 193.150 ;
        RECT 52.300 193.290 52.620 193.350 ;
        RECT 52.775 193.290 53.065 193.335 ;
        RECT 55.520 193.290 55.840 193.350 ;
        RECT 69.780 193.290 70.100 193.350 ;
        RECT 52.300 193.150 58.510 193.290 ;
        RECT 52.300 193.090 52.620 193.150 ;
        RECT 52.775 193.105 53.065 193.150 ;
        RECT 55.520 193.090 55.840 193.150 ;
        RECT 43.575 192.950 43.865 192.995 ;
        RECT 26.080 192.810 28.610 192.950 ;
        RECT 26.080 192.750 26.400 192.810 ;
        RECT 27.460 192.610 27.780 192.670 ;
        RECT 28.470 192.655 28.610 192.810 ;
        RECT 28.855 192.810 29.255 192.950 ;
        RECT 38.975 192.810 41.490 192.950 ;
        RECT 41.810 192.810 43.865 192.950 ;
        RECT 28.855 192.765 29.145 192.810 ;
        RECT 38.975 192.765 39.265 192.810 ;
        RECT 24.330 192.470 27.780 192.610 ;
        RECT 23.715 192.270 24.005 192.315 ;
        RECT 24.330 192.270 24.470 192.470 ;
        RECT 27.460 192.410 27.780 192.470 ;
        RECT 28.395 192.425 28.685 192.655 ;
        RECT 35.740 192.610 36.060 192.670 ;
        RECT 35.740 192.470 38.270 192.610 ;
        RECT 35.740 192.410 36.060 192.470 ;
        RECT 23.715 192.130 24.470 192.270 ;
        RECT 24.700 192.270 25.020 192.330 ;
        RECT 27.935 192.270 28.225 192.315 ;
        RECT 32.060 192.270 32.380 192.330 ;
        RECT 24.700 192.130 32.380 192.270 ;
        RECT 23.715 192.085 24.005 192.130 ;
        RECT 24.700 192.070 25.020 192.130 ;
        RECT 27.935 192.085 28.225 192.130 ;
        RECT 32.060 192.070 32.380 192.130 ;
        RECT 37.120 192.270 37.440 192.330 ;
        RECT 37.595 192.270 37.885 192.315 ;
        RECT 37.120 192.130 37.885 192.270 ;
        RECT 38.130 192.270 38.270 192.470 ;
        RECT 38.500 192.410 38.820 192.670 ;
        RECT 39.420 192.655 39.740 192.670 ;
        RECT 39.420 192.610 39.750 192.655 ;
        RECT 39.420 192.470 40.110 192.610 ;
        RECT 39.420 192.425 39.750 192.470 ;
        RECT 39.420 192.410 39.740 192.425 ;
        RECT 38.975 192.270 39.265 192.315 ;
        RECT 38.130 192.130 39.265 192.270 ;
        RECT 39.970 192.270 40.110 192.470 ;
        RECT 40.340 192.410 40.660 192.670 ;
        RECT 41.350 192.655 41.490 192.810 ;
        RECT 43.575 192.765 43.865 192.810 ;
        RECT 44.955 192.950 45.245 192.995 ;
        RECT 50.015 192.950 50.305 192.995 ;
        RECT 57.360 192.950 57.680 193.010 ;
        RECT 44.955 192.810 50.305 192.950 ;
        RECT 44.955 192.765 45.245 192.810 ;
        RECT 50.015 192.765 50.305 192.810 ;
        RECT 51.010 192.810 57.680 192.950 ;
        RECT 41.275 192.425 41.565 192.655 ;
        RECT 42.180 192.610 42.500 192.670 ;
        RECT 42.655 192.610 42.945 192.655 ;
        RECT 42.180 192.470 42.945 192.610 ;
        RECT 42.180 192.410 42.500 192.470 ;
        RECT 42.655 192.425 42.945 192.470 ;
        RECT 46.320 192.410 46.640 192.670 ;
        RECT 51.010 192.655 51.150 192.810 ;
        RECT 57.360 192.750 57.680 192.810 ;
        RECT 50.935 192.425 51.225 192.655 ;
        RECT 40.800 192.270 41.120 192.330 ;
        RECT 45.860 192.270 46.180 192.330 ;
        RECT 39.970 192.130 46.180 192.270 ;
        RECT 37.120 192.070 37.440 192.130 ;
        RECT 37.595 192.085 37.885 192.130 ;
        RECT 38.975 192.085 39.265 192.130 ;
        RECT 40.800 192.070 41.120 192.130 ;
        RECT 45.860 192.070 46.180 192.130 ;
        RECT 25.620 191.930 25.940 191.990 ;
        RECT 26.095 191.930 26.385 191.975 ;
        RECT 25.620 191.790 26.385 191.930 ;
        RECT 25.620 191.730 25.940 191.790 ;
        RECT 26.095 191.745 26.385 191.790 ;
        RECT 26.935 191.930 27.225 191.975 ;
        RECT 30.680 191.930 31.000 191.990 ;
        RECT 26.935 191.790 31.000 191.930 ;
        RECT 26.935 191.745 27.225 191.790 ;
        RECT 30.680 191.730 31.000 191.790 ;
        RECT 41.260 191.730 41.580 191.990 ;
        RECT 41.720 191.730 42.040 191.990 ;
        RECT 44.940 191.930 45.260 191.990 ;
        RECT 51.010 191.930 51.150 192.425 ;
        RECT 56.440 192.410 56.760 192.670 ;
        RECT 56.900 192.610 57.220 192.670 ;
        RECT 58.370 192.655 58.510 193.150 ;
        RECT 59.750 193.150 70.100 193.290 ;
        RECT 57.835 192.610 58.125 192.655 ;
        RECT 56.900 192.470 58.125 192.610 ;
        RECT 56.900 192.410 57.220 192.470 ;
        RECT 57.835 192.425 58.125 192.470 ;
        RECT 58.295 192.425 58.585 192.655 ;
        RECT 54.600 192.270 54.920 192.330 ;
        RECT 57.375 192.270 57.665 192.315 ;
        RECT 54.600 192.130 57.665 192.270 ;
        RECT 57.910 192.270 58.050 192.425 ;
        RECT 59.750 192.270 59.890 193.150 ;
        RECT 69.780 193.090 70.100 193.150 ;
        RECT 73.460 193.090 73.780 193.350 ;
        RECT 75.315 193.290 75.605 193.335 ;
        RECT 81.740 193.290 82.060 193.350 ;
        RECT 75.315 193.150 82.060 193.290 ;
        RECT 75.315 193.105 75.605 193.150 ;
        RECT 81.740 193.090 82.060 193.150 ;
        RECT 62.880 192.950 63.200 193.010 ;
        RECT 60.670 192.810 63.200 192.950 ;
        RECT 60.120 192.610 60.440 192.670 ;
        RECT 60.670 192.655 60.810 192.810 ;
        RECT 62.880 192.750 63.200 192.810 ;
        RECT 73.015 192.950 73.305 192.995 ;
        RECT 73.550 192.950 73.690 193.090 ;
        RECT 73.015 192.810 73.690 192.950 ;
        RECT 77.615 192.950 77.905 192.995 ;
        RECT 81.280 192.950 81.600 193.010 ;
        RECT 95.170 192.995 95.310 193.490 ;
        RECT 96.460 193.430 96.780 193.490 ;
        RECT 99.680 193.430 100.000 193.490 ;
        RECT 101.520 193.630 101.840 193.690 ;
        RECT 101.995 193.630 102.285 193.675 ;
        RECT 101.520 193.490 102.285 193.630 ;
        RECT 101.520 193.430 101.840 193.490 ;
        RECT 101.995 193.445 102.285 193.490 ;
        RECT 102.900 193.630 103.220 193.690 ;
        RECT 114.860 193.630 115.180 193.690 ;
        RECT 102.900 193.490 115.180 193.630 ;
        RECT 102.900 193.430 103.220 193.490 ;
        RECT 114.860 193.430 115.180 193.490 ;
        RECT 118.080 193.430 118.400 193.690 ;
        RECT 124.980 193.630 125.300 193.690 ;
        RECT 125.455 193.630 125.745 193.675 ;
        RECT 124.980 193.490 125.745 193.630 ;
        RECT 124.980 193.430 125.300 193.490 ;
        RECT 125.455 193.445 125.745 193.490 ;
        RECT 131.880 193.430 132.200 193.690 ;
        RECT 132.340 193.630 132.660 193.690 ;
        RECT 133.735 193.630 134.025 193.675 ;
        RECT 132.340 193.490 134.025 193.630 ;
        RECT 132.340 193.430 132.660 193.490 ;
        RECT 133.735 193.445 134.025 193.490 ;
        RECT 95.580 193.290 95.870 193.335 ;
        RECT 97.680 193.290 97.970 193.335 ;
        RECT 99.250 193.290 99.540 193.335 ;
        RECT 95.580 193.150 99.540 193.290 ;
        RECT 95.580 193.105 95.870 193.150 ;
        RECT 97.680 193.105 97.970 193.150 ;
        RECT 99.250 193.105 99.540 193.150 ;
        RECT 108.460 193.290 108.750 193.335 ;
        RECT 110.560 193.290 110.850 193.335 ;
        RECT 112.130 193.290 112.420 193.335 ;
        RECT 108.460 193.150 112.420 193.290 ;
        RECT 108.460 193.105 108.750 193.150 ;
        RECT 110.560 193.105 110.850 193.150 ;
        RECT 112.130 193.105 112.420 193.150 ;
        RECT 77.615 192.810 81.600 192.950 ;
        RECT 73.015 192.765 73.305 192.810 ;
        RECT 77.615 192.765 77.905 192.810 ;
        RECT 81.280 192.750 81.600 192.810 ;
        RECT 95.095 192.765 95.385 192.995 ;
        RECT 95.975 192.950 96.265 192.995 ;
        RECT 97.165 192.950 97.455 192.995 ;
        RECT 99.685 192.950 99.975 192.995 ;
        RECT 95.975 192.810 99.975 192.950 ;
        RECT 95.975 192.765 96.265 192.810 ;
        RECT 97.165 192.765 97.455 192.810 ;
        RECT 99.685 192.765 99.975 192.810 ;
        RECT 103.360 192.950 103.680 193.010 ;
        RECT 105.215 192.950 105.505 192.995 ;
        RECT 107.500 192.950 107.820 193.010 ;
        RECT 103.360 192.810 107.820 192.950 ;
        RECT 103.360 192.750 103.680 192.810 ;
        RECT 105.215 192.765 105.505 192.810 ;
        RECT 107.500 192.750 107.820 192.810 ;
        RECT 107.960 192.750 108.280 193.010 ;
        RECT 108.855 192.950 109.145 192.995 ;
        RECT 110.045 192.950 110.335 192.995 ;
        RECT 112.565 192.950 112.855 192.995 ;
        RECT 108.855 192.810 112.855 192.950 ;
        RECT 108.855 192.765 109.145 192.810 ;
        RECT 110.045 192.765 110.335 192.810 ;
        RECT 112.565 192.765 112.855 192.810 ;
        RECT 120.840 192.750 121.160 193.010 ;
        RECT 127.280 192.750 127.600 193.010 ;
        RECT 131.970 192.950 132.110 193.430 ;
        RECT 132.340 192.950 132.660 193.010 ;
        RECT 131.970 192.810 136.710 192.950 ;
        RECT 132.340 192.750 132.660 192.810 ;
        RECT 60.595 192.610 60.885 192.655 ;
        RECT 60.120 192.470 60.885 192.610 ;
        RECT 60.120 192.410 60.440 192.470 ;
        RECT 60.595 192.425 60.885 192.470 ;
        RECT 61.515 192.610 61.805 192.655 ;
        RECT 61.960 192.610 62.280 192.670 ;
        RECT 61.515 192.470 62.280 192.610 ;
        RECT 61.515 192.425 61.805 192.470 ;
        RECT 61.960 192.410 62.280 192.470 ;
        RECT 69.780 192.610 70.100 192.670 ;
        RECT 71.160 192.610 71.480 192.670 ;
        RECT 73.475 192.610 73.765 192.655 ;
        RECT 69.780 192.470 73.765 192.610 ;
        RECT 69.780 192.410 70.100 192.470 ;
        RECT 71.160 192.410 71.480 192.470 ;
        RECT 73.475 192.425 73.765 192.470 ;
        RECT 94.160 192.610 94.480 192.670 ;
        RECT 95.540 192.610 95.860 192.670 ;
        RECT 94.160 192.470 95.860 192.610 ;
        RECT 94.160 192.410 94.480 192.470 ;
        RECT 95.540 192.410 95.860 192.470 ;
        RECT 118.540 192.610 118.860 192.670 ;
        RECT 122.235 192.610 122.525 192.655 ;
        RECT 118.540 192.470 122.525 192.610 ;
        RECT 118.540 192.410 118.860 192.470 ;
        RECT 122.235 192.425 122.525 192.470 ;
        RECT 130.960 192.410 131.280 192.670 ;
        RECT 133.720 192.610 134.040 192.670 ;
        RECT 136.570 192.655 136.710 192.810 ;
        RECT 134.655 192.610 134.945 192.655 ;
        RECT 133.720 192.470 134.945 192.610 ;
        RECT 133.720 192.410 134.040 192.470 ;
        RECT 134.655 192.425 134.945 192.470 ;
        RECT 136.495 192.425 136.785 192.655 ;
        RECT 57.910 192.130 59.890 192.270 ;
        RECT 80.820 192.270 81.140 192.330 ;
        RECT 81.295 192.270 81.585 192.315 ;
        RECT 86.800 192.270 87.120 192.330 ;
        RECT 80.820 192.130 87.120 192.270 ;
        RECT 54.600 192.070 54.920 192.130 ;
        RECT 57.375 192.085 57.665 192.130 ;
        RECT 80.820 192.070 81.140 192.130 ;
        RECT 81.295 192.085 81.585 192.130 ;
        RECT 86.800 192.070 87.120 192.130 ;
        RECT 96.430 192.270 96.720 192.315 ;
        RECT 104.295 192.270 104.585 192.315 ;
        RECT 108.420 192.270 108.740 192.330 ;
        RECT 109.200 192.270 109.490 192.315 ;
        RECT 96.430 192.130 102.670 192.270 ;
        RECT 96.430 192.085 96.720 192.130 ;
        RECT 44.940 191.790 51.150 191.930 ;
        RECT 54.140 191.930 54.460 191.990 ;
        RECT 59.200 191.930 59.520 191.990 ;
        RECT 59.675 191.930 59.965 191.975 ;
        RECT 54.140 191.790 59.965 191.930 ;
        RECT 44.940 191.730 45.260 191.790 ;
        RECT 54.140 191.730 54.460 191.790 ;
        RECT 59.200 191.730 59.520 191.790 ;
        RECT 59.675 191.745 59.965 191.790 ;
        RECT 61.500 191.930 61.820 191.990 ;
        RECT 66.100 191.930 66.420 191.990 ;
        RECT 61.500 191.790 66.420 191.930 ;
        RECT 61.500 191.730 61.820 191.790 ;
        RECT 66.100 191.730 66.420 191.790 ;
        RECT 90.940 191.930 91.260 191.990 ;
        RECT 102.530 191.975 102.670 192.130 ;
        RECT 104.295 192.130 108.190 192.270 ;
        RECT 104.295 192.085 104.585 192.130 ;
        RECT 91.415 191.930 91.705 191.975 ;
        RECT 90.940 191.790 91.705 191.930 ;
        RECT 90.940 191.730 91.260 191.790 ;
        RECT 91.415 191.745 91.705 191.790 ;
        RECT 102.455 191.745 102.745 191.975 ;
        RECT 104.755 191.930 105.045 191.975 ;
        RECT 106.580 191.930 106.900 191.990 ;
        RECT 104.755 191.790 106.900 191.930 ;
        RECT 108.050 191.930 108.190 192.130 ;
        RECT 108.420 192.130 109.490 192.270 ;
        RECT 108.420 192.070 108.740 192.130 ;
        RECT 109.200 192.085 109.490 192.130 ;
        RECT 130.515 192.270 130.805 192.315 ;
        RECT 135.115 192.270 135.405 192.315 ;
        RECT 130.515 192.130 135.405 192.270 ;
        RECT 130.515 192.085 130.805 192.130 ;
        RECT 135.115 192.085 135.405 192.130 ;
        RECT 135.575 192.085 135.865 192.315 ;
        RECT 116.240 191.930 116.560 191.990 ;
        RECT 108.050 191.790 116.560 191.930 ;
        RECT 104.755 191.745 105.045 191.790 ;
        RECT 106.580 191.730 106.900 191.790 ;
        RECT 116.240 191.730 116.560 191.790 ;
        RECT 119.920 191.730 120.240 191.990 ;
        RECT 120.395 191.930 120.685 191.975 ;
        RECT 127.740 191.930 128.060 191.990 ;
        RECT 120.395 191.790 128.060 191.930 ;
        RECT 120.395 191.745 120.685 191.790 ;
        RECT 127.740 191.730 128.060 191.790 ;
        RECT 130.040 191.930 130.360 191.990 ;
        RECT 135.650 191.930 135.790 192.085 ;
        RECT 130.040 191.790 135.790 191.930 ;
        RECT 130.040 191.730 130.360 191.790 ;
        RECT 17.270 191.110 146.990 191.590 ;
        RECT 35.280 190.910 35.600 190.970 ;
        RECT 36.200 190.910 36.520 190.970 ;
        RECT 35.280 190.770 36.520 190.910 ;
        RECT 35.280 190.710 35.600 190.770 ;
        RECT 36.200 190.710 36.520 190.770 ;
        RECT 44.020 190.910 44.340 190.970 ;
        RECT 65.180 190.910 65.500 190.970 ;
        RECT 44.020 190.770 65.500 190.910 ;
        RECT 44.020 190.710 44.340 190.770 ;
        RECT 65.180 190.710 65.500 190.770 ;
        RECT 66.115 190.910 66.405 190.955 ;
        RECT 71.620 190.910 71.940 190.970 ;
        RECT 66.115 190.770 71.940 190.910 ;
        RECT 66.115 190.725 66.405 190.770 ;
        RECT 71.620 190.710 71.940 190.770 ;
        RECT 72.080 190.955 72.400 190.970 ;
        RECT 72.080 190.910 72.515 190.955 ;
        RECT 73.460 190.910 73.780 190.970 ;
        RECT 81.740 190.910 82.060 190.970 ;
        RECT 72.080 190.770 73.780 190.910 ;
        RECT 72.080 190.725 72.515 190.770 ;
        RECT 72.080 190.710 72.400 190.725 ;
        RECT 73.460 190.710 73.780 190.770 ;
        RECT 80.910 190.770 82.060 190.910 ;
        RECT 35.740 190.570 36.060 190.630 ;
        RECT 38.515 190.570 38.805 190.615 ;
        RECT 41.720 190.570 42.040 190.630 ;
        RECT 35.740 190.430 37.350 190.570 ;
        RECT 35.740 190.370 36.060 190.430 ;
        RECT 24.715 190.045 25.005 190.275 ;
        RECT 25.620 190.230 25.940 190.290 ;
        RECT 35.280 190.230 35.600 190.290 ;
        RECT 37.210 190.275 37.350 190.430 ;
        RECT 38.515 190.430 39.190 190.570 ;
        RECT 38.515 190.385 38.805 190.430 ;
        RECT 39.050 190.275 39.190 190.430 ;
        RECT 40.430 190.430 42.040 190.570 ;
        RECT 36.215 190.230 36.505 190.275 ;
        RECT 25.620 190.090 35.600 190.230 ;
        RECT 24.790 189.890 24.930 190.045 ;
        RECT 25.620 190.030 25.940 190.090 ;
        RECT 35.280 190.030 35.600 190.090 ;
        RECT 35.830 190.090 36.505 190.230 ;
        RECT 35.830 189.950 35.970 190.090 ;
        RECT 36.215 190.045 36.505 190.090 ;
        RECT 36.675 190.045 36.965 190.275 ;
        RECT 37.135 190.045 37.425 190.275 ;
        RECT 38.975 190.045 39.265 190.275 ;
        RECT 26.080 189.890 26.400 189.950 ;
        RECT 24.790 189.750 26.400 189.890 ;
        RECT 26.080 189.690 26.400 189.750 ;
        RECT 35.740 189.690 36.060 189.950 ;
        RECT 36.750 189.890 36.890 190.045 ;
        RECT 39.880 190.030 40.200 190.290 ;
        RECT 40.430 190.275 40.570 190.430 ;
        RECT 41.720 190.370 42.040 190.430 ;
        RECT 56.915 190.570 57.205 190.615 ;
        RECT 59.675 190.570 59.965 190.615 ;
        RECT 60.120 190.570 60.440 190.630 ;
        RECT 63.800 190.570 64.120 190.630 ;
        RECT 64.275 190.570 64.565 190.615 ;
        RECT 56.915 190.430 60.440 190.570 ;
        RECT 56.915 190.385 57.205 190.430 ;
        RECT 59.675 190.385 59.965 190.430 ;
        RECT 60.120 190.370 60.440 190.430 ;
        RECT 61.130 190.430 63.110 190.570 ;
        RECT 40.355 190.045 40.645 190.275 ;
        RECT 40.815 190.230 41.105 190.275 ;
        RECT 41.260 190.230 41.580 190.290 ;
        RECT 42.640 190.230 42.960 190.290 ;
        RECT 40.815 190.090 42.960 190.230 ;
        RECT 40.815 190.045 41.105 190.090 ;
        RECT 41.260 190.030 41.580 190.090 ;
        RECT 42.640 190.030 42.960 190.090 ;
        RECT 43.575 190.230 43.865 190.275 ;
        RECT 47.700 190.230 48.020 190.290 ;
        RECT 43.575 190.090 48.020 190.230 ;
        RECT 43.575 190.045 43.865 190.090 ;
        RECT 47.700 190.030 48.020 190.090 ;
        RECT 50.935 190.230 51.225 190.275 ;
        RECT 52.760 190.230 53.080 190.290 ;
        RECT 50.935 190.090 53.080 190.230 ;
        RECT 50.935 190.045 51.225 190.090 ;
        RECT 52.760 190.030 53.080 190.090 ;
        RECT 54.155 190.230 54.445 190.275 ;
        RECT 55.520 190.230 55.840 190.290 ;
        RECT 54.155 190.090 55.840 190.230 ;
        RECT 54.155 190.045 54.445 190.090 ;
        RECT 39.420 189.890 39.740 189.950 ;
        RECT 36.750 189.750 39.740 189.890 ;
        RECT 39.420 189.690 39.740 189.750 ;
        RECT 47.255 189.890 47.545 189.935 ;
        RECT 54.230 189.890 54.370 190.045 ;
        RECT 55.520 190.030 55.840 190.090 ;
        RECT 56.455 190.230 56.745 190.275 ;
        RECT 57.360 190.230 57.680 190.290 ;
        RECT 56.455 190.090 57.680 190.230 ;
        RECT 56.455 190.045 56.745 190.090 ;
        RECT 57.360 190.030 57.680 190.090 ;
        RECT 58.755 190.045 59.045 190.275 ;
        RECT 47.255 189.750 54.370 189.890 ;
        RECT 47.255 189.705 47.545 189.750 ;
        RECT 34.820 189.550 35.140 189.610 ;
        RECT 36.660 189.550 36.980 189.610 ;
        RECT 34.820 189.410 36.980 189.550 ;
        RECT 34.820 189.350 35.140 189.410 ;
        RECT 36.660 189.350 36.980 189.410 ;
        RECT 46.320 189.550 46.640 189.610 ;
        RECT 58.830 189.550 58.970 190.045 ;
        RECT 60.580 190.030 60.900 190.290 ;
        RECT 59.660 189.890 59.980 189.950 ;
        RECT 61.130 189.935 61.270 190.430 ;
        RECT 61.960 190.030 62.280 190.290 ;
        RECT 61.055 189.890 61.345 189.935 ;
        RECT 59.660 189.750 61.345 189.890 ;
        RECT 59.660 189.690 59.980 189.750 ;
        RECT 61.055 189.705 61.345 189.750 ;
        RECT 62.050 189.550 62.190 190.030 ;
        RECT 46.320 189.410 62.190 189.550 ;
        RECT 62.970 189.550 63.110 190.430 ;
        RECT 63.800 190.430 64.565 190.570 ;
        RECT 63.800 190.370 64.120 190.430 ;
        RECT 64.275 190.385 64.565 190.430 ;
        RECT 64.735 190.570 65.025 190.615 ;
        RECT 65.640 190.570 65.960 190.630 ;
        RECT 67.495 190.570 67.785 190.615 ;
        RECT 64.735 190.430 67.785 190.570 ;
        RECT 64.735 190.385 65.025 190.430 ;
        RECT 65.640 190.370 65.960 190.430 ;
        RECT 67.495 190.385 67.785 190.430 ;
        RECT 69.795 190.570 70.085 190.615 ;
        RECT 71.175 190.570 71.465 190.615 ;
        RECT 69.795 190.430 70.470 190.570 ;
        RECT 69.795 190.385 70.085 190.430 ;
        RECT 70.330 190.290 70.470 190.430 ;
        RECT 71.175 190.430 74.150 190.570 ;
        RECT 71.175 190.385 71.465 190.430 ;
        RECT 63.340 190.030 63.660 190.290 ;
        RECT 65.180 190.030 65.500 190.290 ;
        RECT 66.560 190.030 66.880 190.290 ;
        RECT 69.335 190.220 69.625 190.275 ;
        RECT 69.335 190.080 70.010 190.220 ;
        RECT 69.335 190.045 69.625 190.080 ;
        RECT 66.100 189.890 66.420 189.950 ;
        RECT 68.415 189.890 68.705 189.935 ;
        RECT 66.100 189.750 68.705 189.890 ;
        RECT 69.870 189.890 70.010 190.080 ;
        RECT 70.240 190.030 70.560 190.290 ;
        RECT 70.715 190.230 71.005 190.275 ;
        RECT 73.475 190.230 73.765 190.275 ;
        RECT 70.715 190.090 73.765 190.230 ;
        RECT 70.715 190.045 71.005 190.090 ;
        RECT 73.475 190.045 73.765 190.090 ;
        RECT 74.010 189.950 74.150 190.430 ;
        RECT 80.910 190.275 81.050 190.770 ;
        RECT 81.740 190.710 82.060 190.770 ;
        RECT 90.940 190.710 91.260 190.970 ;
        RECT 94.620 190.910 94.940 190.970 ;
        RECT 95.555 190.910 95.845 190.955 ;
        RECT 94.620 190.770 95.845 190.910 ;
        RECT 94.620 190.710 94.940 190.770 ;
        RECT 95.555 190.725 95.845 190.770 ;
        RECT 106.580 190.710 106.900 190.970 ;
        RECT 108.420 190.710 108.740 190.970 ;
        RECT 110.275 190.910 110.565 190.955 ;
        RECT 111.640 190.910 111.960 190.970 ;
        RECT 110.275 190.770 111.960 190.910 ;
        RECT 110.275 190.725 110.565 190.770 ;
        RECT 111.640 190.710 111.960 190.770 ;
        RECT 116.240 190.710 116.560 190.970 ;
        RECT 118.540 190.710 118.860 190.970 ;
        RECT 127.740 190.710 128.060 190.970 ;
        RECT 133.720 190.710 134.040 190.970 ;
        RECT 134.180 190.710 134.500 190.970 ;
        RECT 81.295 190.570 81.585 190.615 ;
        RECT 82.200 190.570 82.520 190.630 ;
        RECT 81.295 190.430 82.520 190.570 ;
        RECT 81.295 190.385 81.585 190.430 ;
        RECT 82.200 190.370 82.520 190.430 ;
        RECT 107.960 190.570 108.280 190.630 ;
        RECT 123.600 190.570 123.920 190.630 ;
        RECT 107.960 190.430 123.920 190.570 ;
        RECT 107.960 190.370 108.280 190.430 ;
        RECT 79.915 190.045 80.205 190.275 ;
        RECT 80.835 190.045 81.125 190.275 ;
        RECT 81.755 190.045 82.045 190.275 ;
        RECT 90.495 190.230 90.785 190.275 ;
        RECT 96.460 190.230 96.780 190.290 ;
        RECT 90.495 190.090 96.780 190.230 ;
        RECT 90.495 190.045 90.785 190.090 ;
        RECT 72.080 189.890 72.400 189.950 ;
        RECT 73.920 189.890 74.240 189.950 ;
        RECT 76.235 189.890 76.525 189.935 ;
        RECT 69.870 189.750 72.400 189.890 ;
        RECT 66.100 189.690 66.420 189.750 ;
        RECT 68.415 189.705 68.705 189.750 ;
        RECT 72.080 189.690 72.400 189.750 ;
        RECT 73.090 189.750 76.525 189.890 ;
        RECT 79.990 189.890 80.130 190.045 ;
        RECT 81.280 189.890 81.600 189.950 ;
        RECT 79.990 189.750 81.600 189.890 ;
        RECT 73.090 189.550 73.230 189.750 ;
        RECT 73.920 189.690 74.240 189.750 ;
        RECT 76.235 189.705 76.525 189.750 ;
        RECT 81.280 189.690 81.600 189.750 ;
        RECT 62.970 189.410 73.230 189.550 ;
        RECT 73.460 189.550 73.780 189.610 ;
        RECT 81.830 189.550 81.970 190.045 ;
        RECT 96.460 190.030 96.780 190.090 ;
        RECT 96.920 190.230 97.240 190.290 ;
        RECT 97.395 190.230 97.685 190.275 ;
        RECT 99.695 190.230 99.985 190.275 ;
        RECT 96.920 190.090 97.685 190.230 ;
        RECT 96.920 190.030 97.240 190.090 ;
        RECT 97.395 190.045 97.685 190.090 ;
        RECT 97.930 190.090 99.985 190.230 ;
        RECT 97.930 189.950 98.070 190.090 ;
        RECT 99.695 190.045 99.985 190.090 ;
        RECT 101.980 190.230 102.300 190.290 ;
        RECT 103.375 190.230 103.665 190.275 ;
        RECT 101.980 190.090 103.665 190.230 ;
        RECT 101.980 190.030 102.300 190.090 ;
        RECT 103.375 190.045 103.665 190.090 ;
        RECT 110.735 190.230 111.025 190.275 ;
        RECT 112.575 190.230 112.865 190.275 ;
        RECT 110.735 190.090 112.865 190.230 ;
        RECT 110.735 190.045 111.025 190.090 ;
        RECT 112.575 190.045 112.865 190.090 ;
        RECT 114.860 190.230 115.180 190.290 ;
        RECT 115.335 190.230 115.625 190.275 ;
        RECT 114.860 190.090 115.625 190.230 ;
        RECT 114.860 190.030 115.180 190.090 ;
        RECT 115.335 190.045 115.625 190.090 ;
        RECT 117.160 190.230 117.480 190.290 ;
        RECT 120.930 190.275 121.070 190.430 ;
        RECT 123.600 190.370 123.920 190.430 ;
        RECT 118.095 190.230 118.385 190.275 ;
        RECT 117.160 190.090 118.385 190.230 ;
        RECT 117.160 190.030 117.480 190.090 ;
        RECT 118.095 190.045 118.385 190.090 ;
        RECT 120.855 190.045 121.145 190.275 ;
        RECT 122.190 190.230 122.480 190.275 ;
        RECT 124.060 190.230 124.380 190.290 ;
        RECT 122.190 190.090 124.380 190.230 ;
        RECT 127.830 190.230 127.970 190.710 ;
        RECT 128.660 190.570 128.980 190.630 ;
        RECT 132.815 190.570 133.105 190.615 ;
        RECT 128.660 190.430 133.105 190.570 ;
        RECT 128.660 190.370 128.980 190.430 ;
        RECT 132.815 190.385 133.105 190.430 ;
        RECT 130.975 190.230 131.265 190.275 ;
        RECT 127.830 190.090 131.265 190.230 ;
        RECT 122.190 190.045 122.480 190.090 ;
        RECT 124.060 190.030 124.380 190.090 ;
        RECT 130.975 190.045 131.265 190.090 ;
        RECT 131.880 190.030 132.200 190.290 ;
        RECT 139.815 190.230 140.105 190.275 ;
        RECT 140.620 190.230 140.940 190.290 ;
        RECT 139.815 190.090 140.940 190.230 ;
        RECT 139.815 190.045 140.105 190.090 ;
        RECT 140.620 190.030 140.940 190.090 ;
        RECT 91.875 189.705 92.165 189.935 ;
        RECT 73.460 189.410 81.970 189.550 ;
        RECT 91.950 189.550 92.090 189.705 ;
        RECT 97.840 189.690 98.160 189.950 ;
        RECT 98.775 189.890 99.065 189.935 ;
        RECT 100.140 189.890 100.460 189.950 ;
        RECT 98.775 189.750 100.460 189.890 ;
        RECT 98.775 189.705 99.065 189.750 ;
        RECT 100.140 189.690 100.460 189.750 ;
        RECT 107.500 189.890 107.820 189.950 ;
        RECT 111.195 189.890 111.485 189.935 ;
        RECT 107.500 189.750 111.485 189.890 ;
        RECT 107.500 189.690 107.820 189.750 ;
        RECT 111.195 189.705 111.485 189.750 ;
        RECT 119.475 189.705 119.765 189.935 ;
        RECT 121.735 189.890 122.025 189.935 ;
        RECT 122.925 189.890 123.215 189.935 ;
        RECT 125.445 189.890 125.735 189.935 ;
        RECT 121.735 189.750 125.735 189.890 ;
        RECT 121.735 189.705 122.025 189.750 ;
        RECT 122.925 189.705 123.215 189.750 ;
        RECT 125.445 189.705 125.735 189.750 ;
        RECT 136.505 189.890 136.795 189.935 ;
        RECT 139.025 189.890 139.315 189.935 ;
        RECT 140.215 189.890 140.505 189.935 ;
        RECT 136.505 189.750 140.505 189.890 ;
        RECT 136.505 189.705 136.795 189.750 ;
        RECT 139.025 189.705 139.315 189.750 ;
        RECT 140.215 189.705 140.505 189.750 ;
        RECT 141.095 189.705 141.385 189.935 ;
        RECT 103.360 189.550 103.680 189.610 ;
        RECT 91.950 189.410 103.680 189.550 ;
        RECT 46.320 189.350 46.640 189.410 ;
        RECT 73.460 189.350 73.780 189.410 ;
        RECT 103.360 189.350 103.680 189.410 ;
        RECT 116.240 189.550 116.560 189.610 ;
        RECT 119.550 189.550 119.690 189.705 ;
        RECT 120.840 189.550 121.160 189.610 ;
        RECT 116.240 189.410 121.160 189.550 ;
        RECT 116.240 189.350 116.560 189.410 ;
        RECT 120.840 189.350 121.160 189.410 ;
        RECT 121.340 189.550 121.630 189.595 ;
        RECT 123.440 189.550 123.730 189.595 ;
        RECT 125.010 189.550 125.300 189.595 ;
        RECT 121.340 189.410 125.300 189.550 ;
        RECT 121.340 189.365 121.630 189.410 ;
        RECT 123.440 189.365 123.730 189.410 ;
        RECT 125.010 189.365 125.300 189.410 ;
        RECT 136.940 189.550 137.230 189.595 ;
        RECT 138.510 189.550 138.800 189.595 ;
        RECT 140.610 189.550 140.900 189.595 ;
        RECT 136.940 189.410 140.900 189.550 ;
        RECT 136.940 189.365 137.230 189.410 ;
        RECT 138.510 189.365 138.800 189.410 ;
        RECT 140.610 189.365 140.900 189.410 ;
        RECT 25.175 189.210 25.465 189.255 ;
        RECT 29.300 189.210 29.620 189.270 ;
        RECT 25.175 189.070 29.620 189.210 ;
        RECT 25.175 189.025 25.465 189.070 ;
        RECT 29.300 189.010 29.620 189.070 ;
        RECT 39.420 189.210 39.740 189.270 ;
        RECT 42.195 189.210 42.485 189.255 ;
        RECT 39.420 189.070 42.485 189.210 ;
        RECT 39.420 189.010 39.740 189.070 ;
        RECT 42.195 189.025 42.485 189.070 ;
        RECT 58.280 189.010 58.600 189.270 ;
        RECT 60.120 189.210 60.440 189.270 ;
        RECT 60.595 189.210 60.885 189.255 ;
        RECT 60.120 189.070 60.885 189.210 ;
        RECT 60.120 189.010 60.440 189.070 ;
        RECT 60.595 189.025 60.885 189.070 ;
        RECT 62.420 189.210 62.740 189.270 ;
        RECT 62.895 189.210 63.185 189.255 ;
        RECT 62.420 189.070 63.185 189.210 ;
        RECT 62.420 189.010 62.740 189.070 ;
        RECT 62.895 189.025 63.185 189.070 ;
        RECT 70.700 189.010 71.020 189.270 ;
        RECT 71.160 189.210 71.480 189.270 ;
        RECT 72.095 189.210 72.385 189.255 ;
        RECT 71.160 189.070 72.385 189.210 ;
        RECT 71.160 189.010 71.480 189.070 ;
        RECT 72.095 189.025 72.385 189.070 ;
        RECT 72.540 189.210 72.860 189.270 ;
        RECT 73.015 189.210 73.305 189.255 ;
        RECT 72.540 189.070 73.305 189.210 ;
        RECT 72.540 189.010 72.860 189.070 ;
        RECT 73.015 189.025 73.305 189.070 ;
        RECT 85.880 189.210 86.200 189.270 ;
        RECT 88.655 189.210 88.945 189.255 ;
        RECT 85.880 189.070 88.945 189.210 ;
        RECT 85.880 189.010 86.200 189.070 ;
        RECT 88.655 189.025 88.945 189.070 ;
        RECT 102.440 189.210 102.760 189.270 ;
        RECT 102.915 189.210 103.205 189.255 ;
        RECT 102.440 189.070 103.205 189.210 ;
        RECT 102.440 189.010 102.760 189.070 ;
        RECT 102.915 189.025 103.205 189.070 ;
        RECT 128.200 189.010 128.520 189.270 ;
        RECT 137.400 189.210 137.720 189.270 ;
        RECT 141.170 189.210 141.310 189.705 ;
        RECT 137.400 189.070 141.310 189.210 ;
        RECT 137.400 189.010 137.720 189.070 ;
        RECT 17.270 188.390 146.990 188.870 ;
        RECT 23.335 188.190 23.625 188.235 ;
        RECT 32.060 188.190 32.380 188.250 ;
        RECT 23.335 188.050 32.380 188.190 ;
        RECT 23.335 188.005 23.625 188.050 ;
        RECT 32.060 187.990 32.380 188.050 ;
        RECT 41.735 188.190 42.025 188.235 ;
        RECT 42.180 188.190 42.500 188.250 ;
        RECT 80.820 188.190 81.140 188.250 ;
        RECT 41.735 188.050 42.500 188.190 ;
        RECT 41.735 188.005 42.025 188.050 ;
        RECT 42.180 187.990 42.500 188.050 ;
        RECT 55.150 188.050 81.140 188.190 ;
        RECT 24.700 187.850 25.020 187.910 ;
        RECT 27.920 187.850 28.240 187.910 ;
        RECT 31.140 187.850 31.460 187.910 ;
        RECT 54.140 187.850 54.460 187.910 ;
        RECT 24.700 187.710 31.460 187.850 ;
        RECT 24.700 187.650 25.020 187.710 ;
        RECT 27.920 187.650 28.240 187.710 ;
        RECT 31.140 187.650 31.460 187.710 ;
        RECT 43.190 187.710 54.460 187.850 ;
        RECT 24.790 187.510 24.930 187.650 ;
        RECT 24.330 187.370 24.930 187.510 ;
        RECT 26.555 187.510 26.845 187.555 ;
        RECT 30.220 187.510 30.540 187.570 ;
        RECT 43.190 187.510 43.330 187.710 ;
        RECT 54.140 187.650 54.460 187.710 ;
        RECT 26.555 187.370 30.540 187.510 ;
        RECT 24.330 186.875 24.470 187.370 ;
        RECT 26.555 187.325 26.845 187.370 ;
        RECT 30.220 187.310 30.540 187.370 ;
        RECT 36.290 187.370 43.330 187.510 ;
        RECT 43.560 187.510 43.880 187.570 ;
        RECT 44.035 187.510 44.325 187.555 ;
        RECT 52.760 187.510 53.080 187.570 ;
        RECT 43.560 187.370 53.080 187.510 ;
        RECT 24.715 187.170 25.005 187.215 ;
        RECT 26.080 187.170 26.400 187.230 ;
        RECT 24.715 187.030 26.400 187.170 ;
        RECT 24.715 186.985 25.005 187.030 ;
        RECT 26.080 186.970 26.400 187.030 ;
        RECT 27.000 186.970 27.320 187.230 ;
        RECT 27.475 187.170 27.765 187.215 ;
        RECT 28.395 187.170 28.685 187.215 ;
        RECT 27.475 187.030 28.685 187.170 ;
        RECT 27.475 186.985 27.765 187.030 ;
        RECT 28.395 186.985 28.685 187.030 ;
        RECT 24.255 186.645 24.545 186.875 ;
        RECT 25.620 186.630 25.940 186.890 ;
        RECT 28.470 186.830 28.610 186.985 ;
        RECT 29.300 186.970 29.620 187.230 ;
        RECT 34.835 187.170 35.125 187.215 ;
        RECT 35.280 187.170 35.600 187.230 ;
        RECT 34.835 187.030 35.600 187.170 ;
        RECT 34.835 186.985 35.125 187.030 ;
        RECT 35.280 186.970 35.600 187.030 ;
        RECT 35.740 186.970 36.060 187.230 ;
        RECT 36.290 187.215 36.430 187.370 ;
        RECT 43.560 187.310 43.880 187.370 ;
        RECT 44.035 187.325 44.325 187.370 ;
        RECT 52.760 187.310 53.080 187.370 ;
        RECT 36.215 186.985 36.505 187.215 ;
        RECT 36.660 186.970 36.980 187.230 ;
        RECT 37.580 187.170 37.900 187.230 ;
        RECT 38.500 187.170 38.820 187.230 ;
        RECT 37.580 187.030 38.820 187.170 ;
        RECT 37.580 186.970 37.900 187.030 ;
        RECT 38.500 186.970 38.820 187.030 ;
        RECT 39.435 186.985 39.725 187.215 ;
        RECT 35.830 186.830 35.970 186.970 ;
        RECT 38.975 186.830 39.265 186.875 ;
        RECT 28.470 186.690 35.510 186.830 ;
        RECT 35.830 186.690 39.265 186.830 ;
        RECT 39.510 186.830 39.650 186.985 ;
        RECT 39.880 186.970 40.200 187.230 ;
        RECT 41.735 187.170 42.025 187.215 ;
        RECT 44.480 187.170 44.800 187.230 ;
        RECT 41.735 187.030 44.800 187.170 ;
        RECT 41.735 186.985 42.025 187.030 ;
        RECT 44.480 186.970 44.800 187.030 ;
        RECT 47.700 187.170 48.020 187.230 ;
        RECT 55.150 187.170 55.290 188.050 ;
        RECT 80.820 187.990 81.140 188.050 ;
        RECT 92.795 188.190 93.085 188.235 ;
        RECT 97.840 188.190 98.160 188.250 ;
        RECT 92.795 188.050 98.160 188.190 ;
        RECT 92.795 188.005 93.085 188.050 ;
        RECT 97.840 187.990 98.160 188.050 ;
        RECT 116.715 188.190 117.005 188.235 ;
        RECT 118.540 188.190 118.860 188.250 ;
        RECT 116.715 188.050 118.860 188.190 ;
        RECT 116.715 188.005 117.005 188.050 ;
        RECT 118.540 187.990 118.860 188.050 ;
        RECT 124.060 187.990 124.380 188.250 ;
        RECT 126.820 188.190 127.140 188.250 ;
        RECT 127.295 188.190 127.585 188.235 ;
        RECT 126.820 188.050 127.585 188.190 ;
        RECT 126.820 187.990 127.140 188.050 ;
        RECT 127.295 188.005 127.585 188.050 ;
        RECT 129.135 188.190 129.425 188.235 ;
        RECT 132.800 188.190 133.120 188.250 ;
        RECT 129.135 188.050 133.120 188.190 ;
        RECT 129.135 188.005 129.425 188.050 ;
        RECT 57.820 187.650 58.140 187.910 ;
        RECT 62.880 187.650 63.200 187.910 ;
        RECT 63.340 187.850 63.660 187.910 ;
        RECT 64.735 187.850 65.025 187.895 ;
        RECT 63.340 187.710 65.025 187.850 ;
        RECT 63.340 187.650 63.660 187.710 ;
        RECT 64.735 187.665 65.025 187.710 ;
        RECT 72.095 187.850 72.385 187.895 ;
        RECT 76.680 187.850 76.970 187.895 ;
        RECT 78.250 187.850 78.540 187.895 ;
        RECT 80.350 187.850 80.640 187.895 ;
        RECT 72.095 187.710 75.990 187.850 ;
        RECT 72.095 187.665 72.385 187.710 ;
        RECT 58.295 187.510 58.585 187.555 ;
        RECT 61.055 187.510 61.345 187.555 ;
        RECT 56.990 187.370 58.050 187.510 ;
        RECT 56.990 187.215 57.130 187.370 ;
        RECT 47.700 187.030 55.290 187.170 ;
        RECT 47.700 186.970 48.020 187.030 ;
        RECT 56.915 186.985 57.205 187.215 ;
        RECT 57.375 186.985 57.665 187.215 ;
        RECT 57.910 187.170 58.050 187.370 ;
        RECT 58.295 187.370 61.345 187.510 ;
        RECT 62.970 187.510 63.110 187.650 ;
        RECT 66.560 187.510 66.880 187.570 ;
        RECT 62.970 187.370 66.880 187.510 ;
        RECT 58.295 187.325 58.585 187.370 ;
        RECT 61.055 187.325 61.345 187.370 ;
        RECT 66.560 187.310 66.880 187.370 ;
        RECT 72.540 187.310 72.860 187.570 ;
        RECT 59.660 187.170 59.980 187.230 ;
        RECT 57.910 187.030 59.980 187.170 ;
        RECT 40.340 186.830 40.660 186.890 ;
        RECT 39.510 186.690 40.660 186.830 ;
        RECT 22.400 186.290 22.720 186.550 ;
        RECT 23.255 186.490 23.545 186.535 ;
        RECT 28.395 186.490 28.685 186.535 ;
        RECT 23.255 186.350 28.685 186.490 ;
        RECT 35.370 186.490 35.510 186.690 ;
        RECT 38.975 186.645 39.265 186.690 ;
        RECT 40.340 186.630 40.660 186.690 ;
        RECT 53.220 186.830 53.540 186.890 ;
        RECT 57.450 186.830 57.590 186.985 ;
        RECT 59.660 186.970 59.980 187.030 ;
        RECT 60.120 186.970 60.440 187.230 ;
        RECT 60.580 186.970 60.900 187.230 ;
        RECT 61.500 186.970 61.820 187.230 ;
        RECT 62.420 186.970 62.740 187.230 ;
        RECT 63.355 186.985 63.645 187.215 ;
        RECT 58.280 186.830 58.600 186.890 ;
        RECT 58.755 186.830 59.045 186.875 ;
        RECT 53.220 186.690 59.045 186.830 ;
        RECT 63.430 186.830 63.570 186.985 ;
        RECT 63.800 186.970 64.120 187.230 ;
        RECT 70.700 187.170 71.020 187.230 ;
        RECT 72.095 187.170 72.385 187.215 ;
        RECT 70.700 187.030 72.385 187.170 ;
        RECT 75.850 187.170 75.990 187.710 ;
        RECT 76.680 187.710 80.640 187.850 ;
        RECT 76.680 187.665 76.970 187.710 ;
        RECT 78.250 187.665 78.540 187.710 ;
        RECT 80.350 187.665 80.640 187.710 ;
        RECT 85.000 187.850 85.290 187.895 ;
        RECT 87.100 187.850 87.390 187.895 ;
        RECT 88.670 187.850 88.960 187.895 ;
        RECT 85.000 187.710 88.960 187.850 ;
        RECT 85.000 187.665 85.290 187.710 ;
        RECT 87.100 187.665 87.390 187.710 ;
        RECT 88.670 187.665 88.960 187.710 ;
        RECT 91.415 187.850 91.705 187.895 ;
        RECT 94.620 187.850 94.940 187.910 ;
        RECT 91.415 187.710 94.940 187.850 ;
        RECT 91.415 187.665 91.705 187.710 ;
        RECT 94.620 187.650 94.940 187.710 ;
        RECT 95.540 187.850 95.830 187.895 ;
        RECT 97.110 187.850 97.400 187.895 ;
        RECT 99.210 187.850 99.500 187.895 ;
        RECT 95.540 187.710 99.500 187.850 ;
        RECT 95.540 187.665 95.830 187.710 ;
        RECT 97.110 187.665 97.400 187.710 ;
        RECT 99.210 187.665 99.500 187.710 ;
        RECT 119.460 187.850 119.750 187.895 ;
        RECT 121.030 187.850 121.320 187.895 ;
        RECT 123.130 187.850 123.420 187.895 ;
        RECT 119.460 187.710 123.420 187.850 ;
        RECT 119.460 187.665 119.750 187.710 ;
        RECT 121.030 187.665 121.320 187.710 ;
        RECT 123.130 187.665 123.420 187.710 ;
        RECT 126.360 187.850 126.680 187.910 ;
        RECT 129.210 187.850 129.350 188.005 ;
        RECT 132.800 187.990 133.120 188.050 ;
        RECT 140.620 188.190 140.940 188.250 ;
        RECT 141.095 188.190 141.385 188.235 ;
        RECT 140.620 188.050 141.385 188.190 ;
        RECT 140.620 187.990 140.940 188.050 ;
        RECT 141.095 188.005 141.385 188.050 ;
        RECT 126.360 187.710 129.350 187.850 ;
        RECT 129.580 187.850 129.900 187.910 ;
        RECT 131.420 187.850 131.740 187.910 ;
        RECT 129.580 187.710 131.740 187.850 ;
        RECT 126.360 187.650 126.680 187.710 ;
        RECT 129.580 187.650 129.900 187.710 ;
        RECT 131.420 187.650 131.740 187.710 ;
        RECT 134.220 187.850 134.510 187.895 ;
        RECT 136.320 187.850 136.610 187.895 ;
        RECT 137.890 187.850 138.180 187.895 ;
        RECT 134.220 187.710 138.180 187.850 ;
        RECT 134.220 187.665 134.510 187.710 ;
        RECT 136.320 187.665 136.610 187.710 ;
        RECT 137.890 187.665 138.180 187.710 ;
        RECT 76.245 187.510 76.535 187.555 ;
        RECT 78.765 187.510 79.055 187.555 ;
        RECT 79.955 187.510 80.245 187.555 ;
        RECT 76.245 187.370 80.245 187.510 ;
        RECT 76.245 187.325 76.535 187.370 ;
        RECT 78.765 187.325 79.055 187.370 ;
        RECT 79.955 187.325 80.245 187.370 ;
        RECT 85.395 187.510 85.685 187.555 ;
        RECT 86.585 187.510 86.875 187.555 ;
        RECT 89.105 187.510 89.395 187.555 ;
        RECT 85.395 187.370 89.395 187.510 ;
        RECT 85.395 187.325 85.685 187.370 ;
        RECT 86.585 187.325 86.875 187.370 ;
        RECT 89.105 187.325 89.395 187.370 ;
        RECT 95.105 187.510 95.395 187.555 ;
        RECT 97.625 187.510 97.915 187.555 ;
        RECT 98.815 187.510 99.105 187.555 ;
        RECT 95.105 187.370 99.105 187.510 ;
        RECT 95.105 187.325 95.395 187.370 ;
        RECT 97.625 187.325 97.915 187.370 ;
        RECT 98.815 187.325 99.105 187.370 ;
        RECT 99.680 187.310 100.000 187.570 ;
        RECT 102.440 187.310 102.760 187.570 ;
        RECT 102.915 187.510 103.205 187.555 ;
        RECT 103.360 187.510 103.680 187.570 ;
        RECT 102.915 187.370 103.680 187.510 ;
        RECT 102.915 187.325 103.205 187.370 ;
        RECT 79.500 187.170 79.790 187.215 ;
        RECT 75.850 187.030 79.790 187.170 ;
        RECT 70.700 186.970 71.020 187.030 ;
        RECT 72.095 186.985 72.385 187.030 ;
        RECT 79.500 186.985 79.790 187.030 ;
        RECT 80.835 187.170 81.125 187.215 ;
        RECT 81.280 187.170 81.600 187.230 ;
        RECT 84.515 187.170 84.805 187.215 ;
        RECT 101.060 187.170 101.380 187.230 ;
        RECT 102.990 187.170 103.130 187.325 ;
        RECT 103.360 187.310 103.680 187.370 ;
        RECT 119.025 187.510 119.315 187.555 ;
        RECT 121.545 187.510 121.835 187.555 ;
        RECT 122.735 187.510 123.025 187.555 ;
        RECT 119.025 187.370 123.025 187.510 ;
        RECT 119.025 187.325 119.315 187.370 ;
        RECT 121.545 187.325 121.835 187.370 ;
        RECT 122.735 187.325 123.025 187.370 ;
        RECT 123.600 187.510 123.920 187.570 ;
        RECT 127.280 187.510 127.600 187.570 ;
        RECT 133.735 187.510 134.025 187.555 ;
        RECT 123.600 187.370 134.025 187.510 ;
        RECT 123.600 187.310 123.920 187.370 ;
        RECT 127.280 187.310 127.600 187.370 ;
        RECT 133.735 187.325 134.025 187.370 ;
        RECT 134.615 187.510 134.905 187.555 ;
        RECT 135.805 187.510 136.095 187.555 ;
        RECT 138.325 187.510 138.615 187.555 ;
        RECT 134.615 187.370 138.615 187.510 ;
        RECT 134.615 187.325 134.905 187.370 ;
        RECT 135.805 187.325 136.095 187.370 ;
        RECT 138.325 187.325 138.615 187.370 ;
        RECT 138.870 187.370 143.150 187.510 ;
        RECT 80.835 187.030 86.570 187.170 ;
        RECT 80.835 186.985 81.125 187.030 ;
        RECT 81.280 186.970 81.600 187.030 ;
        RECT 84.515 186.985 84.805 187.030 ;
        RECT 86.430 186.890 86.570 187.030 ;
        RECT 101.060 187.030 103.130 187.170 ;
        RECT 108.895 187.170 109.185 187.215 ;
        RECT 110.260 187.170 110.580 187.230 ;
        RECT 108.895 187.030 110.580 187.170 ;
        RECT 101.060 186.970 101.380 187.030 ;
        RECT 108.895 186.985 109.185 187.030 ;
        RECT 110.260 186.970 110.580 187.030 ;
        RECT 110.720 186.970 111.040 187.230 ;
        RECT 122.220 187.215 122.540 187.230 ;
        RECT 122.220 186.985 122.570 187.215 ;
        RECT 124.995 187.170 125.285 187.215 ;
        RECT 126.835 187.170 127.125 187.215 ;
        RECT 128.200 187.170 128.520 187.230 ;
        RECT 124.995 187.030 126.590 187.170 ;
        RECT 124.995 186.985 125.285 187.030 ;
        RECT 122.220 186.970 122.540 186.985 ;
        RECT 66.560 186.830 66.880 186.890 ;
        RECT 63.430 186.690 66.880 186.830 ;
        RECT 53.220 186.630 53.540 186.690 ;
        RECT 58.280 186.630 58.600 186.690 ;
        RECT 58.755 186.645 59.045 186.690 ;
        RECT 66.560 186.630 66.880 186.690 ;
        RECT 73.460 186.630 73.780 186.890 ;
        RECT 85.880 186.875 86.200 186.890 ;
        RECT 85.850 186.830 86.200 186.875 ;
        RECT 85.685 186.690 86.200 186.830 ;
        RECT 85.850 186.645 86.200 186.690 ;
        RECT 85.880 186.630 86.200 186.645 ;
        RECT 86.340 186.630 86.660 186.890 ;
        RECT 98.470 186.830 98.760 186.875 ;
        RECT 98.470 186.690 100.370 186.830 ;
        RECT 98.470 186.645 98.760 186.690 ;
        RECT 37.580 186.490 37.900 186.550 ;
        RECT 35.370 186.350 37.900 186.490 ;
        RECT 23.255 186.305 23.545 186.350 ;
        RECT 28.395 186.305 28.685 186.350 ;
        RECT 37.580 186.290 37.900 186.350 ;
        RECT 38.040 186.290 38.360 186.550 ;
        RECT 42.655 186.490 42.945 186.535 ;
        RECT 45.400 186.490 45.720 186.550 ;
        RECT 42.655 186.350 45.720 186.490 ;
        RECT 42.655 186.305 42.945 186.350 ;
        RECT 45.400 186.290 45.720 186.350 ;
        RECT 73.920 186.290 74.240 186.550 ;
        RECT 100.230 186.535 100.370 186.690 ;
        RECT 109.355 186.645 109.645 186.875 ;
        RECT 109.815 186.830 110.105 186.875 ;
        RECT 115.780 186.830 116.100 186.890 ;
        RECT 125.440 186.830 125.760 186.890 ;
        RECT 109.815 186.690 116.100 186.830 ;
        RECT 109.815 186.645 110.105 186.690 ;
        RECT 100.155 186.305 100.445 186.535 ;
        RECT 101.995 186.490 102.285 186.535 ;
        RECT 107.500 186.490 107.820 186.550 ;
        RECT 101.995 186.350 107.820 186.490 ;
        RECT 101.995 186.305 102.285 186.350 ;
        RECT 107.500 186.290 107.820 186.350 ;
        RECT 107.975 186.490 108.265 186.535 ;
        RECT 108.420 186.490 108.740 186.550 ;
        RECT 107.975 186.350 108.740 186.490 ;
        RECT 109.430 186.490 109.570 186.645 ;
        RECT 115.780 186.630 116.100 186.690 ;
        RECT 122.080 186.690 125.760 186.830 ;
        RECT 112.100 186.490 112.420 186.550 ;
        RECT 122.080 186.490 122.220 186.690 ;
        RECT 125.440 186.630 125.760 186.690 ;
        RECT 125.900 186.630 126.220 186.890 ;
        RECT 126.450 186.830 126.590 187.030 ;
        RECT 126.835 187.030 128.520 187.170 ;
        RECT 126.835 186.985 127.125 187.030 ;
        RECT 128.200 186.970 128.520 187.030 ;
        RECT 128.675 186.985 128.965 187.215 ;
        RECT 127.740 186.830 128.060 186.890 ;
        RECT 126.450 186.690 128.060 186.830 ;
        RECT 128.750 186.830 128.890 186.985 ;
        RECT 129.120 186.970 129.440 187.230 ;
        RECT 129.580 186.970 129.900 187.230 ;
        RECT 131.880 186.970 132.200 187.230 ;
        RECT 133.810 187.170 133.950 187.325 ;
        RECT 137.400 187.170 137.720 187.230 ;
        RECT 133.810 187.030 137.720 187.170 ;
        RECT 137.400 186.970 137.720 187.030 ;
        RECT 129.670 186.830 129.810 186.970 ;
        RECT 130.500 186.875 130.820 186.890 ;
        RECT 128.750 186.690 129.810 186.830 ;
        RECT 127.740 186.630 128.060 186.690 ;
        RECT 130.385 186.645 130.820 186.875 ;
        RECT 130.975 186.645 131.265 186.875 ;
        RECT 131.435 186.830 131.725 186.875 ;
        RECT 132.340 186.830 132.660 186.890 ;
        RECT 131.435 186.690 132.660 186.830 ;
        RECT 131.435 186.645 131.725 186.690 ;
        RECT 130.500 186.630 130.820 186.645 ;
        RECT 109.430 186.350 122.220 186.490 ;
        RECT 129.120 186.490 129.440 186.550 ;
        RECT 131.050 186.490 131.190 186.645 ;
        RECT 132.340 186.630 132.660 186.690 ;
        RECT 132.815 186.830 133.105 186.875 ;
        RECT 134.960 186.830 135.250 186.875 ;
        RECT 132.815 186.690 135.250 186.830 ;
        RECT 132.815 186.645 133.105 186.690 ;
        RECT 134.960 186.645 135.250 186.690 ;
        RECT 135.560 186.830 135.880 186.890 ;
        RECT 138.870 186.830 139.010 187.370 ;
        RECT 142.000 186.970 142.320 187.230 ;
        RECT 143.010 187.215 143.150 187.370 ;
        RECT 142.935 186.985 143.225 187.215 ;
        RECT 143.840 186.970 144.160 187.230 ;
        RECT 142.475 186.830 142.765 186.875 ;
        RECT 135.560 186.690 139.010 186.830 ;
        RECT 139.330 186.690 142.765 186.830 ;
        RECT 135.560 186.630 135.880 186.690 ;
        RECT 129.120 186.350 131.190 186.490 ;
        RECT 132.430 186.490 132.570 186.630 ;
        RECT 139.330 186.490 139.470 186.690 ;
        RECT 142.475 186.645 142.765 186.690 ;
        RECT 132.430 186.350 139.470 186.490 ;
        RECT 107.975 186.305 108.265 186.350 ;
        RECT 108.420 186.290 108.740 186.350 ;
        RECT 112.100 186.290 112.420 186.350 ;
        RECT 129.120 186.290 129.440 186.350 ;
        RECT 140.620 186.290 140.940 186.550 ;
        RECT 17.270 185.670 146.990 186.150 ;
        RECT 30.220 185.515 30.540 185.530 ;
        RECT 26.555 185.285 26.845 185.515 ;
        RECT 30.155 185.285 30.540 185.515 ;
        RECT 20.990 185.130 21.280 185.175 ;
        RECT 22.400 185.130 22.720 185.190 ;
        RECT 20.990 184.990 22.720 185.130 ;
        RECT 26.630 185.130 26.770 185.285 ;
        RECT 30.220 185.270 30.540 185.285 ;
        RECT 32.060 185.270 32.380 185.530 ;
        RECT 38.960 185.470 39.280 185.530 ;
        RECT 38.130 185.330 39.280 185.470 ;
        RECT 27.000 185.130 27.320 185.190 ;
        RECT 28.015 185.130 28.305 185.175 ;
        RECT 26.630 184.990 27.320 185.130 ;
        RECT 20.990 184.945 21.280 184.990 ;
        RECT 22.400 184.930 22.720 184.990 ;
        RECT 27.000 184.930 27.320 184.990 ;
        RECT 27.550 184.990 28.305 185.130 ;
        RECT 26.080 184.790 26.400 184.850 ;
        RECT 27.550 184.790 27.690 184.990 ;
        RECT 28.015 184.945 28.305 184.990 ;
        RECT 31.140 184.930 31.460 185.190 ;
        RECT 26.080 184.650 27.690 184.790 ;
        RECT 26.080 184.590 26.400 184.650 ;
        RECT 31.615 184.605 31.905 184.835 ;
        RECT 37.135 184.790 37.425 184.835 ;
        RECT 37.580 184.790 37.900 184.850 ;
        RECT 38.130 184.835 38.270 185.330 ;
        RECT 38.960 185.270 39.280 185.330 ;
        RECT 39.880 185.470 40.200 185.530 ;
        RECT 40.815 185.470 41.105 185.515 ;
        RECT 39.880 185.330 41.105 185.470 ;
        RECT 39.880 185.270 40.200 185.330 ;
        RECT 40.815 185.285 41.105 185.330 ;
        RECT 60.120 185.470 60.440 185.530 ;
        RECT 61.515 185.470 61.805 185.515 ;
        RECT 60.120 185.330 61.805 185.470 ;
        RECT 60.120 185.270 60.440 185.330 ;
        RECT 61.515 185.285 61.805 185.330 ;
        RECT 61.960 185.470 62.280 185.530 ;
        RECT 63.800 185.470 64.120 185.530 ;
        RECT 110.260 185.470 110.580 185.530 ;
        RECT 113.940 185.470 114.260 185.530 ;
        RECT 61.960 185.330 64.490 185.470 ;
        RECT 61.960 185.270 62.280 185.330 ;
        RECT 63.800 185.270 64.120 185.330 ;
        RECT 38.500 185.130 38.820 185.190 ;
        RECT 44.940 185.130 45.260 185.190 ;
        RECT 38.500 184.990 41.490 185.130 ;
        RECT 38.500 184.930 38.820 184.990 ;
        RECT 39.050 184.835 39.190 184.990 ;
        RECT 41.350 184.835 41.490 184.990 ;
        RECT 42.270 184.990 45.260 185.130 ;
        RECT 42.270 184.835 42.410 184.990 ;
        RECT 44.940 184.930 45.260 184.990 ;
        RECT 60.580 185.130 60.900 185.190 ;
        RECT 62.895 185.130 63.185 185.175 ;
        RECT 60.580 184.990 63.185 185.130 ;
        RECT 60.580 184.930 60.900 184.990 ;
        RECT 62.895 184.945 63.185 184.990 ;
        RECT 64.350 185.130 64.490 185.330 ;
        RECT 110.260 185.330 114.260 185.470 ;
        RECT 110.260 185.270 110.580 185.330 ;
        RECT 113.940 185.270 114.260 185.330 ;
        RECT 124.075 185.470 124.365 185.515 ;
        RECT 125.900 185.470 126.220 185.530 ;
        RECT 129.580 185.470 129.900 185.530 ;
        RECT 131.880 185.470 132.200 185.530 ;
        RECT 124.075 185.330 126.220 185.470 ;
        RECT 124.075 185.285 124.365 185.330 ;
        RECT 125.900 185.270 126.220 185.330 ;
        RECT 126.910 185.330 129.900 185.470 ;
        RECT 66.100 185.130 66.420 185.190 ;
        RECT 64.350 184.990 66.420 185.130 ;
        RECT 37.135 184.650 37.900 184.790 ;
        RECT 37.135 184.605 37.425 184.650 ;
        RECT 19.655 184.265 19.945 184.495 ;
        RECT 20.535 184.450 20.825 184.495 ;
        RECT 21.725 184.450 22.015 184.495 ;
        RECT 24.245 184.450 24.535 184.495 ;
        RECT 20.535 184.310 24.535 184.450 ;
        RECT 20.535 184.265 20.825 184.310 ;
        RECT 21.725 184.265 22.015 184.310 ;
        RECT 24.245 184.265 24.535 184.310 ;
        RECT 19.730 183.770 19.870 184.265 ;
        RECT 20.140 184.110 20.430 184.155 ;
        RECT 22.240 184.110 22.530 184.155 ;
        RECT 23.810 184.110 24.100 184.155 ;
        RECT 20.140 183.970 24.100 184.110 ;
        RECT 20.140 183.925 20.430 183.970 ;
        RECT 22.240 183.925 22.530 183.970 ;
        RECT 23.810 183.925 24.100 183.970 ;
        RECT 26.540 184.110 26.860 184.170 ;
        RECT 28.855 184.110 29.145 184.155 ;
        RECT 31.690 184.110 31.830 184.605 ;
        RECT 37.580 184.590 37.900 184.650 ;
        RECT 38.055 184.605 38.345 184.835 ;
        RECT 38.975 184.605 39.265 184.835 ;
        RECT 39.895 184.605 40.185 184.835 ;
        RECT 41.275 184.605 41.565 184.835 ;
        RECT 42.195 184.605 42.485 184.835 ;
        RECT 42.640 184.790 42.960 184.850 ;
        RECT 44.495 184.790 44.785 184.835 ;
        RECT 42.640 184.650 44.785 184.790 ;
        RECT 34.820 184.450 35.140 184.510 ;
        RECT 38.515 184.450 38.805 184.495 ;
        RECT 34.820 184.310 38.805 184.450 ;
        RECT 39.970 184.450 40.110 184.605 ;
        RECT 40.340 184.450 40.660 184.510 ;
        RECT 42.270 184.450 42.410 184.605 ;
        RECT 42.640 184.590 42.960 184.650 ;
        RECT 44.495 184.605 44.785 184.650 ;
        RECT 45.400 184.590 45.720 184.850 ;
        RECT 45.860 184.590 46.180 184.850 ;
        RECT 61.055 184.605 61.345 184.835 ;
        RECT 39.970 184.310 42.410 184.450 ;
        RECT 61.130 184.450 61.270 184.605 ;
        RECT 61.960 184.590 62.280 184.850 ;
        RECT 63.340 184.790 63.660 184.850 ;
        RECT 64.350 184.835 64.490 184.990 ;
        RECT 66.100 184.930 66.420 184.990 ;
        RECT 126.360 184.930 126.680 185.190 ;
        RECT 63.815 184.790 64.105 184.835 ;
        RECT 63.340 184.650 64.105 184.790 ;
        RECT 63.340 184.590 63.660 184.650 ;
        RECT 63.815 184.605 64.105 184.650 ;
        RECT 64.275 184.605 64.565 184.835 ;
        RECT 65.195 184.605 65.485 184.835 ;
        RECT 65.655 184.790 65.945 184.835 ;
        RECT 66.560 184.790 66.880 184.850 ;
        RECT 65.655 184.650 66.880 184.790 ;
        RECT 65.655 184.605 65.945 184.650 ;
        RECT 63.430 184.450 63.570 184.590 ;
        RECT 61.130 184.310 63.570 184.450 ;
        RECT 65.270 184.450 65.410 184.605 ;
        RECT 66.560 184.590 66.880 184.650 ;
        RECT 72.540 184.790 72.860 184.850 ;
        RECT 78.075 184.790 78.365 184.835 ;
        RECT 72.540 184.650 78.365 184.790 ;
        RECT 72.540 184.590 72.860 184.650 ;
        RECT 78.075 184.605 78.365 184.650 ;
        RECT 78.995 184.605 79.285 184.835 ;
        RECT 88.610 184.790 88.900 184.835 ;
        RECT 94.620 184.790 94.940 184.850 ;
        RECT 88.610 184.650 94.940 184.790 ;
        RECT 88.610 184.605 88.900 184.650 ;
        RECT 73.000 184.450 73.320 184.510 ;
        RECT 74.395 184.450 74.685 184.495 ;
        RECT 65.270 184.310 74.685 184.450 ;
        RECT 34.820 184.250 35.140 184.310 ;
        RECT 38.515 184.265 38.805 184.310 ;
        RECT 40.340 184.250 40.660 184.310 ;
        RECT 73.000 184.250 73.320 184.310 ;
        RECT 74.395 184.265 74.685 184.310 ;
        RECT 77.615 184.450 77.905 184.495 ;
        RECT 79.070 184.450 79.210 184.605 ;
        RECT 94.620 184.590 94.940 184.650 ;
        RECT 98.300 184.590 98.620 184.850 ;
        RECT 99.680 184.790 100.000 184.850 ;
        RECT 106.595 184.790 106.885 184.835 ;
        RECT 107.960 184.790 108.280 184.850 ;
        RECT 99.680 184.650 108.280 184.790 ;
        RECT 99.680 184.590 100.000 184.650 ;
        RECT 106.595 184.605 106.885 184.650 ;
        RECT 107.960 184.590 108.280 184.650 ;
        RECT 110.260 184.790 110.580 184.850 ;
        RECT 110.735 184.790 111.025 184.835 ;
        RECT 110.260 184.650 111.025 184.790 ;
        RECT 110.260 184.590 110.580 184.650 ;
        RECT 110.735 184.605 111.025 184.650 ;
        RECT 111.180 184.590 111.500 184.850 ;
        RECT 124.995 184.605 125.285 184.835 ;
        RECT 125.915 184.790 126.205 184.835 ;
        RECT 126.910 184.790 127.050 185.330 ;
        RECT 129.580 185.270 129.900 185.330 ;
        RECT 130.590 185.330 132.200 185.470 ;
        RECT 127.455 185.130 127.745 185.175 ;
        RECT 129.120 185.130 129.440 185.190 ;
        RECT 127.455 184.990 129.440 185.130 ;
        RECT 127.455 184.945 127.745 184.990 ;
        RECT 129.120 184.930 129.440 184.990 ;
        RECT 125.915 184.650 127.050 184.790 ;
        RECT 125.915 184.605 126.205 184.650 ;
        RECT 128.675 184.605 128.965 184.835 ;
        RECT 129.655 184.790 129.945 184.835 ;
        RECT 130.590 184.790 130.730 185.330 ;
        RECT 131.880 185.270 132.200 185.330 ;
        RECT 132.800 185.270 133.120 185.530 ;
        RECT 135.115 185.470 135.405 185.515 ;
        RECT 135.560 185.470 135.880 185.530 ;
        RECT 135.115 185.330 135.880 185.470 ;
        RECT 135.115 185.285 135.405 185.330 ;
        RECT 135.560 185.270 135.880 185.330 ;
        RECT 132.890 185.130 133.030 185.270 ;
        RECT 143.840 185.130 144.160 185.190 ;
        RECT 131.050 184.990 144.160 185.130 ;
        RECT 131.050 184.835 131.190 184.990 ;
        RECT 143.840 184.930 144.160 184.990 ;
        RECT 129.655 184.650 130.730 184.790 ;
        RECT 129.655 184.605 129.945 184.650 ;
        RECT 130.975 184.605 131.265 184.835 ;
        RECT 131.420 184.790 131.740 184.850 ;
        RECT 131.895 184.790 132.185 184.835 ;
        RECT 131.420 184.650 132.185 184.790 ;
        RECT 77.615 184.310 79.210 184.450 ;
        RECT 86.340 184.450 86.660 184.510 ;
        RECT 87.275 184.450 87.565 184.495 ;
        RECT 86.340 184.310 87.565 184.450 ;
        RECT 77.615 184.265 77.905 184.310 ;
        RECT 86.340 184.250 86.660 184.310 ;
        RECT 87.275 184.265 87.565 184.310 ;
        RECT 88.155 184.450 88.445 184.495 ;
        RECT 89.345 184.450 89.635 184.495 ;
        RECT 91.865 184.450 92.155 184.495 ;
        RECT 88.155 184.310 92.155 184.450 ;
        RECT 88.155 184.265 88.445 184.310 ;
        RECT 89.345 184.265 89.635 184.310 ;
        RECT 91.865 184.265 92.155 184.310 ;
        RECT 95.080 184.450 95.400 184.510 ;
        RECT 99.770 184.450 99.910 184.590 ;
        RECT 95.080 184.310 99.910 184.450 ;
        RECT 95.080 184.250 95.400 184.310 ;
        RECT 101.535 184.265 101.825 184.495 ;
        RECT 26.540 183.970 31.830 184.110 ;
        RECT 39.880 184.110 40.200 184.170 ;
        RECT 44.955 184.110 45.245 184.155 ;
        RECT 39.880 183.970 45.245 184.110 ;
        RECT 26.540 183.910 26.860 183.970 ;
        RECT 28.855 183.925 29.145 183.970 ;
        RECT 39.880 183.910 40.200 183.970 ;
        RECT 44.955 183.925 45.245 183.970 ;
        RECT 87.760 184.110 88.050 184.155 ;
        RECT 89.860 184.110 90.150 184.155 ;
        RECT 91.430 184.110 91.720 184.155 ;
        RECT 87.760 183.970 91.720 184.110 ;
        RECT 87.760 183.925 88.050 183.970 ;
        RECT 89.860 183.925 90.150 183.970 ;
        RECT 91.430 183.925 91.720 183.970 ;
        RECT 94.175 184.110 94.465 184.155 ;
        RECT 96.920 184.110 97.240 184.170 ;
        RECT 101.610 184.110 101.750 184.265 ;
        RECT 105.200 184.250 105.520 184.510 ;
        RECT 123.600 184.450 123.920 184.510 ;
        RECT 125.070 184.450 125.210 184.605 ;
        RECT 128.200 184.450 128.520 184.510 ;
        RECT 123.600 184.310 128.520 184.450 ;
        RECT 123.600 184.250 123.920 184.310 ;
        RECT 128.200 184.250 128.520 184.310 ;
        RECT 94.175 183.970 101.750 184.110 ;
        RECT 112.115 184.110 112.405 184.155 ;
        RECT 115.320 184.110 115.640 184.170 ;
        RECT 128.750 184.110 128.890 184.605 ;
        RECT 131.420 184.590 131.740 184.650 ;
        RECT 131.895 184.605 132.185 184.650 ;
        RECT 133.720 184.590 134.040 184.850 ;
        RECT 134.195 184.790 134.485 184.835 ;
        RECT 134.640 184.790 134.960 184.850 ;
        RECT 134.195 184.650 134.960 184.790 ;
        RECT 134.195 184.605 134.485 184.650 ;
        RECT 134.640 184.590 134.960 184.650 ;
        RECT 136.480 184.590 136.800 184.850 ;
        RECT 137.400 184.590 137.720 184.850 ;
        RECT 137.860 184.590 138.180 184.850 ;
        RECT 138.780 184.835 139.100 184.850 ;
        RECT 138.750 184.605 139.100 184.835 ;
        RECT 138.780 184.590 139.100 184.605 ;
        RECT 130.500 184.450 130.820 184.510 ;
        RECT 132.815 184.450 133.105 184.495 ;
        RECT 130.500 184.310 133.105 184.450 ;
        RECT 130.500 184.250 130.820 184.310 ;
        RECT 132.815 184.265 133.105 184.310 ;
        RECT 133.260 184.450 133.580 184.510 ;
        RECT 137.950 184.450 138.090 184.590 ;
        RECT 133.260 184.310 138.090 184.450 ;
        RECT 138.295 184.450 138.585 184.495 ;
        RECT 139.485 184.450 139.775 184.495 ;
        RECT 142.005 184.450 142.295 184.495 ;
        RECT 138.295 184.310 142.295 184.450 ;
        RECT 133.260 184.250 133.580 184.310 ;
        RECT 138.295 184.265 138.585 184.310 ;
        RECT 139.485 184.265 139.775 184.310 ;
        RECT 142.005 184.265 142.295 184.310 ;
        RECT 112.115 183.970 115.640 184.110 ;
        RECT 94.175 183.925 94.465 183.970 ;
        RECT 96.920 183.910 97.240 183.970 ;
        RECT 112.115 183.925 112.405 183.970 ;
        RECT 115.320 183.910 115.640 183.970 ;
        RECT 127.370 183.970 128.890 184.110 ;
        RECT 25.160 183.770 25.480 183.830 ;
        RECT 19.730 183.630 25.480 183.770 ;
        RECT 25.160 183.570 25.480 183.630 ;
        RECT 25.620 183.770 25.940 183.830 ;
        RECT 27.935 183.770 28.225 183.815 ;
        RECT 25.620 183.630 28.225 183.770 ;
        RECT 25.620 183.570 25.940 183.630 ;
        RECT 27.935 183.585 28.225 183.630 ;
        RECT 29.300 183.570 29.620 183.830 ;
        RECT 29.760 183.770 30.080 183.830 ;
        RECT 30.235 183.770 30.525 183.815 ;
        RECT 29.760 183.630 30.525 183.770 ;
        RECT 29.760 183.570 30.080 183.630 ;
        RECT 30.235 183.585 30.525 183.630 ;
        RECT 38.500 183.770 38.820 183.830 ;
        RECT 41.275 183.770 41.565 183.815 ;
        RECT 38.500 183.630 41.565 183.770 ;
        RECT 38.500 183.570 38.820 183.630 ;
        RECT 41.275 183.585 41.565 183.630 ;
        RECT 43.560 183.570 43.880 183.830 ;
        RECT 78.060 183.570 78.380 183.830 ;
        RECT 95.095 183.770 95.385 183.815 ;
        RECT 96.000 183.770 96.320 183.830 ;
        RECT 95.095 183.630 96.320 183.770 ;
        RECT 95.095 183.585 95.385 183.630 ;
        RECT 96.000 183.570 96.320 183.630 ;
        RECT 97.380 183.770 97.700 183.830 ;
        RECT 98.775 183.770 99.065 183.815 ;
        RECT 97.380 183.630 99.065 183.770 ;
        RECT 97.380 183.570 97.700 183.630 ;
        RECT 98.775 183.585 99.065 183.630 ;
        RECT 102.455 183.770 102.745 183.815 ;
        RECT 102.900 183.770 103.220 183.830 ;
        RECT 102.455 183.630 103.220 183.770 ;
        RECT 102.455 183.585 102.745 183.630 ;
        RECT 102.900 183.570 103.220 183.630 ;
        RECT 105.660 183.770 105.980 183.830 ;
        RECT 109.355 183.770 109.645 183.815 ;
        RECT 105.660 183.630 109.645 183.770 ;
        RECT 105.660 183.570 105.980 183.630 ;
        RECT 109.355 183.585 109.645 183.630 ;
        RECT 126.820 183.770 127.140 183.830 ;
        RECT 127.370 183.815 127.510 183.970 ;
        RECT 127.295 183.770 127.585 183.815 ;
        RECT 126.820 183.630 127.585 183.770 ;
        RECT 126.820 183.570 127.140 183.630 ;
        RECT 127.295 183.585 127.585 183.630 ;
        RECT 127.740 183.770 128.060 183.830 ;
        RECT 128.215 183.770 128.505 183.815 ;
        RECT 127.740 183.630 128.505 183.770 ;
        RECT 128.750 183.770 128.890 183.970 ;
        RECT 129.595 184.110 129.885 184.155 ;
        RECT 130.040 184.110 130.360 184.170 ;
        RECT 129.595 183.970 130.360 184.110 ;
        RECT 129.595 183.925 129.885 183.970 ;
        RECT 130.040 183.910 130.360 183.970 ;
        RECT 132.340 184.110 132.660 184.170 ;
        RECT 135.560 184.110 135.880 184.170 ;
        RECT 132.340 183.970 135.880 184.110 ;
        RECT 132.340 183.910 132.660 183.970 ;
        RECT 135.560 183.910 135.880 183.970 ;
        RECT 137.900 184.110 138.190 184.155 ;
        RECT 140.000 184.110 140.290 184.155 ;
        RECT 141.570 184.110 141.860 184.155 ;
        RECT 137.900 183.970 141.860 184.110 ;
        RECT 137.900 183.925 138.190 183.970 ;
        RECT 140.000 183.925 140.290 183.970 ;
        RECT 141.570 183.925 141.860 183.970 ;
        RECT 131.880 183.770 132.200 183.830 ;
        RECT 136.020 183.770 136.340 183.830 ;
        RECT 128.750 183.630 136.340 183.770 ;
        RECT 127.740 183.570 128.060 183.630 ;
        RECT 128.215 183.585 128.505 183.630 ;
        RECT 131.880 183.570 132.200 183.630 ;
        RECT 136.020 183.570 136.340 183.630 ;
        RECT 136.480 183.770 136.800 183.830 ;
        RECT 144.315 183.770 144.605 183.815 ;
        RECT 136.480 183.630 144.605 183.770 ;
        RECT 136.480 183.570 136.800 183.630 ;
        RECT 144.315 183.585 144.605 183.630 ;
        RECT 17.270 182.950 146.990 183.430 ;
        RECT 21.955 182.750 22.245 182.795 ;
        RECT 25.620 182.750 25.940 182.810 ;
        RECT 21.955 182.610 25.940 182.750 ;
        RECT 21.955 182.565 22.245 182.610 ;
        RECT 25.620 182.550 25.940 182.610 ;
        RECT 44.955 182.750 45.245 182.795 ;
        RECT 45.860 182.750 46.180 182.810 ;
        RECT 44.955 182.610 46.180 182.750 ;
        RECT 44.955 182.565 45.245 182.610 ;
        RECT 45.860 182.550 46.180 182.610 ;
        RECT 65.180 182.750 65.500 182.810 ;
        RECT 66.560 182.750 66.880 182.810 ;
        RECT 65.180 182.610 66.880 182.750 ;
        RECT 65.180 182.550 65.500 182.610 ;
        RECT 66.560 182.550 66.880 182.610 ;
        RECT 73.000 182.550 73.320 182.810 ;
        RECT 93.255 182.750 93.545 182.795 ;
        RECT 98.300 182.750 98.620 182.810 ;
        RECT 93.255 182.610 98.620 182.750 ;
        RECT 93.255 182.565 93.545 182.610 ;
        RECT 98.300 182.550 98.620 182.610 ;
        RECT 114.875 182.750 115.165 182.795 ;
        RECT 115.320 182.750 115.640 182.810 ;
        RECT 114.875 182.610 115.640 182.750 ;
        RECT 114.875 182.565 115.165 182.610 ;
        RECT 115.320 182.550 115.640 182.610 ;
        RECT 123.600 182.550 123.920 182.810 ;
        RECT 129.120 182.750 129.440 182.810 ;
        RECT 133.735 182.750 134.025 182.795 ;
        RECT 129.120 182.610 134.025 182.750 ;
        RECT 129.120 182.550 129.440 182.610 ;
        RECT 133.735 182.565 134.025 182.610 ;
        RECT 135.035 182.610 137.170 182.750 ;
        RECT 24.700 182.410 24.990 182.455 ;
        RECT 26.270 182.410 26.560 182.455 ;
        RECT 28.370 182.410 28.660 182.455 ;
        RECT 24.700 182.270 28.660 182.410 ;
        RECT 24.700 182.225 24.990 182.270 ;
        RECT 26.270 182.225 26.560 182.270 ;
        RECT 28.370 182.225 28.660 182.270 ;
        RECT 38.500 182.210 38.820 182.470 ;
        RECT 38.975 182.410 39.265 182.455 ;
        RECT 39.880 182.410 40.200 182.470 ;
        RECT 46.335 182.410 46.625 182.455 ;
        RECT 38.975 182.270 40.200 182.410 ;
        RECT 38.975 182.225 39.265 182.270 ;
        RECT 39.880 182.210 40.200 182.270 ;
        RECT 41.810 182.270 46.625 182.410 ;
        RECT 41.810 182.115 41.950 182.270 ;
        RECT 24.265 182.070 24.555 182.115 ;
        RECT 26.785 182.070 27.075 182.115 ;
        RECT 27.975 182.070 28.265 182.115 ;
        RECT 24.265 181.930 28.265 182.070 ;
        RECT 24.265 181.885 24.555 181.930 ;
        RECT 26.785 181.885 27.075 181.930 ;
        RECT 27.975 181.885 28.265 181.930 ;
        RECT 41.735 181.885 42.025 182.115 ;
        RECT 43.560 181.870 43.880 182.130 ;
        RECT 25.160 181.730 25.480 181.790 ;
        RECT 28.855 181.730 29.145 181.775 ;
        RECT 25.160 181.590 29.145 181.730 ;
        RECT 25.160 181.530 25.480 181.590 ;
        RECT 28.855 181.545 29.145 181.590 ;
        RECT 38.040 181.530 38.360 181.790 ;
        RECT 39.420 181.530 39.740 181.790 ;
        RECT 42.195 181.730 42.485 181.775 ;
        RECT 43.100 181.730 43.420 181.790 ;
        RECT 45.490 181.775 45.630 182.270 ;
        RECT 46.335 182.225 46.625 182.270 ;
        RECT 49.080 182.410 49.370 182.455 ;
        RECT 50.650 182.410 50.940 182.455 ;
        RECT 52.750 182.410 53.040 182.455 ;
        RECT 49.080 182.270 53.040 182.410 ;
        RECT 49.080 182.225 49.370 182.270 ;
        RECT 50.650 182.225 50.940 182.270 ;
        RECT 52.750 182.225 53.040 182.270 ;
        RECT 58.280 182.410 58.600 182.470 ;
        RECT 67.955 182.410 68.245 182.455 ;
        RECT 72.555 182.410 72.845 182.455 ;
        RECT 58.280 182.270 68.245 182.410 ;
        RECT 58.280 182.210 58.600 182.270 ;
        RECT 67.955 182.225 68.245 182.270 ;
        RECT 68.490 182.270 72.845 182.410 ;
        RECT 48.645 182.070 48.935 182.115 ;
        RECT 51.165 182.070 51.455 182.115 ;
        RECT 52.355 182.070 52.645 182.115 ;
        RECT 68.490 182.070 68.630 182.270 ;
        RECT 72.555 182.225 72.845 182.270 ;
        RECT 48.645 181.930 52.645 182.070 ;
        RECT 48.645 181.885 48.935 181.930 ;
        RECT 51.165 181.885 51.455 181.930 ;
        RECT 52.355 181.885 52.645 181.930 ;
        RECT 66.650 181.930 68.630 182.070 ;
        RECT 70.715 182.070 71.005 182.115 ;
        RECT 73.090 182.070 73.230 182.550 ;
        RECT 75.760 182.410 76.050 182.455 ;
        RECT 77.330 182.410 77.620 182.455 ;
        RECT 79.430 182.410 79.720 182.455 ;
        RECT 75.760 182.270 79.720 182.410 ;
        RECT 75.760 182.225 76.050 182.270 ;
        RECT 77.330 182.225 77.620 182.270 ;
        RECT 79.430 182.225 79.720 182.270 ;
        RECT 86.840 182.410 87.130 182.455 ;
        RECT 88.940 182.410 89.230 182.455 ;
        RECT 90.510 182.410 90.800 182.455 ;
        RECT 86.840 182.270 90.800 182.410 ;
        RECT 86.840 182.225 87.130 182.270 ;
        RECT 88.940 182.225 89.230 182.270 ;
        RECT 90.510 182.225 90.800 182.270 ;
        RECT 108.460 182.410 108.750 182.455 ;
        RECT 110.560 182.410 110.850 182.455 ;
        RECT 112.130 182.410 112.420 182.455 ;
        RECT 133.260 182.410 133.580 182.470 ;
        RECT 108.460 182.270 112.420 182.410 ;
        RECT 108.460 182.225 108.750 182.270 ;
        RECT 110.560 182.225 110.850 182.270 ;
        RECT 112.130 182.225 112.420 182.270 ;
        RECT 131.510 182.270 133.580 182.410 ;
        RECT 70.715 181.930 73.230 182.070 ;
        RECT 75.325 182.070 75.615 182.115 ;
        RECT 77.845 182.070 78.135 182.115 ;
        RECT 79.035 182.070 79.325 182.115 ;
        RECT 75.325 181.930 79.325 182.070 ;
        RECT 66.650 181.790 66.790 181.930 ;
        RECT 70.715 181.885 71.005 181.930 ;
        RECT 75.325 181.885 75.615 181.930 ;
        RECT 77.845 181.885 78.135 181.930 ;
        RECT 79.035 181.885 79.325 181.930 ;
        RECT 87.235 182.070 87.525 182.115 ;
        RECT 88.425 182.070 88.715 182.115 ;
        RECT 90.945 182.070 91.235 182.115 ;
        RECT 87.235 181.930 91.235 182.070 ;
        RECT 87.235 181.885 87.525 181.930 ;
        RECT 88.425 181.885 88.715 181.930 ;
        RECT 90.945 181.885 91.235 181.930 ;
        RECT 96.000 181.870 96.320 182.130 ;
        RECT 96.935 182.070 97.225 182.115 ;
        RECT 98.300 182.070 98.620 182.130 ;
        RECT 101.060 182.070 101.380 182.130 ;
        RECT 96.935 181.930 101.380 182.070 ;
        RECT 96.935 181.885 97.225 181.930 ;
        RECT 98.300 181.870 98.620 181.930 ;
        RECT 101.060 181.870 101.380 181.930 ;
        RECT 102.900 181.870 103.220 182.130 ;
        RECT 103.835 182.070 104.125 182.115 ;
        RECT 103.835 181.930 107.730 182.070 ;
        RECT 103.835 181.885 104.125 181.930 ;
        RECT 44.495 181.730 44.785 181.775 ;
        RECT 42.195 181.590 44.785 181.730 ;
        RECT 42.195 181.545 42.485 181.590 ;
        RECT 43.100 181.530 43.420 181.590 ;
        RECT 44.495 181.545 44.785 181.590 ;
        RECT 45.415 181.730 45.705 181.775 ;
        RECT 48.160 181.730 48.480 181.790 ;
        RECT 45.415 181.590 48.480 181.730 ;
        RECT 45.415 181.545 45.705 181.590 ;
        RECT 48.160 181.530 48.480 181.590 ;
        RECT 52.760 181.730 53.080 181.790 ;
        RECT 53.235 181.730 53.525 181.775 ;
        RECT 66.560 181.730 66.880 181.790 ;
        RECT 52.760 181.590 53.525 181.730 ;
        RECT 52.760 181.530 53.080 181.590 ;
        RECT 53.235 181.545 53.525 181.590 ;
        RECT 65.730 181.590 66.880 181.730 ;
        RECT 27.630 181.390 27.920 181.435 ;
        RECT 29.300 181.390 29.620 181.450 ;
        RECT 27.630 181.250 29.620 181.390 ;
        RECT 27.630 181.205 27.920 181.250 ;
        RECT 29.300 181.190 29.620 181.250 ;
        RECT 43.560 181.390 43.880 181.450 ;
        RECT 51.840 181.435 52.160 181.450 ;
        RECT 44.035 181.390 44.325 181.435 ;
        RECT 43.560 181.250 44.325 181.390 ;
        RECT 43.560 181.190 43.880 181.250 ;
        RECT 44.035 181.205 44.325 181.250 ;
        RECT 51.840 181.205 52.190 181.435 ;
        RECT 61.040 181.390 61.360 181.450 ;
        RECT 65.035 181.390 65.325 181.435 ;
        RECT 65.730 181.390 65.870 181.590 ;
        RECT 66.560 181.530 66.880 181.590 ;
        RECT 68.400 181.530 68.720 181.790 ;
        RECT 69.335 181.545 69.625 181.775 ;
        RECT 71.635 181.730 71.925 181.775 ;
        RECT 72.540 181.730 72.860 181.790 ;
        RECT 71.635 181.590 72.860 181.730 ;
        RECT 71.635 181.545 71.925 181.590 ;
        RECT 61.040 181.250 65.870 181.390 ;
        RECT 66.100 181.390 66.420 181.450 ;
        RECT 67.035 181.390 67.325 181.435 ;
        RECT 66.100 181.250 67.325 181.390 ;
        RECT 51.840 181.190 52.160 181.205 ;
        RECT 61.040 181.190 61.360 181.250 ;
        RECT 65.035 181.205 65.325 181.250 ;
        RECT 66.100 181.190 66.420 181.250 ;
        RECT 67.035 181.205 67.325 181.250 ;
        RECT 67.940 181.190 68.260 181.450 ;
        RECT 69.410 181.390 69.550 181.545 ;
        RECT 72.540 181.530 72.860 181.590 ;
        RECT 79.915 181.730 80.205 181.775 ;
        RECT 83.580 181.730 83.900 181.790 ;
        RECT 86.340 181.730 86.660 181.790 ;
        RECT 79.915 181.590 86.660 181.730 ;
        RECT 79.915 181.545 80.205 181.590 ;
        RECT 83.580 181.530 83.900 181.590 ;
        RECT 86.340 181.530 86.660 181.590 ;
        RECT 105.660 181.530 105.980 181.790 ;
        RECT 106.580 181.530 106.900 181.790 ;
        RECT 107.590 181.730 107.730 181.930 ;
        RECT 107.960 181.870 108.280 182.130 ;
        RECT 108.855 182.070 109.145 182.115 ;
        RECT 110.045 182.070 110.335 182.115 ;
        RECT 112.565 182.070 112.855 182.115 ;
        RECT 108.855 181.930 112.855 182.070 ;
        RECT 108.855 181.885 109.145 181.930 ;
        RECT 110.045 181.885 110.335 181.930 ;
        RECT 112.565 181.885 112.855 181.930 ;
        RECT 114.400 181.730 114.720 181.790 ;
        RECT 107.590 181.590 114.720 181.730 ;
        RECT 114.400 181.530 114.720 181.590 ;
        RECT 123.155 181.545 123.445 181.775 ;
        RECT 123.600 181.730 123.920 181.790 ;
        RECT 124.075 181.730 124.365 181.775 ;
        RECT 123.600 181.590 124.365 181.730 ;
        RECT 68.490 181.250 69.550 181.390 ;
        RECT 74.380 181.390 74.700 181.450 ;
        RECT 78.580 181.390 78.870 181.435 ;
        RECT 74.380 181.250 78.870 181.390 ;
        RECT 40.340 180.850 40.660 181.110 ;
        RECT 40.815 181.050 41.105 181.095 ;
        RECT 41.260 181.050 41.580 181.110 ;
        RECT 40.815 180.910 41.580 181.050 ;
        RECT 40.815 180.865 41.105 180.910 ;
        RECT 41.260 180.850 41.580 180.910 ;
        RECT 63.340 181.050 63.660 181.110 ;
        RECT 64.275 181.050 64.565 181.095 ;
        RECT 63.340 180.910 64.565 181.050 ;
        RECT 63.340 180.850 63.660 180.910 ;
        RECT 64.275 180.865 64.565 180.910 ;
        RECT 67.480 181.050 67.800 181.110 ;
        RECT 68.490 181.050 68.630 181.250 ;
        RECT 74.380 181.190 74.700 181.250 ;
        RECT 78.580 181.205 78.870 181.250 ;
        RECT 87.690 181.390 87.980 181.435 ;
        RECT 106.135 181.390 106.425 181.435 ;
        RECT 109.200 181.390 109.490 181.435 ;
        RECT 87.690 181.250 93.930 181.390 ;
        RECT 87.690 181.205 87.980 181.250 ;
        RECT 67.480 180.910 68.630 181.050 ;
        RECT 67.480 180.850 67.800 180.910 ;
        RECT 68.860 180.850 69.180 181.110 ;
        RECT 93.790 181.095 93.930 181.250 ;
        RECT 106.135 181.250 109.490 181.390 ;
        RECT 123.230 181.390 123.370 181.545 ;
        RECT 123.600 181.530 123.920 181.590 ;
        RECT 124.075 181.545 124.365 181.590 ;
        RECT 128.200 181.730 128.520 181.790 ;
        RECT 131.510 181.775 131.650 182.270 ;
        RECT 133.260 182.210 133.580 182.270 ;
        RECT 135.035 182.070 135.175 182.610 ;
        RECT 136.020 182.410 136.340 182.470 ;
        RECT 136.020 182.270 136.710 182.410 ;
        RECT 136.020 182.210 136.340 182.270 ;
        RECT 134.730 181.930 135.175 182.070 ;
        RECT 130.515 181.730 130.805 181.775 ;
        RECT 128.200 181.590 130.805 181.730 ;
        RECT 128.200 181.530 128.520 181.590 ;
        RECT 130.515 181.545 130.805 181.590 ;
        RECT 131.435 181.545 131.725 181.775 ;
        RECT 131.880 181.530 132.200 181.790 ;
        RECT 132.815 181.730 133.105 181.775 ;
        RECT 133.260 181.730 133.580 181.790 ;
        RECT 132.815 181.590 133.580 181.730 ;
        RECT 132.815 181.545 133.105 181.590 ;
        RECT 133.260 181.530 133.580 181.590 ;
        RECT 133.720 181.530 134.040 181.790 ;
        RECT 134.180 181.730 134.500 181.790 ;
        RECT 134.730 181.775 134.870 181.930 ;
        RECT 134.655 181.730 134.945 181.775 ;
        RECT 134.180 181.590 134.945 181.730 ;
        RECT 134.180 181.530 134.500 181.590 ;
        RECT 134.655 181.545 134.945 181.590 ;
        RECT 135.560 181.730 135.880 181.790 ;
        RECT 136.035 181.730 136.325 181.775 ;
        RECT 135.560 181.590 136.325 181.730 ;
        RECT 136.570 181.730 136.710 182.270 ;
        RECT 137.030 182.070 137.170 182.610 ;
        RECT 138.780 182.550 139.100 182.810 ;
        RECT 137.860 182.410 138.180 182.470 ;
        RECT 137.860 182.270 140.390 182.410 ;
        RECT 137.860 182.210 138.180 182.270 ;
        RECT 139.715 182.070 140.005 182.115 ;
        RECT 137.030 181.930 140.005 182.070 ;
        RECT 139.715 181.885 140.005 181.930 ;
        RECT 140.250 182.070 140.390 182.270 ;
        RECT 141.095 182.070 141.385 182.115 ;
        RECT 140.250 181.930 141.385 182.070 ;
        RECT 137.415 181.730 137.705 181.775 ;
        RECT 136.570 181.590 137.705 181.730 ;
        RECT 135.560 181.530 135.880 181.590 ;
        RECT 136.035 181.545 136.325 181.590 ;
        RECT 137.415 181.545 137.705 181.590 ;
        RECT 125.440 181.390 125.760 181.450 ;
        RECT 132.355 181.390 132.645 181.435 ;
        RECT 136.955 181.390 137.245 181.435 ;
        RECT 123.230 181.250 131.650 181.390 ;
        RECT 106.135 181.205 106.425 181.250 ;
        RECT 109.200 181.205 109.490 181.250 ;
        RECT 125.440 181.190 125.760 181.250 ;
        RECT 93.715 180.865 94.005 181.095 ;
        RECT 95.540 180.850 95.860 181.110 ;
        RECT 96.000 181.050 96.320 181.110 ;
        RECT 100.615 181.050 100.905 181.095 ;
        RECT 96.000 180.910 100.905 181.050 ;
        RECT 96.000 180.850 96.320 180.910 ;
        RECT 100.615 180.865 100.905 180.910 ;
        RECT 102.455 181.050 102.745 181.095 ;
        RECT 113.940 181.050 114.260 181.110 ;
        RECT 102.455 180.910 114.260 181.050 ;
        RECT 102.455 180.865 102.745 180.910 ;
        RECT 113.940 180.850 114.260 180.910 ;
        RECT 124.060 181.050 124.380 181.110 ;
        RECT 126.360 181.050 126.680 181.110 ;
        RECT 128.200 181.050 128.520 181.110 ;
        RECT 124.060 180.910 128.520 181.050 ;
        RECT 124.060 180.850 124.380 180.910 ;
        RECT 126.360 180.850 126.680 180.910 ;
        RECT 128.200 180.850 128.520 180.910 ;
        RECT 128.660 181.050 128.980 181.110 ;
        RECT 130.975 181.050 131.265 181.095 ;
        RECT 128.660 180.910 131.265 181.050 ;
        RECT 131.510 181.050 131.650 181.250 ;
        RECT 132.355 181.250 137.245 181.390 ;
        RECT 137.490 181.390 137.630 181.545 ;
        RECT 137.860 181.530 138.180 181.790 ;
        RECT 140.250 181.775 140.390 181.930 ;
        RECT 141.095 181.885 141.385 181.930 ;
        RECT 140.175 181.545 140.465 181.775 ;
        RECT 140.620 181.530 140.940 181.790 ;
        RECT 141.555 181.545 141.845 181.775 ;
        RECT 138.320 181.390 138.640 181.450 ;
        RECT 141.630 181.390 141.770 181.545 ;
        RECT 137.490 181.250 141.770 181.390 ;
        RECT 132.355 181.205 132.645 181.250 ;
        RECT 136.955 181.205 137.245 181.250 ;
        RECT 138.320 181.190 138.640 181.250 ;
        RECT 132.800 181.050 133.120 181.110 ;
        RECT 131.510 180.910 133.120 181.050 ;
        RECT 128.660 180.850 128.980 180.910 ;
        RECT 130.975 180.865 131.265 180.910 ;
        RECT 132.800 180.850 133.120 180.910 ;
        RECT 17.270 180.230 146.990 180.710 ;
        RECT 37.120 179.830 37.440 180.090 ;
        RECT 38.040 179.830 38.360 180.090 ;
        RECT 39.880 180.030 40.200 180.090 ;
        RECT 40.355 180.030 40.645 180.075 ;
        RECT 39.880 179.890 40.645 180.030 ;
        RECT 39.880 179.830 40.200 179.890 ;
        RECT 40.355 179.845 40.645 179.890 ;
        RECT 43.560 179.830 43.880 180.090 ;
        RECT 51.840 180.030 52.160 180.090 ;
        RECT 52.315 180.030 52.605 180.075 ;
        RECT 51.840 179.890 52.605 180.030 ;
        RECT 51.840 179.830 52.160 179.890 ;
        RECT 52.315 179.845 52.605 179.890 ;
        RECT 56.900 180.030 57.220 180.090 ;
        RECT 67.480 180.030 67.800 180.090 ;
        RECT 56.900 179.890 67.800 180.030 ;
        RECT 56.900 179.830 57.220 179.890 ;
        RECT 67.480 179.830 67.800 179.890 ;
        RECT 67.940 180.030 68.260 180.090 ;
        RECT 69.335 180.030 69.625 180.075 ;
        RECT 78.060 180.030 78.380 180.090 ;
        RECT 67.940 179.890 69.625 180.030 ;
        RECT 67.940 179.830 68.260 179.890 ;
        RECT 69.335 179.845 69.625 179.890 ;
        RECT 74.470 179.890 78.380 180.030 ;
        RECT 39.435 179.690 39.725 179.735 ;
        RECT 66.100 179.690 66.420 179.750 ;
        RECT 37.670 179.550 39.725 179.690 ;
        RECT 34.820 179.150 35.140 179.410 ;
        RECT 36.200 179.350 36.520 179.410 ;
        RECT 37.150 179.350 37.440 179.395 ;
        RECT 37.670 179.350 37.810 179.550 ;
        RECT 39.435 179.505 39.725 179.550 ;
        RECT 60.670 179.550 66.420 179.690 ;
        RECT 67.570 179.690 67.710 179.830 ;
        RECT 73.015 179.690 73.305 179.735 ;
        RECT 73.460 179.690 73.780 179.750 ;
        RECT 67.570 179.550 73.780 179.690 ;
        RECT 36.200 179.210 37.810 179.350 ;
        RECT 36.200 179.150 36.520 179.210 ;
        RECT 37.150 179.165 37.440 179.210 ;
        RECT 38.500 179.150 38.820 179.410 ;
        RECT 40.340 179.350 40.660 179.410 ;
        RECT 44.955 179.350 45.245 179.395 ;
        RECT 40.340 179.210 45.245 179.350 ;
        RECT 40.340 179.150 40.660 179.210 ;
        RECT 44.955 179.165 45.245 179.210 ;
        RECT 48.160 179.150 48.480 179.410 ;
        RECT 51.395 179.350 51.685 179.395 ;
        RECT 50.090 179.210 51.685 179.350 ;
        RECT 44.480 178.810 44.800 179.070 ;
        RECT 45.400 179.010 45.720 179.070 ;
        RECT 46.335 179.010 46.625 179.055 ;
        RECT 45.400 178.870 46.625 179.010 ;
        RECT 45.400 178.810 45.720 178.870 ;
        RECT 46.335 178.825 46.625 178.870 ;
        RECT 46.780 178.810 47.100 179.070 ;
        RECT 48.620 178.810 48.940 179.070 ;
        RECT 50.090 179.055 50.230 179.210 ;
        RECT 51.395 179.165 51.685 179.210 ;
        RECT 58.280 179.150 58.600 179.410 ;
        RECT 60.670 179.395 60.810 179.550 ;
        RECT 66.100 179.490 66.420 179.550 ;
        RECT 73.015 179.505 73.305 179.550 ;
        RECT 73.460 179.490 73.780 179.550 ;
        RECT 60.595 179.165 60.885 179.395 ;
        RECT 62.895 179.350 63.185 179.395 ;
        RECT 65.195 179.350 65.485 179.395 ;
        RECT 62.895 179.210 65.485 179.350 ;
        RECT 62.895 179.165 63.185 179.210 ;
        RECT 65.195 179.165 65.485 179.210 ;
        RECT 66.560 179.350 66.880 179.410 ;
        RECT 74.470 179.395 74.610 179.890 ;
        RECT 78.060 179.830 78.380 179.890 ;
        RECT 94.620 180.030 94.940 180.090 ;
        RECT 95.095 180.030 95.385 180.075 ;
        RECT 94.620 179.890 95.385 180.030 ;
        RECT 94.620 179.830 94.940 179.890 ;
        RECT 95.095 179.845 95.385 179.890 ;
        RECT 97.380 179.830 97.700 180.090 ;
        RECT 108.420 180.030 108.740 180.090 ;
        RECT 110.720 180.030 111.040 180.090 ;
        RECT 114.860 180.030 115.180 180.090 ;
        RECT 108.420 179.890 109.415 180.030 ;
        RECT 108.420 179.830 108.740 179.890 ;
        RECT 83.580 179.690 83.900 179.750 ;
        RECT 109.275 179.735 109.415 179.890 ;
        RECT 110.720 179.890 115.180 180.030 ;
        RECT 110.720 179.830 111.040 179.890 ;
        RECT 114.860 179.830 115.180 179.890 ;
        RECT 126.360 180.030 126.680 180.090 ;
        RECT 129.120 180.030 129.440 180.090 ;
        RECT 126.360 179.890 127.050 180.030 ;
        RECT 126.360 179.830 126.680 179.890 ;
        RECT 77.690 179.550 83.900 179.690 ;
        RECT 77.690 179.395 77.830 179.550 ;
        RECT 83.580 179.490 83.900 179.550 ;
        RECT 109.200 179.505 109.490 179.735 ;
        RECT 126.910 179.690 127.050 179.890 ;
        RECT 127.830 179.890 129.440 180.030 ;
        RECT 127.295 179.690 127.585 179.735 ;
        RECT 126.910 179.550 127.585 179.690 ;
        RECT 127.295 179.505 127.585 179.550 ;
        RECT 66.560 179.220 73.920 179.350 ;
        RECT 66.560 179.210 74.150 179.220 ;
        RECT 66.560 179.150 66.880 179.210 ;
        RECT 73.780 179.080 74.150 179.210 ;
        RECT 74.395 179.165 74.685 179.395 ;
        RECT 77.615 179.165 77.905 179.395 ;
        RECT 78.060 179.350 78.380 179.410 ;
        RECT 78.895 179.350 79.185 179.395 ;
        RECT 78.060 179.210 79.185 179.350 ;
        RECT 78.060 179.150 78.380 179.210 ;
        RECT 78.895 179.165 79.185 179.210 ;
        RECT 96.920 179.150 97.240 179.410 ;
        RECT 100.600 179.350 100.920 179.410 ;
        RECT 101.075 179.350 101.365 179.395 ;
        RECT 100.600 179.210 101.365 179.350 ;
        RECT 100.600 179.150 100.920 179.210 ;
        RECT 101.075 179.165 101.365 179.210 ;
        RECT 105.215 179.350 105.505 179.395 ;
        RECT 107.960 179.350 108.280 179.410 ;
        RECT 105.215 179.210 108.280 179.350 ;
        RECT 105.215 179.165 105.505 179.210 ;
        RECT 107.960 179.150 108.280 179.210 ;
        RECT 115.320 179.350 115.640 179.410 ;
        RECT 117.620 179.350 117.940 179.410 ;
        RECT 118.095 179.350 118.385 179.395 ;
        RECT 115.320 179.210 118.385 179.350 ;
        RECT 115.320 179.150 115.640 179.210 ;
        RECT 117.620 179.150 117.940 179.210 ;
        RECT 118.095 179.165 118.385 179.210 ;
        RECT 118.540 179.150 118.860 179.410 ;
        RECT 126.360 179.150 126.680 179.410 ;
        RECT 127.830 179.395 127.970 179.890 ;
        RECT 129.120 179.830 129.440 179.890 ;
        RECT 129.580 180.030 129.900 180.090 ;
        RECT 133.260 180.030 133.580 180.090 ;
        RECT 136.035 180.030 136.325 180.075 ;
        RECT 129.580 179.890 132.110 180.030 ;
        RECT 129.580 179.830 129.900 179.890 ;
        RECT 130.500 179.690 130.820 179.750 ;
        RECT 128.750 179.550 130.820 179.690 ;
        RECT 127.755 179.165 128.045 179.395 ;
        RECT 128.200 179.150 128.520 179.410 ;
        RECT 50.015 178.825 50.305 179.055 ;
        RECT 50.460 178.810 50.780 179.070 ;
        RECT 56.900 178.810 57.220 179.070 ;
        RECT 61.040 178.810 61.360 179.070 ;
        RECT 63.340 178.810 63.660 179.070 ;
        RECT 65.640 179.010 65.960 179.070 ;
        RECT 67.955 179.010 68.245 179.055 ;
        RECT 72.095 179.010 72.385 179.055 ;
        RECT 65.640 178.870 68.245 179.010 ;
        RECT 65.640 178.810 65.960 178.870 ;
        RECT 67.955 178.825 68.245 178.870 ;
        RECT 68.950 178.870 72.385 179.010 ;
        RECT 57.835 178.670 58.125 178.715 ;
        RECT 63.430 178.670 63.570 178.810 ;
        RECT 57.835 178.530 63.570 178.670 ;
        RECT 64.735 178.670 65.025 178.715 ;
        RECT 68.400 178.670 68.720 178.730 ;
        RECT 64.735 178.530 68.720 178.670 ;
        RECT 57.835 178.485 58.125 178.530 ;
        RECT 64.735 178.485 65.025 178.530 ;
        RECT 68.400 178.470 68.720 178.530 ;
        RECT 35.295 178.330 35.585 178.375 ;
        RECT 38.960 178.330 39.280 178.390 ;
        RECT 45.860 178.330 46.180 178.390 ;
        RECT 53.220 178.330 53.540 178.390 ;
        RECT 35.295 178.190 53.540 178.330 ;
        RECT 35.295 178.145 35.585 178.190 ;
        RECT 38.960 178.130 39.280 178.190 ;
        RECT 45.860 178.130 46.180 178.190 ;
        RECT 53.220 178.130 53.540 178.190 ;
        RECT 58.280 178.130 58.600 178.390 ;
        RECT 58.740 178.330 59.060 178.390 ;
        RECT 59.215 178.330 59.505 178.375 ;
        RECT 58.740 178.190 59.505 178.330 ;
        RECT 58.740 178.130 59.060 178.190 ;
        RECT 59.215 178.145 59.505 178.190 ;
        RECT 65.180 178.330 65.500 178.390 ;
        RECT 68.950 178.330 69.090 178.870 ;
        RECT 72.095 178.825 72.385 178.870 ;
        RECT 74.010 178.715 74.150 179.080 ;
        RECT 78.495 179.010 78.785 179.055 ;
        RECT 79.685 179.010 79.975 179.055 ;
        RECT 82.205 179.010 82.495 179.055 ;
        RECT 78.495 178.870 82.495 179.010 ;
        RECT 78.495 178.825 78.785 178.870 ;
        RECT 79.685 178.825 79.975 178.870 ;
        RECT 82.205 178.825 82.495 178.870 ;
        RECT 98.300 178.810 98.620 179.070 ;
        RECT 108.855 179.010 109.145 179.055 ;
        RECT 110.045 179.010 110.335 179.055 ;
        RECT 112.565 179.010 112.855 179.055 ;
        RECT 108.855 178.870 112.855 179.010 ;
        RECT 108.855 178.825 109.145 178.870 ;
        RECT 110.045 178.825 110.335 178.870 ;
        RECT 112.565 178.825 112.855 178.870 ;
        RECT 73.935 178.485 74.225 178.715 ;
        RECT 74.380 178.470 74.700 178.730 ;
        RECT 78.100 178.670 78.390 178.715 ;
        RECT 80.200 178.670 80.490 178.715 ;
        RECT 81.770 178.670 82.060 178.715 ;
        RECT 78.100 178.530 82.060 178.670 ;
        RECT 78.100 178.485 78.390 178.530 ;
        RECT 80.200 178.485 80.490 178.530 ;
        RECT 81.770 178.485 82.060 178.530 ;
        RECT 108.460 178.670 108.750 178.715 ;
        RECT 110.560 178.670 110.850 178.715 ;
        RECT 112.130 178.670 112.420 178.715 ;
        RECT 115.410 178.670 115.550 179.150 ;
        RECT 116.255 178.825 116.545 179.055 ;
        RECT 119.475 179.010 119.765 179.055 ;
        RECT 128.750 179.010 128.890 179.550 ;
        RECT 130.500 179.490 130.820 179.550 ;
        RECT 129.195 179.165 129.485 179.395 ;
        RECT 119.475 178.870 128.890 179.010 ;
        RECT 129.210 179.010 129.350 179.165 ;
        RECT 131.420 179.010 131.740 179.070 ;
        RECT 129.210 178.870 131.740 179.010 ;
        RECT 119.475 178.825 119.765 178.870 ;
        RECT 108.460 178.530 112.420 178.670 ;
        RECT 108.460 178.485 108.750 178.530 ;
        RECT 110.560 178.485 110.850 178.530 ;
        RECT 112.130 178.485 112.420 178.530 ;
        RECT 112.650 178.530 115.550 178.670 ;
        RECT 116.330 178.670 116.470 178.825 ;
        RECT 130.130 178.730 130.270 178.870 ;
        RECT 131.420 178.810 131.740 178.870 ;
        RECT 118.080 178.670 118.400 178.730 ;
        RECT 116.330 178.530 118.400 178.670 ;
        RECT 65.180 178.190 69.090 178.330 ;
        RECT 65.180 178.130 65.500 178.190 ;
        RECT 84.500 178.130 84.820 178.390 ;
        RECT 107.040 178.330 107.360 178.390 ;
        RECT 112.650 178.330 112.790 178.530 ;
        RECT 118.080 178.470 118.400 178.530 ;
        RECT 126.375 178.670 126.665 178.715 ;
        RECT 129.580 178.670 129.900 178.730 ;
        RECT 126.375 178.530 129.900 178.670 ;
        RECT 126.375 178.485 126.665 178.530 ;
        RECT 129.580 178.470 129.900 178.530 ;
        RECT 130.040 178.470 130.360 178.730 ;
        RECT 107.040 178.190 112.790 178.330 ;
        RECT 128.215 178.330 128.505 178.375 ;
        RECT 130.960 178.330 131.280 178.390 ;
        RECT 128.215 178.190 131.280 178.330 ;
        RECT 131.510 178.330 131.650 178.810 ;
        RECT 131.970 178.670 132.110 179.890 ;
        RECT 133.260 179.890 136.325 180.030 ;
        RECT 133.260 179.830 133.580 179.890 ;
        RECT 136.035 179.845 136.325 179.890 ;
        RECT 143.840 179.690 144.160 179.750 ;
        RECT 137.030 179.550 144.160 179.690 ;
        RECT 132.355 179.165 132.645 179.395 ;
        RECT 132.800 179.350 133.120 179.410 ;
        RECT 133.275 179.350 133.565 179.395 ;
        RECT 132.800 179.210 133.565 179.350 ;
        RECT 132.430 179.010 132.570 179.165 ;
        RECT 132.800 179.150 133.120 179.210 ;
        RECT 133.275 179.165 133.565 179.210 ;
        RECT 133.720 179.150 134.040 179.410 ;
        RECT 134.180 179.150 134.500 179.410 ;
        RECT 134.640 179.150 134.960 179.410 ;
        RECT 137.030 179.395 137.170 179.550 ;
        RECT 143.840 179.490 144.160 179.550 ;
        RECT 136.955 179.165 137.245 179.395 ;
        RECT 138.320 179.150 138.640 179.410 ;
        RECT 139.255 179.350 139.545 179.395 ;
        RECT 140.620 179.350 140.940 179.410 ;
        RECT 139.145 179.210 140.940 179.350 ;
        RECT 139.255 179.165 139.545 179.210 ;
        RECT 133.810 179.010 133.950 179.150 ;
        RECT 135.100 179.010 135.420 179.070 ;
        RECT 137.875 179.010 138.165 179.055 ;
        RECT 139.330 179.010 139.470 179.165 ;
        RECT 140.620 179.150 140.940 179.210 ;
        RECT 132.430 178.870 133.030 179.010 ;
        RECT 133.810 178.870 134.825 179.010 ;
        RECT 132.890 178.730 133.030 178.870 ;
        RECT 132.340 178.670 132.660 178.730 ;
        RECT 131.970 178.530 132.660 178.670 ;
        RECT 132.340 178.470 132.660 178.530 ;
        RECT 132.800 178.470 133.120 178.730 ;
        RECT 134.685 178.670 134.825 178.870 ;
        RECT 135.100 178.870 139.470 179.010 ;
        RECT 135.100 178.810 135.420 178.870 ;
        RECT 137.875 178.825 138.165 178.870 ;
        RECT 136.940 178.670 137.260 178.730 ;
        RECT 138.335 178.670 138.625 178.715 ;
        RECT 134.685 178.530 138.625 178.670 ;
        RECT 136.940 178.470 137.260 178.530 ;
        RECT 138.335 178.485 138.625 178.530 ;
        RECT 135.100 178.330 135.420 178.390 ;
        RECT 131.510 178.190 135.420 178.330 ;
        RECT 107.040 178.130 107.360 178.190 ;
        RECT 128.215 178.145 128.505 178.190 ;
        RECT 130.960 178.130 131.280 178.190 ;
        RECT 135.100 178.130 135.420 178.190 ;
        RECT 135.560 178.130 135.880 178.390 ;
        RECT 17.270 177.510 146.990 177.990 ;
        RECT 34.835 177.310 35.125 177.355 ;
        RECT 36.200 177.310 36.520 177.370 ;
        RECT 34.835 177.170 36.520 177.310 ;
        RECT 34.835 177.125 35.125 177.170 ;
        RECT 36.200 177.110 36.520 177.170 ;
        RECT 36.675 177.310 36.965 177.355 ;
        RECT 37.120 177.310 37.440 177.370 ;
        RECT 36.675 177.170 37.440 177.310 ;
        RECT 36.675 177.125 36.965 177.170 ;
        RECT 37.120 177.110 37.440 177.170 ;
        RECT 39.420 177.310 39.740 177.370 ;
        RECT 43.575 177.310 43.865 177.355 ;
        RECT 39.420 177.170 43.865 177.310 ;
        RECT 39.420 177.110 39.740 177.170 ;
        RECT 43.575 177.125 43.865 177.170 ;
        RECT 44.480 177.310 44.800 177.370 ;
        RECT 45.875 177.310 46.165 177.355 ;
        RECT 44.480 177.170 46.165 177.310 ;
        RECT 44.480 177.110 44.800 177.170 ;
        RECT 45.875 177.125 46.165 177.170 ;
        RECT 47.255 177.310 47.545 177.355 ;
        RECT 47.700 177.310 48.020 177.370 ;
        RECT 47.255 177.170 48.020 177.310 ;
        RECT 47.255 177.125 47.545 177.170 ;
        RECT 47.700 177.110 48.020 177.170 ;
        RECT 48.175 177.310 48.465 177.355 ;
        RECT 48.620 177.310 48.940 177.370 ;
        RECT 48.175 177.170 48.940 177.310 ;
        RECT 48.175 177.125 48.465 177.170 ;
        RECT 48.620 177.110 48.940 177.170 ;
        RECT 65.640 177.110 65.960 177.370 ;
        RECT 95.080 177.310 95.400 177.370 ;
        RECT 93.330 177.170 95.400 177.310 ;
        RECT 29.300 176.970 29.620 177.030 ;
        RECT 33.455 176.970 33.745 177.015 ;
        RECT 38.500 176.970 38.820 177.030 ;
        RECT 46.780 176.970 47.100 177.030 ;
        RECT 49.095 176.970 49.385 177.015 ;
        RECT 27.550 176.830 33.210 176.970 ;
        RECT 27.550 176.675 27.690 176.830 ;
        RECT 29.300 176.770 29.620 176.830 ;
        RECT 27.475 176.445 27.765 176.675 ;
        RECT 33.070 176.630 33.210 176.830 ;
        RECT 33.455 176.830 38.820 176.970 ;
        RECT 33.455 176.785 33.745 176.830 ;
        RECT 38.500 176.770 38.820 176.830 ;
        RECT 41.810 176.830 46.090 176.970 ;
        RECT 34.375 176.630 34.665 176.675 ;
        RECT 33.070 176.490 34.665 176.630 ;
        RECT 24.715 176.290 25.005 176.335 ;
        RECT 24.715 176.150 25.850 176.290 ;
        RECT 24.715 176.105 25.005 176.150 ;
        RECT 25.710 175.995 25.850 176.150 ;
        RECT 26.540 176.090 26.860 176.350 ;
        RECT 30.695 176.105 30.985 176.335 ;
        RECT 32.535 176.260 32.825 176.335 ;
        RECT 33.070 176.260 33.210 176.490 ;
        RECT 34.375 176.445 34.665 176.490 ;
        RECT 34.835 176.445 35.125 176.675 ;
        RECT 33.900 176.290 34.220 176.350 ;
        RECT 34.910 176.290 35.050 176.445 ;
        RECT 36.215 176.290 36.505 176.335 ;
        RECT 32.535 176.120 33.210 176.260 ;
        RECT 33.530 176.150 34.220 176.290 ;
        RECT 32.535 176.105 32.825 176.120 ;
        RECT 25.635 175.950 25.925 175.995 ;
        RECT 27.460 175.950 27.780 176.010 ;
        RECT 25.635 175.810 27.780 175.950 ;
        RECT 25.635 175.765 25.925 175.810 ;
        RECT 27.460 175.750 27.780 175.810 ;
        RECT 21.020 175.610 21.340 175.670 ;
        RECT 24.255 175.610 24.545 175.655 ;
        RECT 21.020 175.470 24.545 175.610 ;
        RECT 21.020 175.410 21.340 175.470 ;
        RECT 24.255 175.425 24.545 175.470 ;
        RECT 28.840 175.610 29.160 175.670 ;
        RECT 30.770 175.610 30.910 176.105 ;
        RECT 31.600 175.750 31.920 176.010 ;
        RECT 32.075 175.950 32.365 175.995 ;
        RECT 33.530 175.950 33.670 176.150 ;
        RECT 33.900 176.090 34.220 176.150 ;
        RECT 34.450 176.150 36.505 176.290 ;
        RECT 32.075 175.810 33.670 175.950 ;
        RECT 32.075 175.765 32.365 175.810 ;
        RECT 34.450 175.610 34.590 176.150 ;
        RECT 36.215 176.105 36.505 176.150 ;
        RECT 37.135 176.290 37.425 176.335 ;
        RECT 41.810 176.290 41.950 176.830 ;
        RECT 44.495 176.630 44.785 176.675 ;
        RECT 45.400 176.630 45.720 176.690 ;
        RECT 44.495 176.490 45.720 176.630 ;
        RECT 45.950 176.630 46.090 176.830 ;
        RECT 46.780 176.830 49.385 176.970 ;
        RECT 46.780 176.770 47.100 176.830 ;
        RECT 49.095 176.785 49.385 176.830 ;
        RECT 58.780 176.970 59.070 177.015 ;
        RECT 60.880 176.970 61.170 177.015 ;
        RECT 62.450 176.970 62.740 177.015 ;
        RECT 58.780 176.830 62.740 176.970 ;
        RECT 58.780 176.785 59.070 176.830 ;
        RECT 60.880 176.785 61.170 176.830 ;
        RECT 62.450 176.785 62.740 176.830 ;
        RECT 65.195 176.970 65.485 177.015 ;
        RECT 66.100 176.970 66.420 177.030 ;
        RECT 65.195 176.830 66.420 176.970 ;
        RECT 65.195 176.785 65.485 176.830 ;
        RECT 66.100 176.770 66.420 176.830 ;
        RECT 68.400 176.970 68.690 177.015 ;
        RECT 69.970 176.970 70.260 177.015 ;
        RECT 72.070 176.970 72.360 177.015 ;
        RECT 68.400 176.830 72.360 176.970 ;
        RECT 68.400 176.785 68.690 176.830 ;
        RECT 69.970 176.785 70.260 176.830 ;
        RECT 72.070 176.785 72.360 176.830 ;
        RECT 52.300 176.630 52.620 176.690 ;
        RECT 45.950 176.490 52.620 176.630 ;
        RECT 44.495 176.445 44.785 176.490 ;
        RECT 45.400 176.430 45.720 176.490 ;
        RECT 52.300 176.430 52.620 176.490 ;
        RECT 55.520 176.630 55.840 176.690 ;
        RECT 58.295 176.630 58.585 176.675 ;
        RECT 55.520 176.490 58.585 176.630 ;
        RECT 55.520 176.430 55.840 176.490 ;
        RECT 58.295 176.445 58.585 176.490 ;
        RECT 59.175 176.630 59.465 176.675 ;
        RECT 60.365 176.630 60.655 176.675 ;
        RECT 62.885 176.630 63.175 176.675 ;
        RECT 59.175 176.490 63.175 176.630 ;
        RECT 59.175 176.445 59.465 176.490 ;
        RECT 60.365 176.445 60.655 176.490 ;
        RECT 62.885 176.445 63.175 176.490 ;
        RECT 67.965 176.630 68.255 176.675 ;
        RECT 70.485 176.630 70.775 176.675 ;
        RECT 71.675 176.630 71.965 176.675 ;
        RECT 67.965 176.490 71.965 176.630 ;
        RECT 67.965 176.445 68.255 176.490 ;
        RECT 70.485 176.445 70.775 176.490 ;
        RECT 71.675 176.445 71.965 176.490 ;
        RECT 72.555 176.630 72.845 176.675 ;
        RECT 83.580 176.630 83.900 176.690 ;
        RECT 72.555 176.490 83.900 176.630 ;
        RECT 72.555 176.445 72.845 176.490 ;
        RECT 83.580 176.430 83.900 176.490 ;
        RECT 84.960 176.430 85.280 176.690 ;
        RECT 93.330 176.675 93.470 177.170 ;
        RECT 95.080 177.110 95.400 177.170 ;
        RECT 96.920 177.310 97.240 177.370 ;
        RECT 100.615 177.310 100.905 177.355 ;
        RECT 96.920 177.170 100.905 177.310 ;
        RECT 96.920 177.110 97.240 177.170 ;
        RECT 100.615 177.125 100.905 177.170 ;
        RECT 106.580 177.310 106.900 177.370 ;
        RECT 107.055 177.310 107.345 177.355 ;
        RECT 106.580 177.170 107.345 177.310 ;
        RECT 106.580 177.110 106.900 177.170 ;
        RECT 107.055 177.125 107.345 177.170 ;
        RECT 107.500 177.110 107.820 177.370 ;
        RECT 108.435 177.310 108.725 177.355 ;
        RECT 111.180 177.310 111.500 177.370 ;
        RECT 114.875 177.310 115.165 177.355 ;
        RECT 119.460 177.310 119.780 177.370 ;
        RECT 108.435 177.170 111.500 177.310 ;
        RECT 108.435 177.125 108.725 177.170 ;
        RECT 93.740 176.970 94.030 177.015 ;
        RECT 95.840 176.970 96.130 177.015 ;
        RECT 97.410 176.970 97.700 177.015 ;
        RECT 93.740 176.830 97.700 176.970 ;
        RECT 93.740 176.785 94.030 176.830 ;
        RECT 95.840 176.785 96.130 176.830 ;
        RECT 97.410 176.785 97.700 176.830 ;
        RECT 93.255 176.445 93.545 176.675 ;
        RECT 94.135 176.630 94.425 176.675 ;
        RECT 95.325 176.630 95.615 176.675 ;
        RECT 97.845 176.630 98.135 176.675 ;
        RECT 94.135 176.490 98.135 176.630 ;
        RECT 94.135 176.445 94.425 176.490 ;
        RECT 95.325 176.445 95.615 176.490 ;
        RECT 97.845 176.445 98.135 176.490 ;
        RECT 103.820 176.630 104.140 176.690 ;
        RECT 103.820 176.490 106.810 176.630 ;
        RECT 103.820 176.430 104.140 176.490 ;
        RECT 37.135 176.150 41.950 176.290 ;
        RECT 44.955 176.290 45.245 176.335 ;
        RECT 47.700 176.290 48.020 176.350 ;
        RECT 48.635 176.290 48.925 176.335 ;
        RECT 44.955 176.150 48.925 176.290 ;
        RECT 37.135 176.105 37.425 176.150 ;
        RECT 44.955 176.105 45.245 176.150 ;
        RECT 35.280 175.950 35.600 176.010 ;
        RECT 35.755 175.950 36.045 175.995 ;
        RECT 37.210 175.950 37.350 176.105 ;
        RECT 47.700 176.090 48.020 176.150 ;
        RECT 48.635 176.105 48.925 176.150 ;
        RECT 50.460 176.290 50.780 176.350 ;
        RECT 53.235 176.290 53.525 176.335 ;
        RECT 50.460 176.150 53.525 176.290 ;
        RECT 50.460 176.090 50.780 176.150 ;
        RECT 53.235 176.105 53.525 176.150 ;
        RECT 56.900 176.090 57.220 176.350 ;
        RECT 57.835 176.290 58.125 176.335 ;
        RECT 58.740 176.290 59.060 176.350 ;
        RECT 57.835 176.150 59.060 176.290 ;
        RECT 57.835 176.105 58.125 176.150 ;
        RECT 58.740 176.090 59.060 176.150 ;
        RECT 68.860 176.290 69.180 176.350 ;
        RECT 71.220 176.290 71.510 176.335 ;
        RECT 68.860 176.150 71.510 176.290 ;
        RECT 68.860 176.090 69.180 176.150 ;
        RECT 71.220 176.105 71.510 176.150 ;
        RECT 94.590 176.290 94.880 176.335 ;
        RECT 96.000 176.290 96.320 176.350 ;
        RECT 94.590 176.150 96.320 176.290 ;
        RECT 94.590 176.105 94.880 176.150 ;
        RECT 96.000 176.090 96.320 176.150 ;
        RECT 99.680 176.290 100.000 176.350 ;
        RECT 105.200 176.290 105.520 176.350 ;
        RECT 105.675 176.290 105.965 176.335 ;
        RECT 99.680 176.150 105.965 176.290 ;
        RECT 99.680 176.090 100.000 176.150 ;
        RECT 105.200 176.090 105.520 176.150 ;
        RECT 105.675 176.105 105.965 176.150 ;
        RECT 35.280 175.810 37.350 175.950 ;
        RECT 35.280 175.750 35.600 175.810 ;
        RECT 35.755 175.765 36.045 175.810 ;
        RECT 43.560 175.750 43.880 176.010 ;
        RECT 46.335 175.950 46.625 175.995 ;
        RECT 45.030 175.810 46.625 175.950 ;
        RECT 45.030 175.670 45.170 175.810 ;
        RECT 46.335 175.765 46.625 175.810 ;
        RECT 57.375 175.950 57.665 175.995 ;
        RECT 59.520 175.950 59.810 175.995 ;
        RECT 102.455 175.950 102.745 175.995 ;
        RECT 103.360 175.950 103.680 176.010 ;
        RECT 57.375 175.810 59.810 175.950 ;
        RECT 57.375 175.765 57.665 175.810 ;
        RECT 59.520 175.765 59.810 175.810 ;
        RECT 64.810 175.810 73.920 175.950 ;
        RECT 28.840 175.470 34.590 175.610 ;
        RECT 28.840 175.410 29.160 175.470 ;
        RECT 44.940 175.410 45.260 175.670 ;
        RECT 47.240 175.655 47.560 175.670 ;
        RECT 47.240 175.425 47.625 175.655 ;
        RECT 53.695 175.610 53.985 175.655 ;
        RECT 64.810 175.610 64.950 175.810 ;
        RECT 53.695 175.470 64.950 175.610 ;
        RECT 73.780 175.610 73.920 175.810 ;
        RECT 102.455 175.810 103.680 175.950 ;
        RECT 106.670 175.950 106.810 176.490 ;
        RECT 107.105 176.290 107.395 176.335 ;
        RECT 107.590 176.290 107.730 177.110 ;
        RECT 107.960 176.970 108.280 177.030 ;
        RECT 108.510 176.970 108.650 177.125 ;
        RECT 111.180 177.110 111.500 177.170 ;
        RECT 111.730 177.170 115.165 177.310 ;
        RECT 107.960 176.830 108.650 176.970 ;
        RECT 107.960 176.770 108.280 176.830 ;
        RECT 108.420 176.630 108.740 176.690 ;
        RECT 111.730 176.630 111.870 177.170 ;
        RECT 114.875 177.125 115.165 177.170 ;
        RECT 115.410 177.170 119.780 177.310 ;
        RECT 113.940 176.770 114.260 177.030 ;
        RECT 108.050 176.490 111.870 176.630 ;
        RECT 108.050 176.335 108.190 176.490 ;
        RECT 108.420 176.430 108.740 176.490 ;
        RECT 112.100 176.430 112.420 176.690 ;
        RECT 113.495 176.630 113.785 176.675 ;
        RECT 115.410 176.630 115.550 177.170 ;
        RECT 119.460 177.110 119.780 177.170 ;
        RECT 124.995 177.310 125.285 177.355 ;
        RECT 125.900 177.310 126.220 177.370 ;
        RECT 130.040 177.310 130.360 177.370 ;
        RECT 124.995 177.170 126.220 177.310 ;
        RECT 124.995 177.125 125.285 177.170 ;
        RECT 125.900 177.110 126.220 177.170 ;
        RECT 127.370 177.170 130.360 177.310 ;
        RECT 118.540 176.970 118.860 177.030 ;
        RECT 115.870 176.830 118.860 176.970 ;
        RECT 115.870 176.675 116.010 176.830 ;
        RECT 118.540 176.770 118.860 176.830 ;
        RECT 125.440 176.970 125.760 177.030 ;
        RECT 127.370 176.970 127.510 177.170 ;
        RECT 130.040 177.110 130.360 177.170 ;
        RECT 134.180 177.110 134.500 177.370 ;
        RECT 135.575 177.310 135.865 177.355 ;
        RECT 136.020 177.310 136.340 177.370 ;
        RECT 135.575 177.170 136.340 177.310 ;
        RECT 135.575 177.125 135.865 177.170 ;
        RECT 136.020 177.110 136.340 177.170 ;
        RECT 125.440 176.830 127.510 176.970 ;
        RECT 127.740 176.970 128.060 177.030 ;
        RECT 130.960 176.970 131.280 177.030 ;
        RECT 127.740 176.830 131.280 176.970 ;
        RECT 125.440 176.770 125.760 176.830 ;
        RECT 127.740 176.770 128.060 176.830 ;
        RECT 130.960 176.770 131.280 176.830 ;
        RECT 134.640 176.970 134.960 177.030 ;
        RECT 134.640 176.830 136.250 176.970 ;
        RECT 134.640 176.770 134.960 176.830 ;
        RECT 113.495 176.490 115.550 176.630 ;
        RECT 113.495 176.445 113.785 176.490 ;
        RECT 115.795 176.445 116.085 176.675 ;
        RECT 117.620 176.630 117.940 176.690 ;
        RECT 117.250 176.490 117.940 176.630 ;
        RECT 107.105 176.150 107.730 176.290 ;
        RECT 107.105 176.105 107.395 176.150 ;
        RECT 107.975 176.105 108.265 176.335 ;
        RECT 114.860 176.090 115.180 176.350 ;
        RECT 117.250 176.335 117.390 176.490 ;
        RECT 117.620 176.430 117.940 176.490 ;
        RECT 124.060 176.430 124.380 176.690 ;
        RECT 129.690 176.630 129.980 176.675 ;
        RECT 134.195 176.630 134.485 176.675 ;
        RECT 135.560 176.630 135.880 176.690 ;
        RECT 129.690 176.490 133.950 176.630 ;
        RECT 129.690 176.445 129.980 176.490 ;
        RECT 117.175 176.105 117.465 176.335 ;
        RECT 118.540 176.090 118.860 176.350 ;
        RECT 119.000 176.290 119.320 176.350 ;
        RECT 119.935 176.290 120.225 176.335 ;
        RECT 119.000 176.150 120.225 176.290 ;
        RECT 119.000 176.090 119.320 176.150 ;
        RECT 119.935 176.105 120.225 176.150 ;
        RECT 120.855 176.105 121.145 176.335 ;
        RECT 110.720 175.950 111.040 176.010 ;
        RECT 116.240 175.950 116.560 176.010 ;
        RECT 106.670 175.810 116.560 175.950 ;
        RECT 118.630 175.950 118.770 176.090 ;
        RECT 120.930 175.950 121.070 176.105 ;
        RECT 125.440 176.090 125.760 176.350 ;
        RECT 127.740 176.290 128.060 176.350 ;
        RECT 128.675 176.290 128.965 176.335 ;
        RECT 130.515 176.290 130.805 176.335 ;
        RECT 131.420 176.290 131.740 176.350 ;
        RECT 133.810 176.335 133.950 176.490 ;
        RECT 134.195 176.490 135.880 176.630 ;
        RECT 134.195 176.445 134.485 176.490 ;
        RECT 135.560 176.430 135.880 176.490 ;
        RECT 136.110 176.335 136.250 176.830 ;
        RECT 127.740 176.150 128.965 176.290 ;
        RECT 127.740 176.090 128.060 176.150 ;
        RECT 128.675 176.105 128.965 176.150 ;
        RECT 130.130 176.150 130.805 176.290 ;
        RECT 130.130 176.010 130.270 176.150 ;
        RECT 130.515 176.105 130.805 176.150 ;
        RECT 131.050 176.150 131.740 176.290 ;
        RECT 118.630 175.810 121.070 175.950 ;
        RECT 121.760 175.950 122.080 176.010 ;
        RECT 125.915 175.950 126.205 175.995 ;
        RECT 126.820 175.950 127.140 176.010 ;
        RECT 129.135 175.950 129.425 175.995 ;
        RECT 121.760 175.810 129.425 175.950 ;
        RECT 102.455 175.765 102.745 175.810 ;
        RECT 103.360 175.750 103.680 175.810 ;
        RECT 110.720 175.750 111.040 175.810 ;
        RECT 116.240 175.750 116.560 175.810 ;
        RECT 121.760 175.750 122.080 175.810 ;
        RECT 125.915 175.765 126.205 175.810 ;
        RECT 126.820 175.750 127.140 175.810 ;
        RECT 129.135 175.765 129.425 175.810 ;
        RECT 130.040 175.750 130.360 176.010 ;
        RECT 131.050 175.950 131.190 176.150 ;
        RECT 131.420 176.090 131.740 176.150 ;
        RECT 133.735 176.105 134.025 176.335 ;
        RECT 136.035 176.105 136.325 176.335 ;
        RECT 136.940 176.090 137.260 176.350 ;
        RECT 145.220 176.090 145.540 176.350 ;
        RECT 130.590 175.810 131.190 175.950 ;
        RECT 132.800 175.950 133.120 176.010 ;
        RECT 132.800 175.810 144.530 175.950 ;
        RECT 78.060 175.610 78.380 175.670 ;
        RECT 73.780 175.470 78.380 175.610 ;
        RECT 53.695 175.425 53.985 175.470 ;
        RECT 47.240 175.410 47.560 175.425 ;
        RECT 78.060 175.410 78.380 175.470 ;
        RECT 87.260 175.610 87.580 175.670 ;
        RECT 87.735 175.610 88.025 175.655 ;
        RECT 87.260 175.470 88.025 175.610 ;
        RECT 87.260 175.410 87.580 175.470 ;
        RECT 87.735 175.425 88.025 175.470 ;
        RECT 100.155 175.610 100.445 175.655 ;
        RECT 102.915 175.610 103.205 175.655 ;
        RECT 104.280 175.610 104.600 175.670 ;
        RECT 100.155 175.470 104.600 175.610 ;
        RECT 100.155 175.425 100.445 175.470 ;
        RECT 102.915 175.425 103.205 175.470 ;
        RECT 104.280 175.410 104.600 175.470 ;
        RECT 106.135 175.610 106.425 175.655 ;
        RECT 107.500 175.610 107.820 175.670 ;
        RECT 106.135 175.470 107.820 175.610 ;
        RECT 106.135 175.425 106.425 175.470 ;
        RECT 107.500 175.410 107.820 175.470 ;
        RECT 114.400 175.610 114.720 175.670 ;
        RECT 120.395 175.610 120.685 175.655 ;
        RECT 114.400 175.470 120.685 175.610 ;
        RECT 114.400 175.410 114.720 175.470 ;
        RECT 120.395 175.425 120.685 175.470 ;
        RECT 122.680 175.410 123.000 175.670 ;
        RECT 124.520 175.610 124.840 175.670 ;
        RECT 128.200 175.610 128.520 175.670 ;
        RECT 124.520 175.470 128.520 175.610 ;
        RECT 124.520 175.410 124.840 175.470 ;
        RECT 128.200 175.410 128.520 175.470 ;
        RECT 128.660 175.610 128.980 175.670 ;
        RECT 130.590 175.610 130.730 175.810 ;
        RECT 132.800 175.750 133.120 175.810 ;
        RECT 128.660 175.470 130.730 175.610 ;
        RECT 130.975 175.610 131.265 175.655 ;
        RECT 133.720 175.610 134.040 175.670 ;
        RECT 130.975 175.470 134.040 175.610 ;
        RECT 128.660 175.410 128.980 175.470 ;
        RECT 130.975 175.425 131.265 175.470 ;
        RECT 133.720 175.410 134.040 175.470 ;
        RECT 134.180 175.610 134.500 175.670 ;
        RECT 144.390 175.655 144.530 175.810 ;
        RECT 136.035 175.610 136.325 175.655 ;
        RECT 134.180 175.470 136.325 175.610 ;
        RECT 134.180 175.410 134.500 175.470 ;
        RECT 136.035 175.425 136.325 175.470 ;
        RECT 144.315 175.425 144.605 175.655 ;
        RECT 17.270 174.790 146.990 175.270 ;
        RECT 150.360 174.810 151.020 174.990 ;
        RECT 23.715 174.590 24.005 174.635 ;
        RECT 25.175 174.590 25.465 174.635 ;
        RECT 23.715 174.450 25.465 174.590 ;
        RECT 23.715 174.405 24.005 174.450 ;
        RECT 25.175 174.405 25.465 174.450 ;
        RECT 33.900 174.590 34.220 174.650 ;
        RECT 35.740 174.590 36.060 174.650 ;
        RECT 41.720 174.590 42.040 174.650 ;
        RECT 33.900 174.450 42.040 174.590 ;
        RECT 33.900 174.390 34.220 174.450 ;
        RECT 35.740 174.390 36.060 174.450 ;
        RECT 41.720 174.390 42.040 174.450 ;
        RECT 43.560 174.390 43.880 174.650 ;
        RECT 45.400 174.390 45.720 174.650 ;
        RECT 65.180 174.590 65.500 174.650 ;
        RECT 68.415 174.590 68.705 174.635 ;
        RECT 65.180 174.450 68.705 174.590 ;
        RECT 65.180 174.390 65.500 174.450 ;
        RECT 68.415 174.405 68.705 174.450 ;
        RECT 84.055 174.405 84.345 174.635 ;
        RECT 100.140 174.590 100.460 174.650 ;
        RECT 105.200 174.590 105.520 174.650 ;
        RECT 114.415 174.590 114.705 174.635 ;
        RECT 123.600 174.590 123.920 174.650 ;
        RECT 126.360 174.590 126.680 174.650 ;
        RECT 100.140 174.450 104.970 174.590 ;
        RECT 21.940 174.250 22.260 174.310 ;
        RECT 24.715 174.250 25.005 174.295 ;
        RECT 26.540 174.250 26.860 174.310 ;
        RECT 38.515 174.250 38.805 174.295 ;
        RECT 21.940 174.110 25.005 174.250 ;
        RECT 21.940 174.050 22.260 174.110 ;
        RECT 24.715 174.065 25.005 174.110 ;
        RECT 25.480 174.110 29.990 174.250 ;
        RECT 21.495 173.910 21.785 173.955 ;
        RECT 22.415 173.910 22.705 173.955 ;
        RECT 25.480 173.910 25.620 174.110 ;
        RECT 26.540 174.050 26.860 174.110 ;
        RECT 21.495 173.770 22.170 173.910 ;
        RECT 21.495 173.725 21.785 173.770 ;
        RECT 22.030 173.230 22.170 173.770 ;
        RECT 22.415 173.770 25.620 173.910 ;
        RECT 22.415 173.725 22.705 173.770 ;
        RECT 26.095 173.725 26.385 173.955 ;
        RECT 27.015 173.910 27.305 173.955 ;
        RECT 27.460 173.910 27.780 173.970 ;
        RECT 28.840 173.910 29.160 173.970 ;
        RECT 27.015 173.770 27.780 173.910 ;
        RECT 27.015 173.725 27.305 173.770 ;
        RECT 26.170 173.570 26.310 173.725 ;
        RECT 27.460 173.710 27.780 173.770 ;
        RECT 28.010 173.770 29.160 173.910 ;
        RECT 28.010 173.570 28.150 173.770 ;
        RECT 28.840 173.710 29.160 173.770 ;
        RECT 29.300 173.710 29.620 173.970 ;
        RECT 29.850 173.955 29.990 174.110 ;
        RECT 32.150 174.110 38.805 174.250 ;
        RECT 32.150 173.970 32.290 174.110 ;
        RECT 38.515 174.065 38.805 174.110 ;
        RECT 42.195 174.250 42.485 174.295 ;
        RECT 45.490 174.250 45.630 174.390 ;
        RECT 42.195 174.110 45.630 174.250 ;
        RECT 58.280 174.250 58.600 174.310 ;
        RECT 62.740 174.250 63.030 174.295 ;
        RECT 58.280 174.110 63.030 174.250 ;
        RECT 42.195 174.065 42.485 174.110 ;
        RECT 58.280 174.050 58.600 174.110 ;
        RECT 62.740 174.065 63.030 174.110 ;
        RECT 82.370 174.250 82.660 174.295 ;
        RECT 84.130 174.250 84.270 174.405 ;
        RECT 100.140 174.390 100.460 174.450 ;
        RECT 82.370 174.110 84.270 174.250 ;
        RECT 86.815 174.250 87.105 174.295 ;
        RECT 87.260 174.250 87.580 174.310 ;
        RECT 86.815 174.110 87.580 174.250 ;
        RECT 82.370 174.065 82.660 174.110 ;
        RECT 86.815 174.065 87.105 174.110 ;
        RECT 87.260 174.050 87.580 174.110 ;
        RECT 87.720 174.050 88.040 174.310 ;
        RECT 90.495 174.250 90.785 174.295 ;
        RECT 90.940 174.250 91.260 174.310 ;
        RECT 103.820 174.250 104.140 174.310 ;
        RECT 90.495 174.110 104.140 174.250 ;
        RECT 90.495 174.065 90.785 174.110 ;
        RECT 90.940 174.050 91.260 174.110 ;
        RECT 103.820 174.050 104.140 174.110 ;
        RECT 29.775 173.725 30.065 173.955 ;
        RECT 32.060 173.710 32.380 173.970 ;
        RECT 37.595 173.910 37.885 173.955 ;
        RECT 39.420 173.910 39.740 173.970 ;
        RECT 37.595 173.770 39.740 173.910 ;
        RECT 37.595 173.725 37.885 173.770 ;
        RECT 39.420 173.710 39.740 173.770 ;
        RECT 39.895 173.910 40.185 173.955 ;
        RECT 40.340 173.910 40.660 173.970 ;
        RECT 39.895 173.770 41.490 173.910 ;
        RECT 39.895 173.725 40.185 173.770 ;
        RECT 40.340 173.710 40.660 173.770 ;
        RECT 26.170 173.430 28.150 173.570 ;
        RECT 28.380 173.370 28.700 173.630 ;
        RECT 26.080 173.230 26.400 173.290 ;
        RECT 29.390 173.230 29.530 173.710 ;
        RECT 31.600 173.570 31.920 173.630 ;
        RECT 35.280 173.570 35.600 173.630 ;
        RECT 31.600 173.430 35.600 173.570 ;
        RECT 31.600 173.370 31.920 173.430 ;
        RECT 35.280 173.370 35.600 173.430 ;
        RECT 22.030 173.090 29.530 173.230 ;
        RECT 34.820 173.230 35.140 173.290 ;
        RECT 41.350 173.230 41.490 173.770 ;
        RECT 41.735 173.725 42.025 173.955 ;
        RECT 42.655 173.910 42.945 173.955 ;
        RECT 44.020 173.910 44.340 173.970 ;
        RECT 44.495 173.910 44.785 173.955 ;
        RECT 42.655 173.770 44.785 173.910 ;
        RECT 42.655 173.725 42.945 173.770 ;
        RECT 41.810 173.570 41.950 173.725 ;
        RECT 44.020 173.710 44.340 173.770 ;
        RECT 44.495 173.725 44.785 173.770 ;
        RECT 44.940 173.710 45.260 173.970 ;
        RECT 45.415 173.910 45.705 173.955 ;
        RECT 45.860 173.910 46.180 173.970 ;
        RECT 45.415 173.770 46.180 173.910 ;
        RECT 45.415 173.725 45.705 173.770 ;
        RECT 45.860 173.710 46.180 173.770 ;
        RECT 46.320 173.710 46.640 173.970 ;
        RECT 46.795 173.725 47.085 173.955 ;
        RECT 47.240 173.910 47.560 173.970 ;
        RECT 54.140 173.955 54.460 173.970 ;
        RECT 47.715 173.910 48.005 173.955 ;
        RECT 47.240 173.770 48.005 173.910 ;
        RECT 43.100 173.570 43.420 173.630 ;
        RECT 45.030 173.570 45.170 173.710 ;
        RECT 46.870 173.570 47.010 173.725 ;
        RECT 47.240 173.710 47.560 173.770 ;
        RECT 47.715 173.725 48.005 173.770 ;
        RECT 54.140 173.725 54.490 173.955 ;
        RECT 83.120 173.910 83.440 173.970 ;
        RECT 84.975 173.910 85.265 173.955 ;
        RECT 83.120 173.770 85.265 173.910 ;
        RECT 54.140 173.710 54.460 173.725 ;
        RECT 83.120 173.710 83.440 173.770 ;
        RECT 84.975 173.725 85.265 173.770 ;
        RECT 85.435 173.725 85.725 173.955 ;
        RECT 88.180 173.910 88.500 173.970 ;
        RECT 88.655 173.910 88.945 173.955 ;
        RECT 88.180 173.770 88.945 173.910 ;
        RECT 41.810 173.430 47.010 173.570 ;
        RECT 43.100 173.370 43.420 173.430 ;
        RECT 47.330 173.230 47.470 173.710 ;
        RECT 50.945 173.570 51.235 173.615 ;
        RECT 53.465 173.570 53.755 173.615 ;
        RECT 54.655 173.570 54.945 173.615 ;
        RECT 50.945 173.430 54.945 173.570 ;
        RECT 50.945 173.385 51.235 173.430 ;
        RECT 53.465 173.385 53.755 173.430 ;
        RECT 54.655 173.385 54.945 173.430 ;
        RECT 55.520 173.570 55.840 173.630 ;
        RECT 61.515 173.570 61.805 173.615 ;
        RECT 55.520 173.430 61.805 173.570 ;
        RECT 55.520 173.370 55.840 173.430 ;
        RECT 61.515 173.385 61.805 173.430 ;
        RECT 62.395 173.570 62.685 173.615 ;
        RECT 63.585 173.570 63.875 173.615 ;
        RECT 66.105 173.570 66.395 173.615 ;
        RECT 62.395 173.430 66.395 173.570 ;
        RECT 62.395 173.385 62.685 173.430 ;
        RECT 63.585 173.385 63.875 173.430 ;
        RECT 66.105 173.385 66.395 173.430 ;
        RECT 79.005 173.570 79.295 173.615 ;
        RECT 81.525 173.570 81.815 173.615 ;
        RECT 82.715 173.570 83.005 173.615 ;
        RECT 79.005 173.430 83.005 173.570 ;
        RECT 79.005 173.385 79.295 173.430 ;
        RECT 81.525 173.385 81.815 173.430 ;
        RECT 82.715 173.385 83.005 173.430 ;
        RECT 83.580 173.370 83.900 173.630 ;
        RECT 34.820 173.090 41.030 173.230 ;
        RECT 41.350 173.090 47.470 173.230 ;
        RECT 51.380 173.230 51.670 173.275 ;
        RECT 52.950 173.230 53.240 173.275 ;
        RECT 55.050 173.230 55.340 173.275 ;
        RECT 51.380 173.090 55.340 173.230 ;
        RECT 26.080 173.030 26.400 173.090 ;
        RECT 34.820 173.030 35.140 173.090 ;
        RECT 20.575 172.890 20.865 172.935 ;
        RECT 21.480 172.890 21.800 172.950 ;
        RECT 20.575 172.750 21.800 172.890 ;
        RECT 20.575 172.705 20.865 172.750 ;
        RECT 21.480 172.690 21.800 172.750 ;
        RECT 22.875 172.890 23.165 172.935 ;
        RECT 23.320 172.890 23.640 172.950 ;
        RECT 22.875 172.750 23.640 172.890 ;
        RECT 22.875 172.705 23.165 172.750 ;
        RECT 23.320 172.690 23.640 172.750 ;
        RECT 23.795 172.890 24.085 172.935 ;
        RECT 27.000 172.890 27.320 172.950 ;
        RECT 23.795 172.750 27.320 172.890 ;
        RECT 23.795 172.705 24.085 172.750 ;
        RECT 27.000 172.690 27.320 172.750 ;
        RECT 30.680 172.690 31.000 172.950 ;
        RECT 31.600 172.690 31.920 172.950 ;
        RECT 36.675 172.890 36.965 172.935 ;
        RECT 38.040 172.890 38.360 172.950 ;
        RECT 36.675 172.750 38.360 172.890 ;
        RECT 36.675 172.705 36.965 172.750 ;
        RECT 38.040 172.690 38.360 172.750 ;
        RECT 39.420 172.690 39.740 172.950 ;
        RECT 40.890 172.890 41.030 173.090 ;
        RECT 51.380 173.045 51.670 173.090 ;
        RECT 52.950 173.045 53.240 173.090 ;
        RECT 55.050 173.045 55.340 173.090 ;
        RECT 62.000 173.230 62.290 173.275 ;
        RECT 64.100 173.230 64.390 173.275 ;
        RECT 65.670 173.230 65.960 173.275 ;
        RECT 62.000 173.090 65.960 173.230 ;
        RECT 62.000 173.045 62.290 173.090 ;
        RECT 64.100 173.045 64.390 173.090 ;
        RECT 65.670 173.045 65.960 173.090 ;
        RECT 79.440 173.230 79.730 173.275 ;
        RECT 81.010 173.230 81.300 173.275 ;
        RECT 83.110 173.230 83.400 173.275 ;
        RECT 79.440 173.090 83.400 173.230 ;
        RECT 85.510 173.230 85.650 173.725 ;
        RECT 88.180 173.710 88.500 173.770 ;
        RECT 88.655 173.725 88.945 173.770 ;
        RECT 98.760 173.710 99.080 173.970 ;
        RECT 99.680 173.710 100.000 173.970 ;
        RECT 104.830 173.910 104.970 174.450 ;
        RECT 105.200 174.450 105.890 174.590 ;
        RECT 105.200 174.390 105.520 174.450 ;
        RECT 105.750 174.295 105.890 174.450 ;
        RECT 114.415 174.450 126.680 174.590 ;
        RECT 114.415 174.405 114.705 174.450 ;
        RECT 123.600 174.390 123.920 174.450 ;
        RECT 126.360 174.390 126.680 174.450 ;
        RECT 130.590 174.450 135.790 174.590 ;
        RECT 130.590 174.310 130.730 174.450 ;
        RECT 105.720 174.065 106.010 174.295 ;
        RECT 108.420 174.250 108.740 174.310 ;
        RECT 106.715 174.110 110.950 174.250 ;
        RECT 106.715 173.910 106.855 174.110 ;
        RECT 108.420 174.050 108.740 174.110 ;
        RECT 104.830 173.770 106.855 173.910 ;
        RECT 107.055 173.910 107.345 173.955 ;
        RECT 107.960 173.910 108.280 173.970 ;
        RECT 110.810 173.955 110.950 174.110 ;
        RECT 111.180 174.050 111.500 174.310 ;
        RECT 114.875 174.250 115.165 174.295 ;
        RECT 115.320 174.250 115.640 174.310 ;
        RECT 117.620 174.250 117.940 174.310 ;
        RECT 121.760 174.295 122.080 174.310 ;
        RECT 114.875 174.110 117.940 174.250 ;
        RECT 114.875 174.065 115.165 174.110 ;
        RECT 115.320 174.050 115.640 174.110 ;
        RECT 117.620 174.050 117.940 174.110 ;
        RECT 121.695 174.065 122.080 174.295 ;
        RECT 122.695 174.250 122.985 174.295 ;
        RECT 125.440 174.250 125.760 174.310 ;
        RECT 122.695 174.110 125.760 174.250 ;
        RECT 122.695 174.065 122.985 174.110 ;
        RECT 121.760 174.050 122.080 174.065 ;
        RECT 125.440 174.050 125.760 174.110 ;
        RECT 127.280 174.050 127.600 174.310 ;
        RECT 130.500 174.250 130.820 174.310 ;
        RECT 135.650 174.295 135.790 174.450 ;
        RECT 150.360 174.575 152.045 174.810 ;
        RECT 150.360 174.390 151.020 174.575 ;
        RECT 130.130 174.110 130.820 174.250 ;
        RECT 110.735 173.910 111.025 173.955 ;
        RECT 107.055 173.770 108.280 173.910 ;
        RECT 107.055 173.725 107.345 173.770 ;
        RECT 107.960 173.710 108.280 173.770 ;
        RECT 109.890 173.770 111.025 173.910 ;
        RECT 111.270 173.910 111.410 174.050 ;
        RECT 113.020 173.910 113.340 173.970 ;
        RECT 117.175 173.910 117.465 173.955 ;
        RECT 111.270 173.770 113.340 173.910 ;
        RECT 85.880 173.570 86.200 173.630 ;
        RECT 87.275 173.570 87.565 173.615 ;
        RECT 85.880 173.430 87.565 173.570 ;
        RECT 85.880 173.370 86.200 173.430 ;
        RECT 87.275 173.385 87.565 173.430 ;
        RECT 102.465 173.570 102.755 173.615 ;
        RECT 104.985 173.570 105.275 173.615 ;
        RECT 106.175 173.570 106.465 173.615 ;
        RECT 102.465 173.430 106.465 173.570 ;
        RECT 102.465 173.385 102.755 173.430 ;
        RECT 104.985 173.385 105.275 173.430 ;
        RECT 106.175 173.385 106.465 173.430 ;
        RECT 88.640 173.230 88.960 173.290 ;
        RECT 85.510 173.090 88.960 173.230 ;
        RECT 79.440 173.045 79.730 173.090 ;
        RECT 81.010 173.045 81.300 173.090 ;
        RECT 83.110 173.045 83.400 173.090 ;
        RECT 88.640 173.030 88.960 173.090 ;
        RECT 99.235 173.230 99.525 173.275 ;
        RECT 102.900 173.230 103.190 173.275 ;
        RECT 104.470 173.230 104.760 173.275 ;
        RECT 106.570 173.230 106.860 173.275 ;
        RECT 99.235 173.090 102.670 173.230 ;
        RECT 99.235 173.045 99.525 173.090 ;
        RECT 46.320 172.890 46.640 172.950 ;
        RECT 40.890 172.750 46.640 172.890 ;
        RECT 46.320 172.690 46.640 172.750 ;
        RECT 47.240 172.690 47.560 172.950 ;
        RECT 47.700 172.890 48.020 172.950 ;
        RECT 48.635 172.890 48.925 172.935 ;
        RECT 47.700 172.750 48.925 172.890 ;
        RECT 47.700 172.690 48.020 172.750 ;
        RECT 48.635 172.705 48.925 172.750 ;
        RECT 76.695 172.890 76.985 172.935 ;
        RECT 84.960 172.890 85.280 172.950 ;
        RECT 76.695 172.750 85.280 172.890 ;
        RECT 102.530 172.890 102.670 173.090 ;
        RECT 102.900 173.090 106.860 173.230 ;
        RECT 102.900 173.045 103.190 173.090 ;
        RECT 104.470 173.045 104.760 173.090 ;
        RECT 106.570 173.045 106.860 173.090 ;
        RECT 106.120 172.890 106.440 172.950 ;
        RECT 102.530 172.750 106.440 172.890 ;
        RECT 76.695 172.705 76.985 172.750 ;
        RECT 84.960 172.690 85.280 172.750 ;
        RECT 106.120 172.690 106.440 172.750 ;
        RECT 107.515 172.890 107.805 172.935 ;
        RECT 108.420 172.890 108.740 172.950 ;
        RECT 107.515 172.750 108.740 172.890 ;
        RECT 109.890 172.890 110.030 173.770 ;
        RECT 110.735 173.725 111.025 173.770 ;
        RECT 113.020 173.710 113.340 173.770 ;
        RECT 114.950 173.770 117.465 173.910 ;
        RECT 114.950 173.630 115.090 173.770 ;
        RECT 117.175 173.725 117.465 173.770 ;
        RECT 123.140 173.710 123.460 173.970 ;
        RECT 129.120 173.710 129.440 173.970 ;
        RECT 130.130 173.955 130.270 174.110 ;
        RECT 130.500 174.050 130.820 174.110 ;
        RECT 135.575 174.065 135.865 174.295 ;
        RECT 137.400 174.250 137.720 174.310 ;
        RECT 136.570 174.110 137.720 174.250 ;
        RECT 130.055 173.725 130.345 173.955 ;
        RECT 130.960 173.710 131.280 173.970 ;
        RECT 131.950 173.725 132.240 173.955 ;
        RECT 134.655 173.910 134.945 173.955 ;
        RECT 135.100 173.910 135.420 173.970 ;
        RECT 136.570 173.955 136.710 174.110 ;
        RECT 137.400 174.050 137.720 174.110 ;
        RECT 137.860 173.955 138.180 173.970 ;
        RECT 134.655 173.770 135.420 173.910 ;
        RECT 134.655 173.725 134.945 173.770 ;
        RECT 110.260 173.570 110.580 173.630 ;
        RECT 111.195 173.570 111.485 173.615 ;
        RECT 110.260 173.430 111.485 173.570 ;
        RECT 110.260 173.370 110.580 173.430 ;
        RECT 111.195 173.385 111.485 173.430 ;
        RECT 112.560 173.570 112.880 173.630 ;
        RECT 113.495 173.570 113.785 173.615 ;
        RECT 112.560 173.430 113.785 173.570 ;
        RECT 112.560 173.370 112.880 173.430 ;
        RECT 113.495 173.385 113.785 173.430 ;
        RECT 114.860 173.370 115.180 173.630 ;
        RECT 116.715 173.570 117.005 173.615 ;
        RECT 117.620 173.570 117.940 173.630 ;
        RECT 125.900 173.570 126.220 173.630 ;
        RECT 130.515 173.570 130.805 173.615 ;
        RECT 116.715 173.430 126.220 173.570 ;
        RECT 116.715 173.385 117.005 173.430 ;
        RECT 117.620 173.370 117.940 173.430 ;
        RECT 120.930 173.275 121.070 173.430 ;
        RECT 125.900 173.370 126.220 173.430 ;
        RECT 130.130 173.430 130.805 173.570 ;
        RECT 130.130 173.290 130.270 173.430 ;
        RECT 130.515 173.385 130.805 173.430 ;
        RECT 120.855 173.045 121.145 173.275 ;
        RECT 130.040 173.030 130.360 173.290 ;
        RECT 131.970 173.230 132.110 173.725 ;
        RECT 135.100 173.710 135.420 173.770 ;
        RECT 136.495 173.725 136.785 173.955 ;
        RECT 137.830 173.725 138.180 173.955 ;
        RECT 137.860 173.710 138.180 173.725 ;
        RECT 143.840 173.710 144.160 173.970 ;
        RECT 137.375 173.570 137.665 173.615 ;
        RECT 138.565 173.570 138.855 173.615 ;
        RECT 141.085 173.570 141.375 173.615 ;
        RECT 137.375 173.430 141.375 173.570 ;
        RECT 137.375 173.385 137.665 173.430 ;
        RECT 138.565 173.385 138.855 173.430 ;
        RECT 141.085 173.385 141.375 173.430 ;
        RECT 131.510 173.090 132.110 173.230 ;
        RECT 132.815 173.230 133.105 173.275 ;
        RECT 136.480 173.230 136.800 173.290 ;
        RECT 132.815 173.090 136.800 173.230 ;
        RECT 115.335 172.890 115.625 172.935 ;
        RECT 109.890 172.750 115.625 172.890 ;
        RECT 107.515 172.705 107.805 172.750 ;
        RECT 108.420 172.690 108.740 172.750 ;
        RECT 115.335 172.705 115.625 172.750 ;
        RECT 118.080 172.690 118.400 172.950 ;
        RECT 121.775 172.890 122.065 172.935 ;
        RECT 124.060 172.890 124.380 172.950 ;
        RECT 121.775 172.750 124.380 172.890 ;
        RECT 121.775 172.705 122.065 172.750 ;
        RECT 124.060 172.690 124.380 172.750 ;
        RECT 128.660 172.890 128.980 172.950 ;
        RECT 131.510 172.890 131.650 173.090 ;
        RECT 132.815 173.045 133.105 173.090 ;
        RECT 136.480 173.030 136.800 173.090 ;
        RECT 136.980 173.230 137.270 173.275 ;
        RECT 139.080 173.230 139.370 173.275 ;
        RECT 140.650 173.230 140.940 173.275 ;
        RECT 136.980 173.090 140.940 173.230 ;
        RECT 136.980 173.045 137.270 173.090 ;
        RECT 139.080 173.045 139.370 173.090 ;
        RECT 140.650 173.045 140.940 173.090 ;
        RECT 128.660 172.750 131.650 172.890 ;
        RECT 131.880 172.890 132.200 172.950 ;
        RECT 133.735 172.890 134.025 172.935 ;
        RECT 131.880 172.750 134.025 172.890 ;
        RECT 128.660 172.690 128.980 172.750 ;
        RECT 131.880 172.690 132.200 172.750 ;
        RECT 133.735 172.705 134.025 172.750 ;
        RECT 143.380 172.690 143.700 172.950 ;
        RECT 144.760 172.690 145.080 172.950 ;
        RECT 17.270 172.070 146.990 172.550 ;
        RECT 26.080 171.670 26.400 171.930 ;
        RECT 27.000 171.670 27.320 171.930 ;
        RECT 28.840 171.670 29.160 171.930 ;
        RECT 29.775 171.870 30.065 171.915 ;
        RECT 32.060 171.870 32.380 171.930 ;
        RECT 39.895 171.870 40.185 171.915 ;
        RECT 40.340 171.870 40.660 171.930 ;
        RECT 29.775 171.730 39.190 171.870 ;
        RECT 29.775 171.685 30.065 171.730 ;
        RECT 32.060 171.670 32.380 171.730 ;
        RECT 19.680 171.530 19.970 171.575 ;
        RECT 21.780 171.530 22.070 171.575 ;
        RECT 23.350 171.530 23.640 171.575 ;
        RECT 19.680 171.390 23.640 171.530 ;
        RECT 19.680 171.345 19.970 171.390 ;
        RECT 21.780 171.345 22.070 171.390 ;
        RECT 23.350 171.345 23.640 171.390 ;
        RECT 20.075 171.190 20.365 171.235 ;
        RECT 21.265 171.190 21.555 171.235 ;
        RECT 23.785 171.190 24.075 171.235 ;
        RECT 28.930 171.190 29.070 171.670 ;
        RECT 31.180 171.530 31.470 171.575 ;
        RECT 33.280 171.530 33.570 171.575 ;
        RECT 34.850 171.530 35.140 171.575 ;
        RECT 31.180 171.390 35.140 171.530 ;
        RECT 31.180 171.345 31.470 171.390 ;
        RECT 33.280 171.345 33.570 171.390 ;
        RECT 34.850 171.345 35.140 171.390 ;
        RECT 20.075 171.050 24.075 171.190 ;
        RECT 20.075 171.005 20.365 171.050 ;
        RECT 21.265 171.005 21.555 171.050 ;
        RECT 23.785 171.005 24.075 171.050 ;
        RECT 26.630 171.050 29.070 171.190 ;
        RECT 31.575 171.190 31.865 171.235 ;
        RECT 32.765 171.190 33.055 171.235 ;
        RECT 35.285 171.190 35.575 171.235 ;
        RECT 31.575 171.050 35.575 171.190 ;
        RECT 19.180 170.650 19.500 170.910 ;
        RECT 26.630 170.895 26.770 171.050 ;
        RECT 31.575 171.005 31.865 171.050 ;
        RECT 32.765 171.005 33.055 171.050 ;
        RECT 35.285 171.005 35.575 171.050 ;
        RECT 26.555 170.665 26.845 170.895 ;
        RECT 27.460 170.850 27.780 170.910 ;
        RECT 30.220 170.850 30.540 170.910 ;
        RECT 39.050 170.895 39.190 171.730 ;
        RECT 39.895 171.730 40.660 171.870 ;
        RECT 39.895 171.685 40.185 171.730 ;
        RECT 40.340 171.670 40.660 171.730 ;
        RECT 45.415 171.870 45.705 171.915 ;
        RECT 47.240 171.870 47.560 171.930 ;
        RECT 45.415 171.730 47.560 171.870 ;
        RECT 45.415 171.685 45.705 171.730 ;
        RECT 47.240 171.670 47.560 171.730 ;
        RECT 51.855 171.870 52.145 171.915 ;
        RECT 54.140 171.870 54.460 171.930 ;
        RECT 51.855 171.730 54.460 171.870 ;
        RECT 51.855 171.685 52.145 171.730 ;
        RECT 54.140 171.670 54.460 171.730 ;
        RECT 84.500 171.870 84.820 171.930 ;
        RECT 87.275 171.870 87.565 171.915 ;
        RECT 84.500 171.730 87.565 171.870 ;
        RECT 84.500 171.670 84.820 171.730 ;
        RECT 87.275 171.685 87.565 171.730 ;
        RECT 88.640 171.870 88.960 171.930 ;
        RECT 89.115 171.870 89.405 171.915 ;
        RECT 92.320 171.870 92.640 171.930 ;
        RECT 88.640 171.730 92.640 171.870 ;
        RECT 88.640 171.670 88.960 171.730 ;
        RECT 89.115 171.685 89.405 171.730 ;
        RECT 92.320 171.670 92.640 171.730 ;
        RECT 98.760 171.870 99.080 171.930 ;
        RECT 110.260 171.870 110.580 171.930 ;
        RECT 112.560 171.870 112.880 171.930 ;
        RECT 98.760 171.730 112.880 171.870 ;
        RECT 98.760 171.670 99.080 171.730 ;
        RECT 110.260 171.670 110.580 171.730 ;
        RECT 112.560 171.670 112.880 171.730 ;
        RECT 113.020 171.670 113.340 171.930 ;
        RECT 117.635 171.870 117.925 171.915 ;
        RECT 119.000 171.870 119.320 171.930 ;
        RECT 117.635 171.730 119.320 171.870 ;
        RECT 117.635 171.685 117.925 171.730 ;
        RECT 119.000 171.670 119.320 171.730 ;
        RECT 119.460 171.870 119.780 171.930 ;
        RECT 132.340 171.870 132.660 171.930 ;
        RECT 133.735 171.870 134.025 171.915 ;
        RECT 119.460 171.730 131.650 171.870 ;
        RECT 119.460 171.670 119.780 171.730 ;
        RECT 49.555 171.345 49.845 171.575 ;
        RECT 84.055 171.530 84.345 171.575 ;
        RECT 85.880 171.530 86.200 171.590 ;
        RECT 84.055 171.390 86.200 171.530 ;
        RECT 84.055 171.345 84.345 171.390 ;
        RECT 47.240 170.990 47.560 171.250 ;
        RECT 49.630 171.190 49.770 171.345 ;
        RECT 85.880 171.330 86.200 171.390 ;
        RECT 87.720 171.530 88.040 171.590 ;
        RECT 89.560 171.530 89.880 171.590 ;
        RECT 87.720 171.390 89.880 171.530 ;
        RECT 87.720 171.330 88.040 171.390 ;
        RECT 89.560 171.330 89.880 171.390 ;
        RECT 90.980 171.530 91.270 171.575 ;
        RECT 93.080 171.530 93.370 171.575 ;
        RECT 94.650 171.530 94.940 171.575 ;
        RECT 90.980 171.390 94.940 171.530 ;
        RECT 90.980 171.345 91.270 171.390 ;
        RECT 93.080 171.345 93.370 171.390 ;
        RECT 94.650 171.345 94.940 171.390 ;
        RECT 107.040 171.530 107.360 171.590 ;
        RECT 111.195 171.530 111.485 171.575 ;
        RECT 114.860 171.530 115.180 171.590 ;
        RECT 120.380 171.530 120.700 171.590 ;
        RECT 107.040 171.390 115.180 171.530 ;
        RECT 107.040 171.330 107.360 171.390 ;
        RECT 111.195 171.345 111.485 171.390 ;
        RECT 114.860 171.330 115.180 171.390 ;
        RECT 119.550 171.390 120.700 171.530 ;
        RECT 83.580 171.190 83.900 171.250 ;
        RECT 90.495 171.190 90.785 171.235 ;
        RECT 49.630 171.050 51.150 171.190 ;
        RECT 30.695 170.850 30.985 170.895 ;
        RECT 27.265 170.725 29.150 170.850 ;
        RECT 27.265 170.710 29.375 170.725 ;
        RECT 27.460 170.650 27.780 170.710 ;
        RECT 20.530 170.325 20.820 170.555 ;
        RECT 27.935 170.325 28.225 170.555 ;
        RECT 29.010 170.540 29.375 170.710 ;
        RECT 30.220 170.710 30.985 170.850 ;
        RECT 30.220 170.650 30.540 170.710 ;
        RECT 30.695 170.665 30.985 170.710 ;
        RECT 31.690 170.710 32.750 170.850 ;
        RECT 29.085 170.495 29.375 170.540 ;
        RECT 29.760 170.510 30.080 170.570 ;
        RECT 31.690 170.510 31.830 170.710 ;
        RECT 32.060 170.555 32.380 170.570 ;
        RECT 29.760 170.370 31.830 170.510 ;
        RECT 20.100 170.170 20.420 170.230 ;
        RECT 20.650 170.170 20.790 170.325 ;
        RECT 20.100 170.030 20.790 170.170 ;
        RECT 21.940 170.170 22.260 170.230 ;
        RECT 27.460 170.170 27.780 170.230 ;
        RECT 21.940 170.030 27.780 170.170 ;
        RECT 28.010 170.170 28.150 170.325 ;
        RECT 29.760 170.310 30.080 170.370 ;
        RECT 32.030 170.325 32.380 170.555 ;
        RECT 32.610 170.510 32.750 170.710 ;
        RECT 38.515 170.665 38.805 170.895 ;
        RECT 38.975 170.665 39.265 170.895 ;
        RECT 38.590 170.510 38.730 170.665 ;
        RECT 39.880 170.650 40.200 170.910 ;
        RECT 40.340 170.850 40.660 170.910 ;
        RECT 42.195 170.850 42.485 170.895 ;
        RECT 40.340 170.710 42.485 170.850 ;
        RECT 40.340 170.650 40.660 170.710 ;
        RECT 42.195 170.665 42.485 170.710 ;
        RECT 42.730 170.710 44.710 170.850 ;
        RECT 39.970 170.510 40.110 170.650 ;
        RECT 32.610 170.370 38.270 170.510 ;
        RECT 38.590 170.370 40.110 170.510 ;
        RECT 41.260 170.510 41.580 170.570 ;
        RECT 42.730 170.510 42.870 170.710 ;
        RECT 41.260 170.370 42.870 170.510 ;
        RECT 32.060 170.310 32.380 170.325 ;
        RECT 28.380 170.170 28.700 170.230 ;
        RECT 34.820 170.170 35.140 170.230 ;
        RECT 37.595 170.170 37.885 170.215 ;
        RECT 28.010 170.030 37.885 170.170 ;
        RECT 38.130 170.170 38.270 170.370 ;
        RECT 41.260 170.310 41.580 170.370 ;
        RECT 43.100 170.310 43.420 170.570 ;
        RECT 44.570 170.555 44.710 170.710 ;
        RECT 47.700 170.650 48.020 170.910 ;
        RECT 50.015 170.850 50.305 170.895 ;
        RECT 50.460 170.850 50.780 170.910 ;
        RECT 51.010 170.895 51.150 171.050 ;
        RECT 83.580 171.050 90.785 171.190 ;
        RECT 83.580 170.990 83.900 171.050 ;
        RECT 90.495 171.005 90.785 171.050 ;
        RECT 91.375 171.190 91.665 171.235 ;
        RECT 92.565 171.190 92.855 171.235 ;
        RECT 95.085 171.190 95.375 171.235 ;
        RECT 91.375 171.050 95.375 171.190 ;
        RECT 91.375 171.005 91.665 171.050 ;
        RECT 92.565 171.005 92.855 171.050 ;
        RECT 95.085 171.005 95.375 171.050 ;
        RECT 98.775 171.190 99.065 171.235 ;
        RECT 101.060 171.190 101.380 171.250 ;
        RECT 112.560 171.190 112.880 171.250 ;
        RECT 114.415 171.190 114.705 171.235 ;
        RECT 98.775 171.050 108.190 171.190 ;
        RECT 98.775 171.005 99.065 171.050 ;
        RECT 101.060 170.990 101.380 171.050 ;
        RECT 50.015 170.710 50.780 170.850 ;
        RECT 50.015 170.665 50.305 170.710 ;
        RECT 44.495 170.510 44.785 170.555 ;
        RECT 50.090 170.510 50.230 170.665 ;
        RECT 50.460 170.650 50.780 170.710 ;
        RECT 50.935 170.665 51.225 170.895 ;
        RECT 82.660 170.650 82.980 170.910 ;
        RECT 84.040 170.650 84.360 170.910 ;
        RECT 84.975 170.665 85.265 170.895 ;
        RECT 85.435 170.850 85.725 170.895 ;
        RECT 87.260 170.850 87.580 170.910 ;
        RECT 85.435 170.710 87.580 170.850 ;
        RECT 85.435 170.665 85.725 170.710 ;
        RECT 44.495 170.370 50.230 170.510 ;
        RECT 85.050 170.510 85.190 170.665 ;
        RECT 87.260 170.650 87.580 170.710 ;
        RECT 88.180 170.850 88.500 170.910 ;
        RECT 88.655 170.850 88.945 170.895 ;
        RECT 88.180 170.710 88.945 170.850 ;
        RECT 88.180 170.650 88.500 170.710 ;
        RECT 88.655 170.665 88.945 170.710 ;
        RECT 89.560 170.650 89.880 170.910 ;
        RECT 100.600 170.850 100.920 170.910 ;
        RECT 102.455 170.850 102.745 170.895 ;
        RECT 91.490 170.710 102.745 170.850 ;
        RECT 86.800 170.510 87.120 170.570 ;
        RECT 91.490 170.510 91.630 170.710 ;
        RECT 100.600 170.650 100.920 170.710 ;
        RECT 102.455 170.665 102.745 170.710 ;
        RECT 102.900 170.850 103.220 170.910 ;
        RECT 108.050 170.895 108.190 171.050 ;
        RECT 112.560 171.050 114.705 171.190 ;
        RECT 114.950 171.190 115.090 171.330 ;
        RECT 114.950 171.050 116.010 171.190 ;
        RECT 112.560 170.990 112.880 171.050 ;
        RECT 114.415 171.005 114.705 171.050 ;
        RECT 105.675 170.850 105.965 170.895 ;
        RECT 102.900 170.710 105.965 170.850 ;
        RECT 85.050 170.370 85.650 170.510 ;
        RECT 44.495 170.325 44.785 170.370 ;
        RECT 38.500 170.170 38.820 170.230 ;
        RECT 40.815 170.170 41.105 170.215 ;
        RECT 38.130 170.030 41.105 170.170 ;
        RECT 20.100 169.970 20.420 170.030 ;
        RECT 21.940 169.970 22.260 170.030 ;
        RECT 27.460 169.970 27.780 170.030 ;
        RECT 28.380 169.970 28.700 170.030 ;
        RECT 34.820 169.970 35.140 170.030 ;
        RECT 37.595 169.985 37.885 170.030 ;
        RECT 38.500 169.970 38.820 170.030 ;
        RECT 40.815 169.985 41.105 170.030 ;
        RECT 44.035 170.170 44.325 170.215 ;
        RECT 45.495 170.170 45.785 170.215 ;
        RECT 44.035 170.030 45.785 170.170 ;
        RECT 44.035 169.985 44.325 170.030 ;
        RECT 45.495 169.985 45.785 170.030 ;
        RECT 46.320 169.970 46.640 170.230 ;
        RECT 85.510 170.170 85.650 170.370 ;
        RECT 86.800 170.370 91.630 170.510 ;
        RECT 91.830 170.510 92.120 170.555 ;
        RECT 102.530 170.510 102.670 170.665 ;
        RECT 102.900 170.650 103.220 170.710 ;
        RECT 105.675 170.665 105.965 170.710 ;
        RECT 107.975 170.665 108.265 170.895 ;
        RECT 115.320 170.650 115.640 170.910 ;
        RECT 115.870 170.895 116.010 171.050 ;
        RECT 115.795 170.665 116.085 170.895 ;
        RECT 118.080 170.850 118.400 170.910 ;
        RECT 119.550 170.895 119.690 171.390 ;
        RECT 120.380 171.330 120.700 171.390 ;
        RECT 123.600 171.530 123.920 171.590 ;
        RECT 128.660 171.530 128.980 171.590 ;
        RECT 123.600 171.390 128.980 171.530 ;
        RECT 123.600 171.330 123.920 171.390 ;
        RECT 124.520 171.190 124.840 171.250 ;
        RECT 120.010 171.050 124.840 171.190 ;
        RECT 120.010 170.895 120.150 171.050 ;
        RECT 124.520 170.990 124.840 171.050 ;
        RECT 118.555 170.850 118.845 170.895 ;
        RECT 118.080 170.710 118.845 170.850 ;
        RECT 118.080 170.650 118.400 170.710 ;
        RECT 118.555 170.665 118.845 170.710 ;
        RECT 119.475 170.665 119.765 170.895 ;
        RECT 119.935 170.665 120.225 170.895 ;
        RECT 120.380 170.850 120.700 170.910 ;
        RECT 121.775 170.850 122.065 170.895 ;
        RECT 120.380 170.710 122.065 170.850 ;
        RECT 120.380 170.650 120.700 170.710 ;
        RECT 121.775 170.665 122.065 170.710 ;
        RECT 122.220 170.850 122.540 170.910 ;
        RECT 122.695 170.850 122.985 170.895 ;
        RECT 122.220 170.710 122.985 170.850 ;
        RECT 122.220 170.650 122.540 170.710 ;
        RECT 122.695 170.665 122.985 170.710 ;
        RECT 123.155 170.850 123.445 170.895 ;
        RECT 124.060 170.850 124.380 170.910 ;
        RECT 127.370 170.895 127.510 171.390 ;
        RECT 128.660 171.330 128.980 171.390 ;
        RECT 130.055 171.530 130.345 171.575 ;
        RECT 130.960 171.530 131.280 171.590 ;
        RECT 130.055 171.390 131.280 171.530 ;
        RECT 130.055 171.345 130.345 171.390 ;
        RECT 130.960 171.330 131.280 171.390 ;
        RECT 127.740 170.990 128.060 171.250 ;
        RECT 128.200 170.990 128.520 171.250 ;
        RECT 126.375 170.850 126.665 170.895 ;
        RECT 123.155 170.710 124.380 170.850 ;
        RECT 123.155 170.665 123.445 170.710 ;
        RECT 124.060 170.650 124.380 170.710 ;
        RECT 125.530 170.710 126.665 170.850 ;
        RECT 91.830 170.370 98.070 170.510 ;
        RECT 102.530 170.370 123.370 170.510 ;
        RECT 86.800 170.310 87.120 170.370 ;
        RECT 91.830 170.325 92.120 170.370 ;
        RECT 87.275 170.170 87.565 170.215 ;
        RECT 87.720 170.170 88.040 170.230 ;
        RECT 85.510 170.030 88.040 170.170 ;
        RECT 87.275 169.985 87.565 170.030 ;
        RECT 87.720 169.970 88.040 170.030 ;
        RECT 88.180 169.970 88.500 170.230 ;
        RECT 96.920 170.170 97.240 170.230 ;
        RECT 97.395 170.170 97.685 170.215 ;
        RECT 96.920 170.030 97.685 170.170 ;
        RECT 97.930 170.170 98.070 170.370 ;
        RECT 123.230 170.230 123.370 170.370 ;
        RECT 102.915 170.170 103.205 170.215 ;
        RECT 97.930 170.030 103.205 170.170 ;
        RECT 96.920 169.970 97.240 170.030 ;
        RECT 97.395 169.985 97.685 170.030 ;
        RECT 102.915 169.985 103.205 170.030 ;
        RECT 109.800 170.170 110.120 170.230 ;
        RECT 113.035 170.170 113.325 170.215 ;
        RECT 109.800 170.030 113.325 170.170 ;
        RECT 109.800 169.970 110.120 170.030 ;
        RECT 113.035 169.985 113.325 170.030 ;
        RECT 113.955 170.170 114.245 170.215 ;
        RECT 118.540 170.170 118.860 170.230 ;
        RECT 113.955 170.030 118.860 170.170 ;
        RECT 113.955 169.985 114.245 170.030 ;
        RECT 118.540 169.970 118.860 170.030 ;
        RECT 120.855 170.170 121.145 170.215 ;
        RECT 121.300 170.170 121.620 170.230 ;
        RECT 120.855 170.030 121.620 170.170 ;
        RECT 120.855 169.985 121.145 170.030 ;
        RECT 121.300 169.970 121.620 170.030 ;
        RECT 123.140 169.970 123.460 170.230 ;
        RECT 125.530 170.170 125.670 170.710 ;
        RECT 126.375 170.665 126.665 170.710 ;
        RECT 127.295 170.665 127.585 170.895 ;
        RECT 129.135 170.850 129.425 170.895 ;
        RECT 130.040 170.850 130.360 170.910 ;
        RECT 131.510 170.895 131.650 171.730 ;
        RECT 132.340 171.730 134.025 171.870 ;
        RECT 132.340 171.670 132.660 171.730 ;
        RECT 133.735 171.685 134.025 171.730 ;
        RECT 137.415 171.870 137.705 171.915 ;
        RECT 137.860 171.870 138.180 171.930 ;
        RECT 137.415 171.730 138.180 171.870 ;
        RECT 137.415 171.685 137.705 171.730 ;
        RECT 137.860 171.670 138.180 171.730 ;
        RECT 136.480 171.190 136.800 171.250 ;
        RECT 140.175 171.190 140.465 171.235 ;
        RECT 131.970 171.050 134.870 171.190 ;
        RECT 129.135 170.710 130.360 170.850 ;
        RECT 129.135 170.665 129.425 170.710 ;
        RECT 130.040 170.650 130.360 170.710 ;
        RECT 131.435 170.665 131.725 170.895 ;
        RECT 125.915 170.510 126.205 170.555 ;
        RECT 126.820 170.510 127.140 170.570 ;
        RECT 125.915 170.370 127.140 170.510 ;
        RECT 125.915 170.325 126.205 170.370 ;
        RECT 126.820 170.310 127.140 170.370 ;
        RECT 127.740 170.510 128.060 170.570 ;
        RECT 131.970 170.510 132.110 171.050 ;
        RECT 134.730 170.910 134.870 171.050 ;
        RECT 136.480 171.050 140.465 171.190 ;
        RECT 136.480 170.990 136.800 171.050 ;
        RECT 140.175 171.005 140.465 171.050 ;
        RECT 133.720 170.650 134.040 170.910 ;
        RECT 134.640 170.650 134.960 170.910 ;
        RECT 143.380 170.850 143.700 170.910 ;
        RECT 144.315 170.850 144.605 170.895 ;
        RECT 143.380 170.710 144.605 170.850 ;
        RECT 143.380 170.650 143.700 170.710 ;
        RECT 144.315 170.665 144.605 170.710 ;
        RECT 127.740 170.370 132.110 170.510 ;
        RECT 127.740 170.310 128.060 170.370 ;
        RECT 132.340 170.310 132.660 170.570 ;
        RECT 133.260 170.510 133.580 170.570 ;
        RECT 138.780 170.510 139.100 170.570 ;
        RECT 133.260 170.370 139.100 170.510 ;
        RECT 133.260 170.310 133.580 170.370 ;
        RECT 138.780 170.310 139.100 170.370 ;
        RECT 139.255 170.510 139.545 170.555 ;
        RECT 141.555 170.510 141.845 170.555 ;
        RECT 139.255 170.370 141.845 170.510 ;
        RECT 139.255 170.325 139.545 170.370 ;
        RECT 141.555 170.325 141.845 170.370 ;
        RECT 129.120 170.170 129.440 170.230 ;
        RECT 130.500 170.170 130.820 170.230 ;
        RECT 125.530 170.030 130.820 170.170 ;
        RECT 129.120 169.970 129.440 170.030 ;
        RECT 130.500 169.970 130.820 170.030 ;
        RECT 130.960 170.170 131.280 170.230 ;
        RECT 134.640 170.170 134.960 170.230 ;
        RECT 130.960 170.030 134.960 170.170 ;
        RECT 130.960 169.970 131.280 170.030 ;
        RECT 134.640 169.970 134.960 170.030 ;
        RECT 135.575 170.170 135.865 170.215 ;
        RECT 136.020 170.170 136.340 170.230 ;
        RECT 135.575 170.030 136.340 170.170 ;
        RECT 135.575 169.985 135.865 170.030 ;
        RECT 136.020 169.970 136.340 170.030 ;
        RECT 139.700 169.970 140.020 170.230 ;
        RECT 17.270 169.350 146.990 169.830 ;
        RECT 20.100 168.950 20.420 169.210 ;
        RECT 20.955 169.150 21.245 169.195 ;
        RECT 21.480 169.150 21.800 169.210 ;
        RECT 25.160 169.150 25.480 169.210 ;
        RECT 30.220 169.150 30.540 169.210 ;
        RECT 20.955 169.010 21.800 169.150 ;
        RECT 20.955 168.965 21.245 169.010 ;
        RECT 21.480 168.950 21.800 169.010 ;
        RECT 23.410 169.010 30.540 169.150 ;
        RECT 21.940 168.610 22.260 168.870 ;
        RECT 19.180 168.470 19.500 168.530 ;
        RECT 22.415 168.470 22.705 168.515 ;
        RECT 23.410 168.470 23.550 169.010 ;
        RECT 25.160 168.950 25.480 169.010 ;
        RECT 30.220 168.950 30.540 169.010 ;
        RECT 30.680 169.195 31.000 169.210 ;
        RECT 30.680 168.965 31.065 169.195 ;
        RECT 31.615 169.150 31.905 169.195 ;
        RECT 32.060 169.150 32.380 169.210 ;
        RECT 31.615 169.010 32.380 169.150 ;
        RECT 31.615 168.965 31.905 169.010 ;
        RECT 30.680 168.950 31.000 168.965 ;
        RECT 32.060 168.950 32.380 169.010 ;
        RECT 39.880 169.150 40.200 169.210 ;
        RECT 42.195 169.150 42.485 169.195 ;
        RECT 39.880 169.010 42.485 169.150 ;
        RECT 39.880 168.950 40.200 169.010 ;
        RECT 42.195 168.965 42.485 169.010 ;
        RECT 43.100 169.150 43.420 169.210 ;
        RECT 44.955 169.150 45.245 169.195 ;
        RECT 43.100 169.010 45.245 169.150 ;
        RECT 43.100 168.950 43.420 169.010 ;
        RECT 44.955 168.965 45.245 169.010 ;
        RECT 88.640 168.950 88.960 169.210 ;
        RECT 91.875 169.150 92.165 169.195 ;
        RECT 100.600 169.150 100.920 169.210 ;
        RECT 91.875 169.010 100.920 169.150 ;
        RECT 91.875 168.965 92.165 169.010 ;
        RECT 100.600 168.950 100.920 169.010 ;
        RECT 101.535 169.150 101.825 169.195 ;
        RECT 102.900 169.150 103.220 169.210 ;
        RECT 101.535 169.010 103.220 169.150 ;
        RECT 101.535 168.965 101.825 169.010 ;
        RECT 102.900 168.950 103.220 169.010 ;
        RECT 105.200 169.150 105.520 169.210 ;
        RECT 105.675 169.150 105.965 169.195 ;
        RECT 105.200 169.010 105.965 169.150 ;
        RECT 105.200 168.950 105.520 169.010 ;
        RECT 105.675 168.965 105.965 169.010 ;
        RECT 106.580 169.150 106.900 169.210 ;
        RECT 115.780 169.150 116.100 169.210 ;
        RECT 116.255 169.150 116.545 169.195 ;
        RECT 106.580 169.010 108.420 169.150 ;
        RECT 106.580 168.950 106.900 169.010 ;
        RECT 23.780 168.855 24.100 168.870 ;
        RECT 23.750 168.810 24.100 168.855 ;
        RECT 27.920 168.810 28.240 168.870 ;
        RECT 29.760 168.810 30.080 168.870 ;
        RECT 23.750 168.670 24.250 168.810 ;
        RECT 27.920 168.670 30.080 168.810 ;
        RECT 23.750 168.625 24.100 168.670 ;
        RECT 23.780 168.610 24.100 168.625 ;
        RECT 27.920 168.610 28.240 168.670 ;
        RECT 29.760 168.610 30.080 168.670 ;
        RECT 19.180 168.330 23.550 168.470 ;
        RECT 30.310 168.470 30.450 168.950 ;
        RECT 55.520 168.810 55.840 168.870 ;
        RECT 35.370 168.670 55.840 168.810 ;
        RECT 35.370 168.515 35.510 168.670 ;
        RECT 36.660 168.515 36.980 168.530 ;
        RECT 35.295 168.470 35.585 168.515 ;
        RECT 30.310 168.330 35.585 168.470 ;
        RECT 19.180 168.270 19.500 168.330 ;
        RECT 22.415 168.285 22.705 168.330 ;
        RECT 35.295 168.285 35.585 168.330 ;
        RECT 36.630 168.285 36.980 168.515 ;
        RECT 36.660 168.270 36.980 168.285 ;
        RECT 46.320 168.470 46.640 168.530 ;
        RECT 51.930 168.515 52.070 168.670 ;
        RECT 55.520 168.610 55.840 168.670 ;
        RECT 82.660 168.810 82.980 168.870 ;
        RECT 89.100 168.810 89.420 168.870 ;
        RECT 96.015 168.810 96.305 168.855 ;
        RECT 82.660 168.670 89.420 168.810 ;
        RECT 82.660 168.610 82.980 168.670 ;
        RECT 89.100 168.610 89.420 168.670 ;
        RECT 90.570 168.670 96.305 168.810 ;
        RECT 50.520 168.470 50.810 168.515 ;
        RECT 46.320 168.330 50.810 168.470 ;
        RECT 46.320 168.270 46.640 168.330 ;
        RECT 50.520 168.285 50.810 168.330 ;
        RECT 51.855 168.285 52.145 168.515 ;
        RECT 62.895 168.470 63.185 168.515 ;
        RECT 64.275 168.470 64.565 168.515 ;
        RECT 62.895 168.330 64.565 168.470 ;
        RECT 62.895 168.285 63.185 168.330 ;
        RECT 64.275 168.285 64.565 168.330 ;
        RECT 84.040 168.470 84.360 168.530 ;
        RECT 87.735 168.470 88.025 168.515 ;
        RECT 84.040 168.330 88.025 168.470 ;
        RECT 84.040 168.270 84.360 168.330 ;
        RECT 87.735 168.285 88.025 168.330 ;
        RECT 23.295 168.130 23.585 168.175 ;
        RECT 24.485 168.130 24.775 168.175 ;
        RECT 27.005 168.130 27.295 168.175 ;
        RECT 23.295 167.990 27.295 168.130 ;
        RECT 23.295 167.945 23.585 167.990 ;
        RECT 24.485 167.945 24.775 167.990 ;
        RECT 27.005 167.945 27.295 167.990 ;
        RECT 36.175 168.130 36.465 168.175 ;
        RECT 37.365 168.130 37.655 168.175 ;
        RECT 39.885 168.130 40.175 168.175 ;
        RECT 36.175 167.990 40.175 168.130 ;
        RECT 36.175 167.945 36.465 167.990 ;
        RECT 37.365 167.945 37.655 167.990 ;
        RECT 39.885 167.945 40.175 167.990 ;
        RECT 47.265 168.130 47.555 168.175 ;
        RECT 49.785 168.130 50.075 168.175 ;
        RECT 50.975 168.130 51.265 168.175 ;
        RECT 47.265 167.990 51.265 168.130 ;
        RECT 47.265 167.945 47.555 167.990 ;
        RECT 49.785 167.945 50.075 167.990 ;
        RECT 50.975 167.945 51.265 167.990 ;
        RECT 67.020 167.930 67.340 168.190 ;
        RECT 79.440 167.930 79.760 168.190 ;
        RECT 87.810 168.130 87.950 168.285 ;
        RECT 89.560 168.270 89.880 168.530 ;
        RECT 90.570 168.515 90.710 168.670 ;
        RECT 96.015 168.625 96.305 168.670 ;
        RECT 96.920 168.810 97.240 168.870 ;
        RECT 106.120 168.810 106.440 168.870 ;
        RECT 107.515 168.810 107.805 168.855 ;
        RECT 96.920 168.670 104.970 168.810 ;
        RECT 96.920 168.610 97.240 168.670 ;
        RECT 90.495 168.285 90.785 168.515 ;
        RECT 92.320 168.470 92.640 168.530 ;
        RECT 92.795 168.470 93.085 168.515 ;
        RECT 95.095 168.470 95.385 168.515 ;
        RECT 92.320 168.330 95.385 168.470 ;
        RECT 88.180 168.130 88.500 168.190 ;
        RECT 90.570 168.130 90.710 168.285 ;
        RECT 92.320 168.270 92.640 168.330 ;
        RECT 92.795 168.285 93.085 168.330 ;
        RECT 95.095 168.285 95.385 168.330 ;
        RECT 98.315 168.470 98.605 168.515 ;
        RECT 98.760 168.470 99.080 168.530 ;
        RECT 98.315 168.330 99.080 168.470 ;
        RECT 98.315 168.285 98.605 168.330 ;
        RECT 98.760 168.270 99.080 168.330 ;
        RECT 99.220 168.270 99.540 168.530 ;
        RECT 99.680 168.270 100.000 168.530 ;
        RECT 100.140 168.270 100.460 168.530 ;
        RECT 104.830 168.515 104.970 168.670 ;
        RECT 106.120 168.670 107.805 168.810 ;
        RECT 108.280 168.810 108.420 169.010 ;
        RECT 115.780 169.010 116.545 169.150 ;
        RECT 115.780 168.950 116.100 169.010 ;
        RECT 116.255 168.965 116.545 169.010 ;
        RECT 118.080 168.950 118.400 169.210 ;
        RECT 122.695 169.150 122.985 169.195 ;
        RECT 125.900 169.150 126.220 169.210 ;
        RECT 132.340 169.150 132.660 169.210 ;
        RECT 133.720 169.150 134.040 169.210 ;
        RECT 122.695 169.010 125.670 169.150 ;
        RECT 122.695 168.965 122.985 169.010 ;
        RECT 118.170 168.810 118.310 168.950 ;
        RECT 108.280 168.670 116.010 168.810 ;
        RECT 118.170 168.670 121.070 168.810 ;
        RECT 106.120 168.610 106.440 168.670 ;
        RECT 107.515 168.625 107.805 168.670 ;
        RECT 104.755 168.285 105.045 168.515 ;
        RECT 106.580 168.270 106.900 168.530 ;
        RECT 107.040 168.270 107.360 168.530 ;
        RECT 108.420 168.270 108.740 168.530 ;
        RECT 110.260 168.270 110.580 168.530 ;
        RECT 112.575 168.470 112.865 168.515 ;
        RECT 113.020 168.470 113.340 168.530 ;
        RECT 115.870 168.515 116.010 168.670 ;
        RECT 114.415 168.470 114.705 168.515 ;
        RECT 112.575 168.330 113.340 168.470 ;
        RECT 112.575 168.285 112.865 168.330 ;
        RECT 113.020 168.270 113.340 168.330 ;
        RECT 113.570 168.330 114.705 168.470 ;
        RECT 87.810 167.990 90.710 168.130 ;
        RECT 88.180 167.930 88.500 167.990 ;
        RECT 97.855 167.945 98.145 168.175 ;
        RECT 101.995 168.130 102.285 168.175 ;
        RECT 99.770 167.990 102.285 168.130 ;
        RECT 22.900 167.790 23.190 167.835 ;
        RECT 25.000 167.790 25.290 167.835 ;
        RECT 26.570 167.790 26.860 167.835 ;
        RECT 22.900 167.650 26.860 167.790 ;
        RECT 22.900 167.605 23.190 167.650 ;
        RECT 25.000 167.605 25.290 167.650 ;
        RECT 26.570 167.605 26.860 167.650 ;
        RECT 28.840 167.790 29.160 167.850 ;
        RECT 29.315 167.790 29.605 167.835 ;
        RECT 28.840 167.650 29.605 167.790 ;
        RECT 28.840 167.590 29.160 167.650 ;
        RECT 29.315 167.605 29.605 167.650 ;
        RECT 35.780 167.790 36.070 167.835 ;
        RECT 37.880 167.790 38.170 167.835 ;
        RECT 39.450 167.790 39.740 167.835 ;
        RECT 35.780 167.650 39.740 167.790 ;
        RECT 35.780 167.605 36.070 167.650 ;
        RECT 37.880 167.605 38.170 167.650 ;
        RECT 39.450 167.605 39.740 167.650 ;
        RECT 47.700 167.790 47.990 167.835 ;
        RECT 49.270 167.790 49.560 167.835 ;
        RECT 51.370 167.790 51.660 167.835 ;
        RECT 47.700 167.650 51.660 167.790 ;
        RECT 97.930 167.790 98.070 167.945 ;
        RECT 99.770 167.790 99.910 167.990 ;
        RECT 101.995 167.945 102.285 167.990 ;
        RECT 113.570 167.850 113.710 168.330 ;
        RECT 114.415 168.285 114.705 168.330 ;
        RECT 115.795 168.285 116.085 168.515 ;
        RECT 117.175 168.470 117.465 168.515 ;
        RECT 116.330 168.330 117.465 168.470 ;
        RECT 115.320 168.130 115.640 168.190 ;
        RECT 116.330 168.130 116.470 168.330 ;
        RECT 117.175 168.285 117.465 168.330 ;
        RECT 118.095 168.470 118.385 168.515 ;
        RECT 118.540 168.470 118.860 168.530 ;
        RECT 118.095 168.330 118.860 168.470 ;
        RECT 118.095 168.285 118.385 168.330 ;
        RECT 118.540 168.270 118.860 168.330 ;
        RECT 119.000 168.270 119.320 168.530 ;
        RECT 119.935 168.470 120.225 168.515 ;
        RECT 120.380 168.470 120.700 168.530 ;
        RECT 120.930 168.515 121.070 168.670 ;
        RECT 123.140 168.610 123.460 168.870 ;
        RECT 125.530 168.810 125.670 169.010 ;
        RECT 125.900 169.010 129.810 169.150 ;
        RECT 125.900 168.950 126.220 169.010 ;
        RECT 125.530 168.670 129.350 168.810 ;
        RECT 119.935 168.330 120.700 168.470 ;
        RECT 119.935 168.285 120.225 168.330 ;
        RECT 120.380 168.270 120.700 168.330 ;
        RECT 120.855 168.285 121.145 168.515 ;
        RECT 128.215 168.470 128.505 168.515 ;
        RECT 128.660 168.470 128.980 168.530 ;
        RECT 129.210 168.515 129.350 168.670 ;
        RECT 129.670 168.515 129.810 169.010 ;
        RECT 132.340 169.010 134.040 169.150 ;
        RECT 132.340 168.950 132.660 169.010 ;
        RECT 133.720 168.950 134.040 169.010 ;
        RECT 134.655 169.150 134.945 169.195 ;
        RECT 139.700 169.150 140.020 169.210 ;
        RECT 134.655 169.010 140.020 169.150 ;
        RECT 134.655 168.965 134.945 169.010 ;
        RECT 139.700 168.950 140.020 169.010 ;
        RECT 131.435 168.810 131.725 168.855 ;
        RECT 144.300 168.810 144.620 168.870 ;
        RECT 131.435 168.670 144.620 168.810 ;
        RECT 131.435 168.625 131.725 168.670 ;
        RECT 144.300 168.610 144.620 168.670 ;
        RECT 128.215 168.330 128.980 168.470 ;
        RECT 128.215 168.285 128.505 168.330 ;
        RECT 128.660 168.270 128.980 168.330 ;
        RECT 129.135 168.285 129.425 168.515 ;
        RECT 129.595 168.285 129.885 168.515 ;
        RECT 130.040 168.270 130.360 168.530 ;
        RECT 131.880 168.270 132.200 168.530 ;
        RECT 132.340 168.470 132.660 168.530 ;
        RECT 132.815 168.470 133.105 168.515 ;
        RECT 132.340 168.330 133.105 168.470 ;
        RECT 132.340 168.270 132.660 168.330 ;
        RECT 132.815 168.285 133.105 168.330 ;
        RECT 133.260 168.270 133.580 168.530 ;
        RECT 133.720 168.270 134.040 168.530 ;
        RECT 136.940 168.515 137.260 168.530 ;
        RECT 136.910 168.285 137.260 168.515 ;
        RECT 143.855 168.285 144.145 168.515 ;
        RECT 136.940 168.270 137.260 168.285 ;
        RECT 115.320 167.990 116.470 168.130 ;
        RECT 121.315 168.130 121.605 168.175 ;
        RECT 124.520 168.130 124.840 168.190 ;
        RECT 121.315 167.990 124.840 168.130 ;
        RECT 115.320 167.930 115.640 167.990 ;
        RECT 121.315 167.945 121.605 167.990 ;
        RECT 124.520 167.930 124.840 167.990 ;
        RECT 127.295 168.130 127.585 168.175 ;
        RECT 135.575 168.130 135.865 168.175 ;
        RECT 127.295 167.990 135.865 168.130 ;
        RECT 127.295 167.945 127.585 167.990 ;
        RECT 129.210 167.850 129.350 167.990 ;
        RECT 133.810 167.850 133.950 167.990 ;
        RECT 135.575 167.945 135.865 167.990 ;
        RECT 136.455 168.130 136.745 168.175 ;
        RECT 137.645 168.130 137.935 168.175 ;
        RECT 140.165 168.130 140.455 168.175 ;
        RECT 136.455 167.990 140.455 168.130 ;
        RECT 136.455 167.945 136.745 167.990 ;
        RECT 137.645 167.945 137.935 167.990 ;
        RECT 140.165 167.945 140.455 167.990 ;
        RECT 97.930 167.650 99.910 167.790 ;
        RECT 100.600 167.790 100.920 167.850 ;
        RECT 113.480 167.790 113.800 167.850 ;
        RECT 100.600 167.650 113.800 167.790 ;
        RECT 47.700 167.605 47.990 167.650 ;
        RECT 49.270 167.605 49.560 167.650 ;
        RECT 51.370 167.605 51.660 167.650 ;
        RECT 100.600 167.590 100.920 167.650 ;
        RECT 113.480 167.590 113.800 167.650 ;
        RECT 114.875 167.790 115.165 167.835 ;
        RECT 119.475 167.790 119.765 167.835 ;
        RECT 114.875 167.650 119.230 167.790 ;
        RECT 114.875 167.605 115.165 167.650 ;
        RECT 21.020 167.250 21.340 167.510 ;
        RECT 30.695 167.450 30.985 167.495 ;
        RECT 31.600 167.450 31.920 167.510 ;
        RECT 30.695 167.310 31.920 167.450 ;
        RECT 30.695 167.265 30.985 167.310 ;
        RECT 31.600 167.250 31.920 167.310 ;
        RECT 62.420 167.250 62.740 167.510 ;
        RECT 82.660 167.250 82.980 167.510 ;
        RECT 87.720 167.250 88.040 167.510 ;
        RECT 96.935 167.450 97.225 167.495 ;
        RECT 99.220 167.450 99.540 167.510 ;
        RECT 115.780 167.450 116.100 167.510 ;
        RECT 96.935 167.310 116.100 167.450 ;
        RECT 96.935 167.265 97.225 167.310 ;
        RECT 99.220 167.250 99.540 167.310 ;
        RECT 115.780 167.250 116.100 167.310 ;
        RECT 117.635 167.450 117.925 167.495 ;
        RECT 118.080 167.450 118.400 167.510 ;
        RECT 117.635 167.310 118.400 167.450 ;
        RECT 119.090 167.450 119.230 167.650 ;
        RECT 119.475 167.650 128.890 167.790 ;
        RECT 119.475 167.605 119.765 167.650 ;
        RECT 121.300 167.450 121.620 167.510 ;
        RECT 119.090 167.310 121.620 167.450 ;
        RECT 117.635 167.265 117.925 167.310 ;
        RECT 118.080 167.250 118.400 167.310 ;
        RECT 121.300 167.250 121.620 167.310 ;
        RECT 121.775 167.450 122.065 167.495 ;
        RECT 123.600 167.450 123.920 167.510 ;
        RECT 121.775 167.310 123.920 167.450 ;
        RECT 128.750 167.450 128.890 167.650 ;
        RECT 129.120 167.590 129.440 167.850 ;
        RECT 133.720 167.590 134.040 167.850 ;
        RECT 136.060 167.790 136.350 167.835 ;
        RECT 138.160 167.790 138.450 167.835 ;
        RECT 139.730 167.790 140.020 167.835 ;
        RECT 143.930 167.790 144.070 168.285 ;
        RECT 136.060 167.650 140.020 167.790 ;
        RECT 136.060 167.605 136.350 167.650 ;
        RECT 138.160 167.605 138.450 167.650 ;
        RECT 139.730 167.605 140.020 167.650 ;
        RECT 140.250 167.650 144.070 167.790 ;
        RECT 130.040 167.450 130.360 167.510 ;
        RECT 128.750 167.310 130.360 167.450 ;
        RECT 121.775 167.265 122.065 167.310 ;
        RECT 123.600 167.250 123.920 167.310 ;
        RECT 130.040 167.250 130.360 167.310 ;
        RECT 132.800 167.450 133.120 167.510 ;
        RECT 140.250 167.450 140.390 167.650 ;
        RECT 144.760 167.590 145.080 167.850 ;
        RECT 132.800 167.310 140.390 167.450 ;
        RECT 132.800 167.250 133.120 167.310 ;
        RECT 142.460 167.250 142.780 167.510 ;
        RECT 17.270 166.630 146.990 167.110 ;
        RECT 36.660 166.230 36.980 166.490 ;
        RECT 37.595 166.430 37.885 166.475 ;
        RECT 39.420 166.430 39.740 166.490 ;
        RECT 37.595 166.290 39.740 166.430 ;
        RECT 37.595 166.245 37.885 166.290 ;
        RECT 39.420 166.230 39.740 166.290 ;
        RECT 78.535 166.430 78.825 166.475 ;
        RECT 79.440 166.430 79.760 166.490 ;
        RECT 78.535 166.290 79.760 166.430 ;
        RECT 78.535 166.245 78.825 166.290 ;
        RECT 79.440 166.230 79.760 166.290 ;
        RECT 79.915 166.430 80.205 166.475 ;
        RECT 82.660 166.430 82.980 166.490 ;
        RECT 79.915 166.290 82.980 166.430 ;
        RECT 79.915 166.245 80.205 166.290 ;
        RECT 82.660 166.230 82.980 166.290 ;
        RECT 97.395 166.430 97.685 166.475 ;
        RECT 97.840 166.430 98.160 166.490 ;
        RECT 97.395 166.290 98.160 166.430 ;
        RECT 97.395 166.245 97.685 166.290 ;
        RECT 97.840 166.230 98.160 166.290 ;
        RECT 113.480 166.430 113.800 166.490 ;
        RECT 122.695 166.430 122.985 166.475 ;
        RECT 124.060 166.430 124.380 166.490 ;
        RECT 127.740 166.430 128.060 166.490 ;
        RECT 113.480 166.290 122.450 166.430 ;
        RECT 113.480 166.230 113.800 166.290 ;
        RECT 55.980 166.090 56.300 166.150 ;
        RECT 68.415 166.090 68.705 166.135 ;
        RECT 55.980 165.950 68.705 166.090 ;
        RECT 55.980 165.890 56.300 165.950 ;
        RECT 68.415 165.905 68.705 165.950 ;
        RECT 72.120 166.090 72.410 166.135 ;
        RECT 74.220 166.090 74.510 166.135 ;
        RECT 75.790 166.090 76.080 166.135 ;
        RECT 117.620 166.090 117.940 166.150 ;
        RECT 72.120 165.950 76.080 166.090 ;
        RECT 72.120 165.905 72.410 165.950 ;
        RECT 74.220 165.905 74.510 165.950 ;
        RECT 75.790 165.905 76.080 165.950 ;
        RECT 117.250 165.950 117.940 166.090 ;
        RECT 62.880 165.750 63.200 165.810 ;
        RECT 66.115 165.750 66.405 165.795 ;
        RECT 62.880 165.610 66.405 165.750 ;
        RECT 62.880 165.550 63.200 165.610 ;
        RECT 66.115 165.565 66.405 165.610 ;
        RECT 71.620 165.550 71.940 165.810 ;
        RECT 72.515 165.750 72.805 165.795 ;
        RECT 73.705 165.750 73.995 165.795 ;
        RECT 76.225 165.750 76.515 165.795 ;
        RECT 72.515 165.610 76.515 165.750 ;
        RECT 72.515 165.565 72.805 165.610 ;
        RECT 73.705 165.565 73.995 165.610 ;
        RECT 76.225 165.565 76.515 165.610 ;
        RECT 96.920 165.750 97.240 165.810 ;
        RECT 117.250 165.795 117.390 165.950 ;
        RECT 117.620 165.890 117.940 165.950 ;
        RECT 118.540 166.090 118.860 166.150 ;
        RECT 118.540 165.950 121.990 166.090 ;
        RECT 118.540 165.890 118.860 165.950 ;
        RECT 96.920 165.610 98.530 165.750 ;
        RECT 96.920 165.550 97.240 165.610 ;
        RECT 57.360 165.410 57.680 165.470 ;
        RECT 58.755 165.410 59.045 165.455 ;
        RECT 57.360 165.270 59.045 165.410 ;
        RECT 57.360 165.210 57.680 165.270 ;
        RECT 58.755 165.225 59.045 165.270 ;
        RECT 63.340 165.210 63.660 165.470 ;
        RECT 64.720 165.210 65.040 165.470 ;
        RECT 67.480 165.410 67.800 165.470 ;
        RECT 70.255 165.410 70.545 165.455 ;
        RECT 67.480 165.270 70.545 165.410 ;
        RECT 67.480 165.210 67.800 165.270 ;
        RECT 70.255 165.225 70.545 165.270 ;
        RECT 71.175 165.410 71.465 165.455 ;
        RECT 71.175 165.270 74.150 165.410 ;
        RECT 71.175 165.225 71.465 165.270 ;
        RECT 74.010 165.130 74.150 165.270 ;
        RECT 97.380 165.210 97.700 165.470 ;
        RECT 98.390 165.455 98.530 165.610 ;
        RECT 117.175 165.565 117.465 165.795 ;
        RECT 98.315 165.225 98.605 165.455 ;
        RECT 109.800 165.410 110.120 165.470 ;
        RECT 112.115 165.410 112.405 165.455 ;
        RECT 109.800 165.270 112.405 165.410 ;
        RECT 109.800 165.210 110.120 165.270 ;
        RECT 112.115 165.225 112.405 165.270 ;
        RECT 115.780 165.210 116.100 165.470 ;
        RECT 116.715 165.410 117.005 165.455 ;
        RECT 116.330 165.270 117.005 165.410 ;
        RECT 116.330 165.130 116.470 165.270 ;
        RECT 116.715 165.225 117.005 165.270 ;
        RECT 117.620 165.210 117.940 165.470 ;
        RECT 118.095 165.410 118.385 165.455 ;
        RECT 118.540 165.410 118.860 165.470 ;
        RECT 120.380 165.410 120.700 165.470 ;
        RECT 121.850 165.455 121.990 165.950 ;
        RECT 122.310 165.750 122.450 166.290 ;
        RECT 122.695 166.290 128.060 166.430 ;
        RECT 122.695 166.245 122.985 166.290 ;
        RECT 124.060 166.230 124.380 166.290 ;
        RECT 127.740 166.230 128.060 166.290 ;
        RECT 129.595 166.430 129.885 166.475 ;
        RECT 131.435 166.430 131.725 166.475 ;
        RECT 129.595 166.290 131.190 166.430 ;
        RECT 129.595 166.245 129.885 166.290 ;
        RECT 131.050 166.090 131.190 166.290 ;
        RECT 131.435 166.290 135.790 166.430 ;
        RECT 131.435 166.245 131.725 166.290 ;
        RECT 134.195 166.090 134.485 166.135 ;
        RECT 131.050 165.950 134.485 166.090 ;
        RECT 134.195 165.905 134.485 165.950 ;
        RECT 127.740 165.750 128.060 165.810 ;
        RECT 129.135 165.750 129.425 165.795 ;
        RECT 129.580 165.750 129.900 165.810 ;
        RECT 122.310 165.610 122.910 165.750 ;
        RECT 122.770 165.455 122.910 165.610 ;
        RECT 127.740 165.610 129.900 165.750 ;
        RECT 127.740 165.550 128.060 165.610 ;
        RECT 129.135 165.565 129.425 165.610 ;
        RECT 129.580 165.550 129.900 165.610 ;
        RECT 132.340 165.750 132.660 165.810 ;
        RECT 133.735 165.750 134.025 165.795 ;
        RECT 132.340 165.610 134.025 165.750 ;
        RECT 135.650 165.750 135.790 166.290 ;
        RECT 136.940 166.230 137.260 166.490 ;
        RECT 139.715 165.750 140.005 165.795 ;
        RECT 142.460 165.750 142.780 165.810 ;
        RECT 143.855 165.750 144.145 165.795 ;
        RECT 135.650 165.610 140.005 165.750 ;
        RECT 132.340 165.550 132.660 165.610 ;
        RECT 133.735 165.565 134.025 165.610 ;
        RECT 139.715 165.565 140.005 165.610 ;
        RECT 140.710 165.610 144.145 165.750 ;
        RECT 118.095 165.270 120.700 165.410 ;
        RECT 118.095 165.225 118.385 165.270 ;
        RECT 118.540 165.210 118.860 165.270 ;
        RECT 120.380 165.210 120.700 165.270 ;
        RECT 121.775 165.225 122.065 165.455 ;
        RECT 122.695 165.410 122.985 165.455 ;
        RECT 123.600 165.410 123.920 165.470 ;
        RECT 122.695 165.270 123.920 165.410 ;
        RECT 122.695 165.225 122.985 165.270 ;
        RECT 123.600 165.210 123.920 165.270 ;
        RECT 125.455 165.410 125.745 165.455 ;
        RECT 128.660 165.410 128.980 165.470 ;
        RECT 125.455 165.270 128.980 165.410 ;
        RECT 125.455 165.225 125.745 165.270 ;
        RECT 128.660 165.210 128.980 165.270 ;
        RECT 130.500 165.210 130.820 165.470 ;
        RECT 130.960 165.410 131.280 165.470 ;
        RECT 134.180 165.410 134.500 165.470 ;
        RECT 134.655 165.410 134.945 165.455 ;
        RECT 130.960 165.270 134.945 165.410 ;
        RECT 130.960 165.210 131.280 165.270 ;
        RECT 134.180 165.210 134.500 165.270 ;
        RECT 134.655 165.225 134.945 165.270 ;
        RECT 135.100 165.210 135.420 165.470 ;
        RECT 135.575 165.410 135.865 165.455 ;
        RECT 140.710 165.410 140.850 165.610 ;
        RECT 142.460 165.550 142.780 165.610 ;
        RECT 143.855 165.565 144.145 165.610 ;
        RECT 135.575 165.270 140.850 165.410 ;
        RECT 135.575 165.225 135.865 165.270 ;
        RECT 37.515 165.070 37.805 165.115 ;
        RECT 38.040 165.070 38.360 165.130 ;
        RECT 37.515 164.930 38.360 165.070 ;
        RECT 37.515 164.885 37.805 164.930 ;
        RECT 38.040 164.870 38.360 164.930 ;
        RECT 38.500 164.870 38.820 165.130 ;
        RECT 61.500 165.070 61.820 165.130 ;
        RECT 62.435 165.070 62.725 165.115 ;
        RECT 61.500 164.930 62.725 165.070 ;
        RECT 61.500 164.870 61.820 164.930 ;
        RECT 62.435 164.885 62.725 164.930 ;
        RECT 64.275 165.070 64.565 165.115 ;
        RECT 67.020 165.070 67.340 165.130 ;
        RECT 64.275 164.930 67.340 165.070 ;
        RECT 64.275 164.885 64.565 164.930 ;
        RECT 67.020 164.870 67.340 164.930 ;
        RECT 67.955 164.885 68.245 165.115 ;
        RECT 69.320 165.070 69.640 165.130 ;
        RECT 73.000 165.115 73.320 165.130 ;
        RECT 70.715 165.070 71.005 165.115 ;
        RECT 69.320 164.930 71.005 165.070 ;
        RECT 61.960 164.530 62.280 164.790 ;
        RECT 64.720 164.730 65.040 164.790 ;
        RECT 68.030 164.730 68.170 164.885 ;
        RECT 69.320 164.870 69.640 164.930 ;
        RECT 70.715 164.885 71.005 164.930 ;
        RECT 72.970 164.885 73.320 165.115 ;
        RECT 73.000 164.870 73.320 164.885 ;
        RECT 73.920 164.870 74.240 165.130 ;
        RECT 74.840 165.070 75.160 165.130 ;
        RECT 79.755 165.070 80.045 165.115 ;
        RECT 80.360 165.070 80.680 165.130 ;
        RECT 74.840 164.930 80.680 165.070 ;
        RECT 74.840 164.870 75.160 164.930 ;
        RECT 79.755 164.885 80.045 164.930 ;
        RECT 80.360 164.870 80.680 164.930 ;
        RECT 80.835 165.070 81.125 165.115 ;
        RECT 82.660 165.070 82.980 165.130 ;
        RECT 80.835 164.930 82.980 165.070 ;
        RECT 80.835 164.885 81.125 164.930 ;
        RECT 82.660 164.870 82.980 164.930 ;
        RECT 116.240 164.870 116.560 165.130 ;
        RECT 124.520 165.070 124.840 165.130 ;
        RECT 126.835 165.070 127.125 165.115 ;
        RECT 124.520 164.930 127.125 165.070 ;
        RECT 124.520 164.870 124.840 164.930 ;
        RECT 126.835 164.885 127.125 164.930 ;
        RECT 127.755 165.070 128.045 165.115 ;
        RECT 128.200 165.070 128.520 165.130 ;
        RECT 129.580 165.070 129.900 165.130 ;
        RECT 138.795 165.070 139.085 165.115 ;
        RECT 141.095 165.070 141.385 165.115 ;
        RECT 127.755 164.930 129.350 165.070 ;
        RECT 127.755 164.885 128.045 164.930 ;
        RECT 128.200 164.870 128.520 164.930 ;
        RECT 64.720 164.590 68.170 164.730 ;
        RECT 64.720 164.530 65.040 164.590 ;
        RECT 78.980 164.530 79.300 164.790 ;
        RECT 113.940 164.730 114.260 164.790 ;
        RECT 115.335 164.730 115.625 164.775 ;
        RECT 113.940 164.590 115.625 164.730 ;
        RECT 113.940 164.530 114.260 164.590 ;
        RECT 115.335 164.545 115.625 164.590 ;
        RECT 119.000 164.530 119.320 164.790 ;
        RECT 128.660 164.530 128.980 164.790 ;
        RECT 129.210 164.730 129.350 164.930 ;
        RECT 129.580 164.930 138.550 165.070 ;
        RECT 129.580 164.870 129.900 164.930 ;
        RECT 135.100 164.730 135.420 164.790 ;
        RECT 129.210 164.590 135.420 164.730 ;
        RECT 135.100 164.530 135.420 164.590 ;
        RECT 136.495 164.730 136.785 164.775 ;
        RECT 137.860 164.730 138.180 164.790 ;
        RECT 136.495 164.590 138.180 164.730 ;
        RECT 138.410 164.730 138.550 164.930 ;
        RECT 138.795 164.930 141.385 165.070 ;
        RECT 138.795 164.885 139.085 164.930 ;
        RECT 141.095 164.885 141.385 164.930 ;
        RECT 139.255 164.730 139.545 164.775 ;
        RECT 138.410 164.590 139.545 164.730 ;
        RECT 136.495 164.545 136.785 164.590 ;
        RECT 137.860 164.530 138.180 164.590 ;
        RECT 139.255 164.545 139.545 164.590 ;
        RECT 17.270 163.910 146.990 164.390 ;
        RECT 57.360 163.510 57.680 163.770 ;
        RECT 57.835 163.525 58.125 163.755 ;
        RECT 62.420 163.710 62.740 163.770 ;
        RECT 59.750 163.570 62.740 163.710 ;
        RECT 57.910 163.370 58.050 163.525 ;
        RECT 59.750 163.370 59.890 163.570 ;
        RECT 62.420 163.510 62.740 163.570 ;
        RECT 68.415 163.710 68.705 163.755 ;
        RECT 73.000 163.710 73.320 163.770 ;
        RECT 68.415 163.570 73.320 163.710 ;
        RECT 68.415 163.525 68.705 163.570 ;
        RECT 73.000 163.510 73.320 163.570 ;
        RECT 82.660 163.510 82.980 163.770 ;
        RECT 109.800 163.510 110.120 163.770 ;
        RECT 111.195 163.525 111.485 163.755 ;
        RECT 114.415 163.710 114.705 163.755 ;
        RECT 113.110 163.570 114.705 163.710 ;
        RECT 57.910 163.230 59.890 163.370 ;
        RECT 60.090 163.370 60.380 163.415 ;
        RECT 61.960 163.370 62.280 163.430 ;
        RECT 78.980 163.370 79.300 163.430 ;
        RECT 60.090 163.230 62.280 163.370 ;
        RECT 60.090 163.185 60.380 163.230 ;
        RECT 61.960 163.170 62.280 163.230 ;
        RECT 72.630 163.230 79.300 163.370 ;
        RECT 82.750 163.370 82.890 163.510 ;
        RECT 87.735 163.370 88.025 163.415 ;
        RECT 82.750 163.230 88.025 163.370 ;
        RECT 18.735 163.030 19.025 163.075 ;
        RECT 15.960 162.890 19.025 163.030 ;
        RECT 15.960 162.830 16.280 162.890 ;
        RECT 18.735 162.845 19.025 162.890 ;
        RECT 55.980 162.830 56.300 163.090 ;
        RECT 58.295 162.845 58.585 163.075 ;
        RECT 59.200 163.030 59.520 163.090 ;
        RECT 66.115 163.030 66.405 163.075 ;
        RECT 70.700 163.030 71.020 163.090 ;
        RECT 72.630 163.075 72.770 163.230 ;
        RECT 78.980 163.170 79.300 163.230 ;
        RECT 59.200 162.890 64.030 163.030 ;
        RECT 19.655 162.350 19.945 162.395 ;
        RECT 57.820 162.350 58.140 162.410 ;
        RECT 19.655 162.210 58.140 162.350 ;
        RECT 19.655 162.165 19.945 162.210 ;
        RECT 57.820 162.150 58.140 162.210 ;
        RECT 58.370 162.010 58.510 162.845 ;
        RECT 59.200 162.830 59.520 162.890 ;
        RECT 58.740 162.490 59.060 162.750 ;
        RECT 59.635 162.690 59.925 162.735 ;
        RECT 60.825 162.690 61.115 162.735 ;
        RECT 63.345 162.690 63.635 162.735 ;
        RECT 59.635 162.550 63.635 162.690 ;
        RECT 63.890 162.690 64.030 162.890 ;
        RECT 66.115 162.890 71.020 163.030 ;
        RECT 66.115 162.845 66.405 162.890 ;
        RECT 70.700 162.830 71.020 162.890 ;
        RECT 72.555 162.845 72.845 163.075 ;
        RECT 77.110 163.030 77.400 163.075 ;
        RECT 85.420 163.030 85.740 163.090 ;
        RECT 85.970 163.075 86.110 163.230 ;
        RECT 87.735 163.185 88.025 163.230 ;
        RECT 104.250 163.370 104.540 163.415 ;
        RECT 111.270 163.370 111.410 163.525 ;
        RECT 104.250 163.230 111.410 163.370 ;
        RECT 104.250 163.185 104.540 163.230 ;
        RECT 112.560 163.170 112.880 163.430 ;
        RECT 113.110 163.415 113.250 163.570 ;
        RECT 114.415 163.525 114.705 163.570 ;
        RECT 117.175 163.710 117.465 163.755 ;
        RECT 117.620 163.710 117.940 163.770 ;
        RECT 117.175 163.570 117.940 163.710 ;
        RECT 117.175 163.525 117.465 163.570 ;
        RECT 117.620 163.510 117.940 163.570 ;
        RECT 123.615 163.710 123.905 163.755 ;
        RECT 129.580 163.710 129.900 163.770 ;
        RECT 123.615 163.570 129.900 163.710 ;
        RECT 123.615 163.525 123.905 163.570 ;
        RECT 129.580 163.510 129.900 163.570 ;
        RECT 130.515 163.710 130.805 163.755 ;
        RECT 132.800 163.710 133.120 163.770 ;
        RECT 130.515 163.570 133.120 163.710 ;
        RECT 130.515 163.525 130.805 163.570 ;
        RECT 132.800 163.510 133.120 163.570 ;
        RECT 133.275 163.710 133.565 163.755 ;
        RECT 143.395 163.710 143.685 163.755 ;
        RECT 143.840 163.710 144.160 163.770 ;
        RECT 133.275 163.570 142.230 163.710 ;
        RECT 133.275 163.525 133.565 163.570 ;
        RECT 113.035 163.185 113.325 163.415 ;
        RECT 118.095 163.370 118.385 163.415 ;
        RECT 119.460 163.370 119.780 163.430 ;
        RECT 127.740 163.370 128.060 163.430 ;
        RECT 140.620 163.370 140.940 163.430 ;
        RECT 142.090 163.370 142.230 163.570 ;
        RECT 143.395 163.570 144.160 163.710 ;
        RECT 143.395 163.525 143.685 163.570 ;
        RECT 143.840 163.510 144.160 163.570 ;
        RECT 144.760 163.510 145.080 163.770 ;
        RECT 145.220 163.370 145.540 163.430 ;
        RECT 115.410 163.230 128.060 163.370 ;
        RECT 77.110 162.890 85.740 163.030 ;
        RECT 77.110 162.845 77.400 162.890 ;
        RECT 85.420 162.830 85.740 162.890 ;
        RECT 85.895 162.845 86.185 163.075 ;
        RECT 86.815 162.845 87.105 163.075 ;
        RECT 88.640 163.030 88.960 163.090 ;
        RECT 90.495 163.030 90.785 163.075 ;
        RECT 88.640 162.890 90.785 163.030 ;
        RECT 68.860 162.690 69.180 162.750 ;
        RECT 69.335 162.690 69.625 162.735 ;
        RECT 63.890 162.550 69.625 162.690 ;
        RECT 59.635 162.505 59.925 162.550 ;
        RECT 60.825 162.505 61.115 162.550 ;
        RECT 63.345 162.505 63.635 162.550 ;
        RECT 68.860 162.490 69.180 162.550 ;
        RECT 69.335 162.505 69.625 162.550 ;
        RECT 71.620 162.690 71.940 162.750 ;
        RECT 73.460 162.690 73.780 162.750 ;
        RECT 75.775 162.690 76.065 162.735 ;
        RECT 71.620 162.550 76.065 162.690 ;
        RECT 71.620 162.490 71.940 162.550 ;
        RECT 73.460 162.490 73.780 162.550 ;
        RECT 75.775 162.505 76.065 162.550 ;
        RECT 76.655 162.690 76.945 162.735 ;
        RECT 77.845 162.690 78.135 162.735 ;
        RECT 80.365 162.690 80.655 162.735 ;
        RECT 76.655 162.550 80.655 162.690 ;
        RECT 76.655 162.505 76.945 162.550 ;
        RECT 77.845 162.505 78.135 162.550 ;
        RECT 80.365 162.505 80.655 162.550 ;
        RECT 80.820 162.690 81.140 162.750 ;
        RECT 86.340 162.690 86.660 162.750 ;
        RECT 86.890 162.690 87.030 162.845 ;
        RECT 88.640 162.830 88.960 162.890 ;
        RECT 90.495 162.845 90.785 162.890 ;
        RECT 101.060 163.030 101.380 163.090 ;
        RECT 102.915 163.030 103.205 163.075 ;
        RECT 101.060 162.890 103.205 163.030 ;
        RECT 101.060 162.830 101.380 162.890 ;
        RECT 102.915 162.845 103.205 162.890 ;
        RECT 112.115 162.845 112.405 163.075 ;
        RECT 80.820 162.550 87.030 162.690 ;
        RECT 92.795 162.690 93.085 162.735 ;
        RECT 93.240 162.690 93.560 162.750 ;
        RECT 92.795 162.550 93.560 162.690 ;
        RECT 80.820 162.490 81.140 162.550 ;
        RECT 86.340 162.490 86.660 162.550 ;
        RECT 92.795 162.505 93.085 162.550 ;
        RECT 93.240 162.490 93.560 162.550 ;
        RECT 103.795 162.690 104.085 162.735 ;
        RECT 104.985 162.690 105.275 162.735 ;
        RECT 107.505 162.690 107.795 162.735 ;
        RECT 103.795 162.550 107.795 162.690 ;
        RECT 112.190 162.690 112.330 162.845 ;
        RECT 113.940 162.830 114.260 163.090 ;
        RECT 115.410 162.690 115.550 163.230 ;
        RECT 118.095 163.185 118.385 163.230 ;
        RECT 119.460 163.170 119.780 163.230 ;
        RECT 127.740 163.170 128.060 163.230 ;
        RECT 131.970 163.230 141.770 163.370 ;
        RECT 142.090 163.230 145.540 163.370 ;
        RECT 116.240 162.830 116.560 163.090 ;
        RECT 116.715 162.845 117.005 163.075 ;
        RECT 118.540 163.030 118.860 163.090 ;
        RECT 119.015 163.030 119.305 163.075 ;
        RECT 118.540 162.890 119.305 163.030 ;
        RECT 112.190 162.550 115.550 162.690 ;
        RECT 103.795 162.505 104.085 162.550 ;
        RECT 104.985 162.505 105.275 162.550 ;
        RECT 107.505 162.505 107.795 162.550 ;
        RECT 115.780 162.490 116.100 162.750 ;
        RECT 116.790 162.690 116.930 162.845 ;
        RECT 118.540 162.830 118.860 162.890 ;
        RECT 119.015 162.845 119.305 162.890 ;
        RECT 119.935 163.030 120.225 163.075 ;
        RECT 120.855 163.030 121.145 163.075 ;
        RECT 119.935 162.890 121.145 163.030 ;
        RECT 119.935 162.845 120.225 162.890 ;
        RECT 120.855 162.845 121.145 162.890 ;
        RECT 121.300 163.030 121.620 163.090 ;
        RECT 121.775 163.030 122.065 163.075 ;
        RECT 121.300 162.890 122.065 163.030 ;
        RECT 121.300 162.830 121.620 162.890 ;
        RECT 121.775 162.845 122.065 162.890 ;
        RECT 122.220 162.830 122.540 163.090 ;
        RECT 122.695 163.030 122.985 163.075 ;
        RECT 123.600 163.030 123.920 163.090 ;
        RECT 122.695 162.890 123.920 163.030 ;
        RECT 122.695 162.845 122.985 162.890 ;
        RECT 123.600 162.830 123.920 162.890 ;
        RECT 129.595 163.030 129.885 163.075 ;
        RECT 131.970 163.030 132.110 163.230 ;
        RECT 140.620 163.170 140.940 163.230 ;
        RECT 129.595 162.890 132.110 163.030 ;
        RECT 129.595 162.845 129.885 162.890 ;
        RECT 132.340 162.830 132.660 163.090 ;
        RECT 134.180 162.830 134.500 163.090 ;
        RECT 136.480 162.830 136.800 163.090 ;
        RECT 141.630 163.075 141.770 163.230 ;
        RECT 145.220 163.170 145.540 163.230 ;
        RECT 136.955 163.030 137.245 163.075 ;
        RECT 138.795 163.030 139.085 163.075 ;
        RECT 136.955 162.890 139.085 163.030 ;
        RECT 136.955 162.845 137.245 162.890 ;
        RECT 138.795 162.845 139.085 162.890 ;
        RECT 141.555 162.845 141.845 163.075 ;
        RECT 142.475 163.030 142.765 163.075 ;
        RECT 143.380 163.030 143.700 163.090 ;
        RECT 142.475 162.890 143.700 163.030 ;
        RECT 142.475 162.845 142.765 162.890 ;
        RECT 143.380 162.830 143.700 162.890 ;
        RECT 143.855 163.030 144.145 163.075 ;
        RECT 143.855 162.890 144.990 163.030 ;
        RECT 143.855 162.845 144.145 162.890 ;
        RECT 127.740 162.690 128.060 162.750 ;
        RECT 137.415 162.690 137.705 162.735 ;
        RECT 116.790 162.550 117.390 162.690 ;
        RECT 59.240 162.350 59.530 162.395 ;
        RECT 61.340 162.350 61.630 162.395 ;
        RECT 62.910 162.350 63.200 162.395 ;
        RECT 59.240 162.210 63.200 162.350 ;
        RECT 59.240 162.165 59.530 162.210 ;
        RECT 61.340 162.165 61.630 162.210 ;
        RECT 62.910 162.165 63.200 162.210 ;
        RECT 67.480 162.150 67.800 162.410 ;
        RECT 69.795 162.350 70.085 162.395 ;
        RECT 74.840 162.350 75.160 162.410 ;
        RECT 69.795 162.210 75.160 162.350 ;
        RECT 69.795 162.165 70.085 162.210 ;
        RECT 74.840 162.150 75.160 162.210 ;
        RECT 76.260 162.350 76.550 162.395 ;
        RECT 78.360 162.350 78.650 162.395 ;
        RECT 79.930 162.350 80.220 162.395 ;
        RECT 76.260 162.210 80.220 162.350 ;
        RECT 76.260 162.165 76.550 162.210 ;
        RECT 78.360 162.165 78.650 162.210 ;
        RECT 79.930 162.165 80.220 162.210 ;
        RECT 103.400 162.350 103.690 162.395 ;
        RECT 105.500 162.350 105.790 162.395 ;
        RECT 107.070 162.350 107.360 162.395 ;
        RECT 103.400 162.210 107.360 162.350 ;
        RECT 103.400 162.165 103.690 162.210 ;
        RECT 105.500 162.165 105.790 162.210 ;
        RECT 107.070 162.165 107.360 162.210 ;
        RECT 112.100 162.350 112.420 162.410 ;
        RECT 117.250 162.350 117.390 162.550 ;
        RECT 127.740 162.550 137.705 162.690 ;
        RECT 127.740 162.490 128.060 162.550 ;
        RECT 137.415 162.505 137.705 162.550 ;
        RECT 121.300 162.350 121.620 162.410 ;
        RECT 130.500 162.350 130.820 162.410 ;
        RECT 112.100 162.210 116.930 162.350 ;
        RECT 117.250 162.210 121.620 162.350 ;
        RECT 112.100 162.150 112.420 162.210 ;
        RECT 60.580 162.010 60.900 162.070 ;
        RECT 58.370 161.870 60.900 162.010 ;
        RECT 60.580 161.810 60.900 161.870 ;
        RECT 65.655 162.010 65.945 162.055 ;
        RECT 67.020 162.010 67.340 162.070 ;
        RECT 67.940 162.010 68.260 162.070 ;
        RECT 65.655 161.870 68.260 162.010 ;
        RECT 65.655 161.825 65.945 161.870 ;
        RECT 67.020 161.810 67.340 161.870 ;
        RECT 67.940 161.810 68.260 161.870 ;
        RECT 71.620 161.810 71.940 162.070 ;
        RECT 75.315 162.010 75.605 162.055 ;
        RECT 75.760 162.010 76.080 162.070 ;
        RECT 75.315 161.870 76.080 162.010 ;
        RECT 75.315 161.825 75.605 161.870 ;
        RECT 75.760 161.810 76.080 161.870 ;
        RECT 83.120 161.810 83.440 162.070 ;
        RECT 88.180 161.810 88.500 162.070 ;
        RECT 115.320 161.810 115.640 162.070 ;
        RECT 116.790 162.010 116.930 162.210 ;
        RECT 121.300 162.150 121.620 162.210 ;
        RECT 123.230 162.210 130.820 162.350 ;
        RECT 123.230 162.010 123.370 162.210 ;
        RECT 130.500 162.150 130.820 162.210 ;
        RECT 131.435 162.350 131.725 162.395 ;
        RECT 142.920 162.350 143.240 162.410 ;
        RECT 131.435 162.210 143.240 162.350 ;
        RECT 131.435 162.165 131.725 162.210 ;
        RECT 142.920 162.150 143.240 162.210 ;
        RECT 116.790 161.870 123.370 162.010 ;
        RECT 123.600 162.010 123.920 162.070 ;
        RECT 124.520 162.010 124.840 162.070 ;
        RECT 133.260 162.010 133.580 162.070 ;
        RECT 123.600 161.870 133.580 162.010 ;
        RECT 123.600 161.810 123.920 161.870 ;
        RECT 124.520 161.810 124.840 161.870 ;
        RECT 133.260 161.810 133.580 161.870 ;
        RECT 134.655 162.010 134.945 162.055 ;
        RECT 135.100 162.010 135.420 162.070 ;
        RECT 134.655 161.870 135.420 162.010 ;
        RECT 134.655 161.825 134.945 161.870 ;
        RECT 135.100 161.810 135.420 161.870 ;
        RECT 137.860 162.010 138.180 162.070 ;
        RECT 144.850 162.010 144.990 162.890 ;
        RECT 137.860 161.870 144.990 162.010 ;
        RECT 137.860 161.810 138.180 161.870 ;
        RECT 17.270 161.190 146.990 161.670 ;
        RECT 35.280 160.990 35.600 161.050 ;
        RECT 37.135 160.990 37.425 161.035 ;
        RECT 35.280 160.850 37.425 160.990 ;
        RECT 35.280 160.790 35.600 160.850 ;
        RECT 37.135 160.805 37.425 160.850 ;
        RECT 35.740 160.650 36.060 160.710 ;
        RECT 36.215 160.650 36.505 160.695 ;
        RECT 35.740 160.510 36.505 160.650 ;
        RECT 37.210 160.650 37.350 160.805 ;
        RECT 47.700 160.790 48.020 161.050 ;
        RECT 57.375 160.990 57.665 161.035 ;
        RECT 60.580 160.990 60.900 161.050 ;
        RECT 57.375 160.850 60.900 160.990 ;
        RECT 57.375 160.805 57.665 160.850 ;
        RECT 60.580 160.790 60.900 160.850 ;
        RECT 63.340 160.990 63.660 161.050 ;
        RECT 65.180 160.990 65.500 161.050 ;
        RECT 65.655 160.990 65.945 161.035 ;
        RECT 63.340 160.850 65.945 160.990 ;
        RECT 63.340 160.790 63.660 160.850 ;
        RECT 65.180 160.790 65.500 160.850 ;
        RECT 65.655 160.805 65.945 160.850 ;
        RECT 56.440 160.650 56.760 160.710 ;
        RECT 37.210 160.510 56.760 160.650 ;
        RECT 35.740 160.450 36.060 160.510 ;
        RECT 36.215 160.465 36.505 160.510 ;
        RECT 56.440 160.450 56.760 160.510 ;
        RECT 59.240 160.650 59.530 160.695 ;
        RECT 61.340 160.650 61.630 160.695 ;
        RECT 62.910 160.650 63.200 160.695 ;
        RECT 59.240 160.510 63.200 160.650 ;
        RECT 59.240 160.465 59.530 160.510 ;
        RECT 61.340 160.465 61.630 160.510 ;
        RECT 62.910 160.465 63.200 160.510 ;
        RECT 38.960 160.310 39.280 160.370 ;
        RECT 35.830 160.170 41.030 160.310 ;
        RECT 32.520 159.970 32.840 160.030 ;
        RECT 35.830 160.015 35.970 160.170 ;
        RECT 38.960 160.110 39.280 160.170 ;
        RECT 35.755 159.970 36.045 160.015 ;
        RECT 38.500 159.970 38.820 160.030 ;
        RECT 40.890 160.015 41.030 160.170 ;
        RECT 58.740 160.110 59.060 160.370 ;
        RECT 59.635 160.310 59.925 160.355 ;
        RECT 60.825 160.310 61.115 160.355 ;
        RECT 63.345 160.310 63.635 160.355 ;
        RECT 59.635 160.170 63.635 160.310 ;
        RECT 65.730 160.310 65.870 160.805 ;
        RECT 70.700 160.790 71.020 161.050 ;
        RECT 85.420 160.790 85.740 161.050 ;
        RECT 88.180 160.990 88.500 161.050 ;
        RECT 89.115 160.990 89.405 161.035 ;
        RECT 94.160 160.990 94.480 161.050 ;
        RECT 101.060 160.990 101.380 161.050 ;
        RECT 88.180 160.850 89.405 160.990 ;
        RECT 88.180 160.790 88.500 160.850 ;
        RECT 89.115 160.805 89.405 160.850 ;
        RECT 90.570 160.850 105.890 160.990 ;
        RECT 74.880 160.650 75.170 160.695 ;
        RECT 76.980 160.650 77.270 160.695 ;
        RECT 78.550 160.650 78.840 160.695 ;
        RECT 74.880 160.510 78.840 160.650 ;
        RECT 74.880 160.465 75.170 160.510 ;
        RECT 76.980 160.465 77.270 160.510 ;
        RECT 78.550 160.465 78.840 160.510 ;
        RECT 70.240 160.310 70.560 160.370 ;
        RECT 73.460 160.310 73.780 160.370 ;
        RECT 90.570 160.355 90.710 160.850 ;
        RECT 94.160 160.790 94.480 160.850 ;
        RECT 101.060 160.790 101.380 160.850 ;
        RECT 90.980 160.650 91.270 160.695 ;
        RECT 93.080 160.650 93.370 160.695 ;
        RECT 94.650 160.650 94.940 160.695 ;
        RECT 90.980 160.510 94.940 160.650 ;
        RECT 90.980 160.465 91.270 160.510 ;
        RECT 93.080 160.465 93.370 160.510 ;
        RECT 94.650 160.465 94.940 160.510 ;
        RECT 97.380 160.450 97.700 160.710 ;
        RECT 101.520 160.650 101.810 160.695 ;
        RECT 103.090 160.650 103.380 160.695 ;
        RECT 105.190 160.650 105.480 160.695 ;
        RECT 101.520 160.510 105.480 160.650 ;
        RECT 101.520 160.465 101.810 160.510 ;
        RECT 103.090 160.465 103.380 160.510 ;
        RECT 105.190 160.465 105.480 160.510 ;
        RECT 105.750 160.355 105.890 160.850 ;
        RECT 107.960 160.790 108.280 161.050 ;
        RECT 115.780 160.990 116.100 161.050 ;
        RECT 118.540 160.990 118.860 161.050 ;
        RECT 115.780 160.850 118.860 160.990 ;
        RECT 115.780 160.790 116.100 160.850 ;
        RECT 118.540 160.790 118.860 160.850 ;
        RECT 127.740 160.790 128.060 161.050 ;
        RECT 132.340 160.990 132.660 161.050 ;
        RECT 138.780 160.990 139.100 161.050 ;
        RECT 132.340 160.850 139.100 160.990 ;
        RECT 132.340 160.790 132.660 160.850 ;
        RECT 138.780 160.790 139.100 160.850 ;
        RECT 140.620 160.790 140.940 161.050 ;
        RECT 109.800 160.650 110.120 160.710 ;
        RECT 116.700 160.650 117.020 160.710 ;
        RECT 109.800 160.510 110.490 160.650 ;
        RECT 109.800 160.450 110.120 160.510 ;
        RECT 110.350 160.355 110.490 160.510 ;
        RECT 110.810 160.510 117.020 160.650 ;
        RECT 118.630 160.650 118.770 160.790 ;
        RECT 123.155 160.650 123.445 160.695 ;
        RECT 126.360 160.650 126.680 160.710 ;
        RECT 118.630 160.510 126.680 160.650 ;
        RECT 110.810 160.370 110.950 160.510 ;
        RECT 116.700 160.450 117.020 160.510 ;
        RECT 123.155 160.465 123.445 160.510 ;
        RECT 126.360 160.450 126.680 160.510 ;
        RECT 134.220 160.650 134.510 160.695 ;
        RECT 136.320 160.650 136.610 160.695 ;
        RECT 137.890 160.650 138.180 160.695 ;
        RECT 134.220 160.510 138.180 160.650 ;
        RECT 134.220 160.465 134.510 160.510 ;
        RECT 136.320 160.465 136.610 160.510 ;
        RECT 137.890 160.465 138.180 160.510 ;
        RECT 74.395 160.310 74.685 160.355 ;
        RECT 65.730 160.170 69.090 160.310 ;
        RECT 59.635 160.125 59.925 160.170 ;
        RECT 60.825 160.125 61.115 160.170 ;
        RECT 63.345 160.125 63.635 160.170 ;
        RECT 40.355 159.970 40.645 160.015 ;
        RECT 32.520 159.830 36.045 159.970 ;
        RECT 32.520 159.770 32.840 159.830 ;
        RECT 35.755 159.785 36.045 159.830 ;
        RECT 36.290 159.830 38.820 159.970 ;
        RECT 33.440 159.630 33.760 159.690 ;
        RECT 34.835 159.630 35.125 159.675 ;
        RECT 36.290 159.630 36.430 159.830 ;
        RECT 38.500 159.770 38.820 159.830 ;
        RECT 39.510 159.830 40.645 159.970 ;
        RECT 39.510 159.690 39.650 159.830 ;
        RECT 40.355 159.785 40.645 159.830 ;
        RECT 40.815 159.785 41.105 160.015 ;
        RECT 33.440 159.490 36.430 159.630 ;
        RECT 33.440 159.430 33.760 159.490 ;
        RECT 34.835 159.445 35.125 159.490 ;
        RECT 38.040 159.430 38.360 159.690 ;
        RECT 38.975 159.630 39.265 159.675 ;
        RECT 39.420 159.630 39.740 159.690 ;
        RECT 38.975 159.490 39.740 159.630 ;
        RECT 38.975 159.445 39.265 159.490 ;
        RECT 39.420 159.430 39.740 159.490 ;
        RECT 39.895 159.630 40.185 159.675 ;
        RECT 40.890 159.630 41.030 159.785 ;
        RECT 41.720 159.770 42.040 160.030 ;
        RECT 54.615 159.970 54.905 160.015 ;
        RECT 55.060 159.970 55.380 160.030 ;
        RECT 54.615 159.830 55.380 159.970 ;
        RECT 54.615 159.785 54.905 159.830 ;
        RECT 55.060 159.770 55.380 159.830 ;
        RECT 55.535 159.970 55.825 160.015 ;
        RECT 55.980 159.970 56.300 160.030 ;
        RECT 64.260 159.970 64.580 160.030 ;
        RECT 55.535 159.830 56.300 159.970 ;
        RECT 57.755 159.845 64.580 159.970 ;
        RECT 55.535 159.785 55.825 159.830 ;
        RECT 55.980 159.770 56.300 159.830 ;
        RECT 57.605 159.830 64.580 159.845 ;
        RECT 39.895 159.490 41.030 159.630 ;
        RECT 46.780 159.630 47.100 159.690 ;
        RECT 46.780 159.490 54.830 159.630 ;
        RECT 39.895 159.445 40.185 159.490 ;
        RECT 46.780 159.430 47.100 159.490 ;
        RECT 54.690 159.350 54.830 159.490 ;
        RECT 56.440 159.430 56.760 159.690 ;
        RECT 57.605 159.615 57.895 159.830 ;
        RECT 64.260 159.770 64.580 159.830 ;
        RECT 64.720 159.970 65.040 160.030 ;
        RECT 67.035 159.970 67.325 160.015 ;
        RECT 64.720 159.830 67.325 159.970 ;
        RECT 64.720 159.770 65.040 159.830 ;
        RECT 67.035 159.785 67.325 159.830 ;
        RECT 67.940 159.770 68.260 160.030 ;
        RECT 68.400 159.770 68.720 160.030 ;
        RECT 68.950 160.015 69.090 160.170 ;
        RECT 70.240 160.170 74.685 160.310 ;
        RECT 70.240 160.110 70.560 160.170 ;
        RECT 73.460 160.110 73.780 160.170 ;
        RECT 74.395 160.125 74.685 160.170 ;
        RECT 75.275 160.310 75.565 160.355 ;
        RECT 76.465 160.310 76.755 160.355 ;
        RECT 78.985 160.310 79.275 160.355 ;
        RECT 75.275 160.170 79.275 160.310 ;
        RECT 75.275 160.125 75.565 160.170 ;
        RECT 76.465 160.125 76.755 160.170 ;
        RECT 78.985 160.125 79.275 160.170 ;
        RECT 82.675 160.310 82.965 160.355 ;
        RECT 82.675 160.170 87.030 160.310 ;
        RECT 82.675 160.125 82.965 160.170 ;
        RECT 68.875 159.785 69.165 160.015 ;
        RECT 69.795 159.785 70.085 160.015 ;
        RECT 59.980 159.630 60.270 159.675 ;
        RECT 58.370 159.490 60.270 159.630 ;
        RECT 33.900 159.090 34.220 159.350 ;
        RECT 37.055 159.290 37.345 159.335 ;
        RECT 38.515 159.290 38.805 159.335 ;
        RECT 37.055 159.150 38.805 159.290 ;
        RECT 37.055 159.105 37.345 159.150 ;
        RECT 38.515 159.105 38.805 159.150 ;
        RECT 42.655 159.290 42.945 159.335 ;
        RECT 46.320 159.290 46.640 159.350 ;
        RECT 42.655 159.150 46.640 159.290 ;
        RECT 42.655 159.105 42.945 159.150 ;
        RECT 46.320 159.090 46.640 159.150 ;
        RECT 47.240 159.290 47.560 159.350 ;
        RECT 47.795 159.290 48.085 159.335 ;
        RECT 47.240 159.150 48.085 159.290 ;
        RECT 47.240 159.090 47.560 159.150 ;
        RECT 47.795 159.105 48.085 159.150 ;
        RECT 48.635 159.290 48.925 159.335 ;
        RECT 50.460 159.290 50.780 159.350 ;
        RECT 48.635 159.150 50.780 159.290 ;
        RECT 48.635 159.105 48.925 159.150 ;
        RECT 50.460 159.090 50.780 159.150 ;
        RECT 54.600 159.090 54.920 159.350 ;
        RECT 55.075 159.290 55.365 159.335 ;
        RECT 56.900 159.290 57.220 159.350 ;
        RECT 58.370 159.335 58.510 159.490 ;
        RECT 59.980 159.445 60.270 159.490 ;
        RECT 61.040 159.630 61.360 159.690 ;
        RECT 66.115 159.630 66.405 159.675 ;
        RECT 61.040 159.490 66.405 159.630 ;
        RECT 61.040 159.430 61.360 159.490 ;
        RECT 66.115 159.445 66.405 159.490 ;
        RECT 66.560 159.630 66.880 159.690 ;
        RECT 69.870 159.630 70.010 159.785 ;
        RECT 73.920 159.770 74.240 160.030 ;
        RECT 75.760 160.015 76.080 160.030 ;
        RECT 75.730 159.970 76.080 160.015 ;
        RECT 75.565 159.830 76.080 159.970 ;
        RECT 75.730 159.785 76.080 159.830 ;
        RECT 75.760 159.770 76.080 159.785 ;
        RECT 82.200 159.770 82.520 160.030 ;
        RECT 83.120 159.770 83.440 160.030 ;
        RECT 86.340 159.770 86.660 160.030 ;
        RECT 86.890 160.015 87.030 160.170 ;
        RECT 90.440 160.125 90.730 160.355 ;
        RECT 91.375 160.310 91.665 160.355 ;
        RECT 92.565 160.310 92.855 160.355 ;
        RECT 95.085 160.310 95.375 160.355 ;
        RECT 91.375 160.170 95.375 160.310 ;
        RECT 91.375 160.125 91.665 160.170 ;
        RECT 92.565 160.125 92.855 160.170 ;
        RECT 95.085 160.125 95.375 160.170 ;
        RECT 101.085 160.310 101.375 160.355 ;
        RECT 103.605 160.310 103.895 160.355 ;
        RECT 104.795 160.310 105.085 160.355 ;
        RECT 101.085 160.170 105.085 160.310 ;
        RECT 101.085 160.125 101.375 160.170 ;
        RECT 103.605 160.125 103.895 160.170 ;
        RECT 104.795 160.125 105.085 160.170 ;
        RECT 105.675 160.125 105.965 160.355 ;
        RECT 110.275 160.125 110.565 160.355 ;
        RECT 110.720 160.110 111.040 160.370 ;
        RECT 112.560 160.310 112.880 160.370 ;
        RECT 111.730 160.170 112.880 160.310 ;
        RECT 86.815 159.785 87.105 160.015 ;
        RECT 89.100 159.970 89.420 160.030 ;
        RECT 89.575 159.970 89.865 160.015 ;
        RECT 89.100 159.830 89.865 159.970 ;
        RECT 89.100 159.770 89.420 159.830 ;
        RECT 89.575 159.785 89.865 159.830 ;
        RECT 90.035 159.970 90.325 160.015 ;
        RECT 90.940 159.970 91.260 160.030 ;
        RECT 97.840 159.970 98.160 160.030 ;
        RECT 90.035 159.830 98.160 159.970 ;
        RECT 90.035 159.785 90.325 159.830 ;
        RECT 66.560 159.490 70.010 159.630 ;
        RECT 78.980 159.630 79.300 159.690 ;
        RECT 85.435 159.630 85.725 159.675 ;
        RECT 78.980 159.490 85.725 159.630 ;
        RECT 66.560 159.430 66.880 159.490 ;
        RECT 78.980 159.430 79.300 159.490 ;
        RECT 85.435 159.445 85.725 159.490 ;
        RECT 55.075 159.150 57.220 159.290 ;
        RECT 55.075 159.105 55.365 159.150 ;
        RECT 56.900 159.090 57.220 159.150 ;
        RECT 58.295 159.105 58.585 159.335 ;
        RECT 60.580 159.290 60.900 159.350 ;
        RECT 68.875 159.290 69.165 159.335 ;
        RECT 60.580 159.150 69.165 159.290 ;
        RECT 60.580 159.090 60.900 159.150 ;
        RECT 68.875 159.105 69.165 159.150 ;
        RECT 78.520 159.290 78.840 159.350 ;
        RECT 81.295 159.290 81.585 159.335 ;
        RECT 78.520 159.150 81.585 159.290 ;
        RECT 78.520 159.090 78.840 159.150 ;
        RECT 81.295 159.105 81.585 159.150 ;
        RECT 88.180 159.090 88.500 159.350 ;
        RECT 89.650 159.290 89.790 159.785 ;
        RECT 90.940 159.770 91.260 159.830 ;
        RECT 97.840 159.770 98.160 159.830 ;
        RECT 109.815 159.970 110.105 160.015 ;
        RECT 111.730 159.970 111.870 160.170 ;
        RECT 112.560 160.110 112.880 160.170 ;
        RECT 124.060 160.310 124.380 160.370 ;
        RECT 125.455 160.310 125.745 160.355 ;
        RECT 124.060 160.170 125.745 160.310 ;
        RECT 124.060 160.110 124.380 160.170 ;
        RECT 125.455 160.125 125.745 160.170 ;
        RECT 125.900 160.110 126.220 160.370 ;
        RECT 126.835 160.310 127.125 160.355 ;
        RECT 130.960 160.310 131.280 160.370 ;
        RECT 126.835 160.170 131.280 160.310 ;
        RECT 126.835 160.125 127.125 160.170 ;
        RECT 130.960 160.110 131.280 160.170 ;
        RECT 133.720 160.110 134.040 160.370 ;
        RECT 134.615 160.310 134.905 160.355 ;
        RECT 135.805 160.310 136.095 160.355 ;
        RECT 138.325 160.310 138.615 160.355 ;
        RECT 134.615 160.170 138.615 160.310 ;
        RECT 134.615 160.125 134.905 160.170 ;
        RECT 135.805 160.125 136.095 160.170 ;
        RECT 138.325 160.125 138.615 160.170 ;
        RECT 143.380 160.110 143.700 160.370 ;
        RECT 143.840 160.110 144.160 160.370 ;
        RECT 109.815 159.830 111.870 159.970 ;
        RECT 109.815 159.785 110.105 159.830 ;
        RECT 112.100 159.770 112.420 160.030 ;
        RECT 113.035 159.970 113.325 160.015 ;
        RECT 115.320 159.970 115.640 160.030 ;
        RECT 113.035 159.830 115.640 159.970 ;
        RECT 113.035 159.785 113.325 159.830 ;
        RECT 115.320 159.770 115.640 159.830 ;
        RECT 119.015 159.970 119.305 160.015 ;
        RECT 119.460 159.970 119.780 160.030 ;
        RECT 119.015 159.830 119.780 159.970 ;
        RECT 119.015 159.785 119.305 159.830 ;
        RECT 119.460 159.770 119.780 159.830 ;
        RECT 119.935 159.970 120.225 160.015 ;
        RECT 121.760 159.970 122.080 160.030 ;
        RECT 122.695 159.970 122.985 160.015 ;
        RECT 119.935 159.830 122.985 159.970 ;
        RECT 119.935 159.785 120.225 159.830 ;
        RECT 121.760 159.770 122.080 159.830 ;
        RECT 122.695 159.785 122.985 159.830 ;
        RECT 91.830 159.630 92.120 159.675 ;
        RECT 92.780 159.630 93.100 159.690 ;
        RECT 91.830 159.490 93.100 159.630 ;
        RECT 91.830 159.445 92.120 159.490 ;
        RECT 92.780 159.430 93.100 159.490 ;
        RECT 104.280 159.675 104.600 159.690 ;
        RECT 104.280 159.445 104.630 159.675 ;
        RECT 108.420 159.630 108.740 159.690 ;
        RECT 112.575 159.630 112.865 159.675 ;
        RECT 108.420 159.490 112.865 159.630 ;
        RECT 122.770 159.630 122.910 159.785 ;
        RECT 126.360 159.770 126.680 160.030 ;
        RECT 127.740 159.970 128.060 160.030 ;
        RECT 128.215 159.970 128.505 160.015 ;
        RECT 127.740 159.830 128.505 159.970 ;
        RECT 127.740 159.770 128.060 159.830 ;
        RECT 128.215 159.785 128.505 159.830 ;
        RECT 129.135 159.970 129.425 160.015 ;
        RECT 129.580 159.970 129.900 160.030 ;
        RECT 131.420 159.970 131.740 160.030 ;
        RECT 135.100 160.015 135.420 160.030 ;
        RECT 135.070 159.970 135.420 160.015 ;
        RECT 129.135 159.830 131.740 159.970 ;
        RECT 134.905 159.830 135.420 159.970 ;
        RECT 129.135 159.785 129.425 159.830 ;
        RECT 129.580 159.770 129.900 159.830 ;
        RECT 131.420 159.770 131.740 159.830 ;
        RECT 135.070 159.785 135.420 159.830 ;
        RECT 135.100 159.770 135.420 159.785 ;
        RECT 125.440 159.630 125.760 159.690 ;
        RECT 126.450 159.630 126.590 159.770 ;
        RECT 128.675 159.630 128.965 159.675 ;
        RECT 122.770 159.490 126.130 159.630 ;
        RECT 126.450 159.490 128.965 159.630 ;
        RECT 104.280 159.430 104.600 159.445 ;
        RECT 108.420 159.430 108.740 159.490 ;
        RECT 112.575 159.445 112.865 159.490 ;
        RECT 125.440 159.430 125.760 159.490 ;
        RECT 96.000 159.290 96.320 159.350 ;
        RECT 89.650 159.150 96.320 159.290 ;
        RECT 96.000 159.090 96.320 159.150 ;
        RECT 97.380 159.290 97.700 159.350 ;
        RECT 98.775 159.290 99.065 159.335 ;
        RECT 97.380 159.150 99.065 159.290 ;
        RECT 97.380 159.090 97.700 159.150 ;
        RECT 98.775 159.105 99.065 159.150 ;
        RECT 117.160 159.290 117.480 159.350 ;
        RECT 119.475 159.290 119.765 159.335 ;
        RECT 117.160 159.150 119.765 159.290 ;
        RECT 117.160 159.090 117.480 159.150 ;
        RECT 119.475 159.105 119.765 159.150 ;
        RECT 122.680 159.290 123.000 159.350 ;
        RECT 124.060 159.290 124.380 159.350 ;
        RECT 122.680 159.150 124.380 159.290 ;
        RECT 125.990 159.290 126.130 159.490 ;
        RECT 128.675 159.445 128.965 159.490 ;
        RECT 127.740 159.290 128.060 159.350 ;
        RECT 125.990 159.150 128.060 159.290 ;
        RECT 122.680 159.090 123.000 159.150 ;
        RECT 124.060 159.090 124.380 159.150 ;
        RECT 127.740 159.090 128.060 159.150 ;
        RECT 141.080 159.090 141.400 159.350 ;
        RECT 142.920 159.090 143.240 159.350 ;
        RECT 17.270 158.470 146.990 158.950 ;
        RECT 15.840 158.270 16.260 158.410 ;
        RECT 74.380 158.270 74.700 158.330 ;
        RECT 76.695 158.270 76.985 158.315 ;
        RECT 15.840 158.130 73.920 158.270 ;
        RECT 15.840 157.960 16.260 158.130 ;
        RECT 31.155 157.930 31.445 157.975 ;
        RECT 32.075 157.930 32.365 157.975 ;
        RECT 31.155 157.790 32.365 157.930 ;
        RECT 31.155 157.745 31.445 157.790 ;
        RECT 32.075 157.745 32.365 157.790 ;
        RECT 33.155 157.930 33.445 157.975 ;
        RECT 33.900 157.930 34.220 157.990 ;
        RECT 33.155 157.790 34.220 157.930 ;
        RECT 33.155 157.745 33.445 157.790 ;
        RECT 33.900 157.730 34.220 157.790 ;
        RECT 45.415 157.930 45.705 157.975 ;
        RECT 47.240 157.930 47.560 157.990 ;
        RECT 45.415 157.790 47.560 157.930 ;
        RECT 45.415 157.745 45.705 157.790 ;
        RECT 47.240 157.730 47.560 157.790 ;
        RECT 47.700 157.930 48.020 157.990 ;
        RECT 54.600 157.930 54.920 157.990 ;
        RECT 55.075 157.930 55.365 157.975 ;
        RECT 47.700 157.790 53.910 157.930 ;
        RECT 47.700 157.730 48.020 157.790 ;
        RECT 29.300 157.590 29.620 157.650 ;
        RECT 30.695 157.590 30.985 157.635 ;
        RECT 29.300 157.450 30.985 157.590 ;
        RECT 29.300 157.390 29.620 157.450 ;
        RECT 30.695 157.405 30.985 157.450 ;
        RECT 31.615 157.590 31.905 157.635 ;
        RECT 32.520 157.590 32.840 157.650 ;
        RECT 31.615 157.450 32.840 157.590 ;
        RECT 31.615 157.405 31.905 157.450 ;
        RECT 30.770 157.250 30.910 157.405 ;
        RECT 32.520 157.390 32.840 157.450 ;
        RECT 34.375 157.590 34.665 157.635 ;
        RECT 34.820 157.590 35.140 157.650 ;
        RECT 35.740 157.635 36.060 157.650 ;
        RECT 35.710 157.590 36.060 157.635 ;
        RECT 34.375 157.450 35.140 157.590 ;
        RECT 35.545 157.450 36.060 157.590 ;
        RECT 34.375 157.405 34.665 157.450 ;
        RECT 34.820 157.390 35.140 157.450 ;
        RECT 35.710 157.405 36.060 157.450 ;
        RECT 35.740 157.390 36.060 157.405 ;
        RECT 46.320 157.390 46.640 157.650 ;
        RECT 46.780 157.390 47.100 157.650 ;
        RECT 48.175 157.590 48.465 157.635 ;
        RECT 47.330 157.450 48.465 157.590 ;
        RECT 33.440 157.250 33.760 157.310 ;
        RECT 30.770 157.110 33.760 157.250 ;
        RECT 33.440 157.050 33.760 157.110 ;
        RECT 35.255 157.250 35.545 157.295 ;
        RECT 36.445 157.250 36.735 157.295 ;
        RECT 38.965 157.250 39.255 157.295 ;
        RECT 35.255 157.110 39.255 157.250 ;
        RECT 35.255 157.065 35.545 157.110 ;
        RECT 36.445 157.065 36.735 157.110 ;
        RECT 38.965 157.065 39.255 157.110 ;
        RECT 34.360 156.910 34.680 156.970 ;
        RECT 33.070 156.770 34.680 156.910 ;
        RECT 33.070 156.615 33.210 156.770 ;
        RECT 34.360 156.710 34.680 156.770 ;
        RECT 34.860 156.910 35.150 156.955 ;
        RECT 36.960 156.910 37.250 156.955 ;
        RECT 38.530 156.910 38.820 156.955 ;
        RECT 34.860 156.770 38.820 156.910 ;
        RECT 47.330 156.910 47.470 157.450 ;
        RECT 48.175 157.405 48.465 157.450 ;
        RECT 50.000 157.390 50.320 157.650 ;
        RECT 50.460 157.590 50.780 157.650 ;
        RECT 50.460 157.450 50.975 157.590 ;
        RECT 50.460 157.390 50.780 157.450 ;
        RECT 51.380 157.390 51.700 157.650 ;
        RECT 52.300 157.635 52.620 157.650 ;
        RECT 53.770 157.635 53.910 157.790 ;
        RECT 54.600 157.790 55.365 157.930 ;
        RECT 54.600 157.730 54.920 157.790 ;
        RECT 55.075 157.745 55.365 157.790 ;
        RECT 55.980 157.930 56.300 157.990 ;
        RECT 61.500 157.930 61.820 157.990 ;
        RECT 62.435 157.930 62.725 157.975 ;
        RECT 55.980 157.790 62.725 157.930 ;
        RECT 55.980 157.730 56.300 157.790 ;
        RECT 61.500 157.730 61.820 157.790 ;
        RECT 62.435 157.745 62.725 157.790 ;
        RECT 64.260 157.730 64.580 157.990 ;
        RECT 65.180 157.730 65.500 157.990 ;
        RECT 66.115 157.930 66.405 157.975 ;
        RECT 66.560 157.930 66.880 157.990 ;
        RECT 66.115 157.790 66.880 157.930 ;
        RECT 66.115 157.745 66.405 157.790 ;
        RECT 66.560 157.730 66.880 157.790 ;
        RECT 71.130 157.930 71.420 157.975 ;
        RECT 71.620 157.930 71.940 157.990 ;
        RECT 71.130 157.790 71.940 157.930 ;
        RECT 73.780 157.930 73.920 158.130 ;
        RECT 74.380 158.130 76.985 158.270 ;
        RECT 74.380 158.070 74.700 158.130 ;
        RECT 76.695 158.085 76.985 158.130 ;
        RECT 92.780 158.070 93.100 158.330 ;
        RECT 95.540 158.270 95.860 158.330 ;
        RECT 99.235 158.270 99.525 158.315 ;
        RECT 95.540 158.130 99.525 158.270 ;
        RECT 95.540 158.070 95.860 158.130 ;
        RECT 99.235 158.085 99.525 158.130 ;
        RECT 104.280 158.270 104.600 158.330 ;
        RECT 104.755 158.270 105.045 158.315 ;
        RECT 104.280 158.130 105.045 158.270 ;
        RECT 104.280 158.070 104.600 158.130 ;
        RECT 104.755 158.085 105.045 158.130 ;
        RECT 114.860 158.270 115.180 158.330 ;
        RECT 123.140 158.270 123.460 158.330 ;
        RECT 129.580 158.270 129.900 158.330 ;
        RECT 114.860 158.130 123.460 158.270 ;
        RECT 114.860 158.070 115.180 158.130 ;
        RECT 123.140 158.070 123.460 158.130 ;
        RECT 126.910 158.130 129.900 158.270 ;
        RECT 80.375 157.930 80.665 157.975 ;
        RECT 73.780 157.790 80.665 157.930 ;
        RECT 71.130 157.745 71.420 157.790 ;
        RECT 71.620 157.730 71.940 157.790 ;
        RECT 80.375 157.745 80.665 157.790 ;
        RECT 101.535 157.930 101.825 157.975 ;
        RECT 107.960 157.930 108.280 157.990 ;
        RECT 126.910 157.975 127.050 158.130 ;
        RECT 129.580 158.070 129.900 158.130 ;
        RECT 131.895 158.270 132.185 158.315 ;
        RECT 136.480 158.270 136.800 158.330 ;
        RECT 131.895 158.130 136.800 158.270 ;
        RECT 131.895 158.085 132.185 158.130 ;
        RECT 136.480 158.070 136.800 158.130 ;
        RECT 113.955 157.930 114.245 157.975 ;
        RECT 101.535 157.790 110.950 157.930 ;
        RECT 101.535 157.745 101.825 157.790 ;
        RECT 107.960 157.730 108.280 157.790 ;
        RECT 51.855 157.405 52.145 157.635 ;
        RECT 52.300 157.590 52.630 157.635 ;
        RECT 52.300 157.450 52.815 157.590 ;
        RECT 52.300 157.405 52.630 157.450 ;
        RECT 53.695 157.405 53.985 157.635 ;
        RECT 47.715 157.250 48.005 157.295 ;
        RECT 50.920 157.250 51.240 157.310 ;
        RECT 47.715 157.110 51.240 157.250 ;
        RECT 47.715 157.065 48.005 157.110 ;
        RECT 50.920 157.050 51.240 157.110 ;
        RECT 51.930 157.250 52.070 157.405 ;
        RECT 52.300 157.390 52.620 157.405 ;
        RECT 54.140 157.390 54.460 157.650 ;
        RECT 56.440 157.390 56.760 157.650 ;
        RECT 56.900 157.590 57.220 157.650 ;
        RECT 56.900 157.450 57.415 157.590 ;
        RECT 56.900 157.390 57.220 157.450 ;
        RECT 57.835 157.405 58.125 157.635 ;
        RECT 52.760 157.250 53.080 157.310 ;
        RECT 57.910 157.250 58.050 157.405 ;
        RECT 58.280 157.390 58.600 157.650 ;
        RECT 58.985 157.590 59.275 157.635 ;
        RECT 60.580 157.590 60.900 157.650 ;
        RECT 58.985 157.450 60.900 157.590 ;
        RECT 58.985 157.405 59.275 157.450 ;
        RECT 60.580 157.390 60.900 157.450 ;
        RECT 61.040 157.390 61.360 157.650 ;
        RECT 61.975 157.405 62.265 157.635 ;
        RECT 62.050 157.250 62.190 157.405 ;
        RECT 62.880 157.390 63.200 157.650 ;
        RECT 69.795 157.590 70.085 157.635 ;
        RECT 70.240 157.590 70.560 157.650 ;
        RECT 69.795 157.450 70.560 157.590 ;
        RECT 69.795 157.405 70.085 157.450 ;
        RECT 70.240 157.390 70.560 157.450 ;
        RECT 96.935 157.590 97.225 157.635 ;
        RECT 98.300 157.590 98.620 157.650 ;
        RECT 96.935 157.450 98.620 157.590 ;
        RECT 96.935 157.405 97.225 157.450 ;
        RECT 98.300 157.390 98.620 157.450 ;
        RECT 101.060 157.390 101.380 157.650 ;
        RECT 102.900 157.590 103.220 157.650 ;
        RECT 104.295 157.590 104.585 157.635 ;
        RECT 102.900 157.450 104.585 157.590 ;
        RECT 102.900 157.390 103.220 157.450 ;
        RECT 104.295 157.405 104.585 157.450 ;
        RECT 106.120 157.590 106.440 157.650 ;
        RECT 110.810 157.635 110.950 157.790 ;
        RECT 113.955 157.790 116.930 157.930 ;
        RECT 113.955 157.745 114.245 157.790 ;
        RECT 106.595 157.590 106.885 157.635 ;
        RECT 106.120 157.450 106.885 157.590 ;
        RECT 106.120 157.390 106.440 157.450 ;
        RECT 106.595 157.405 106.885 157.450 ;
        RECT 110.735 157.405 111.025 157.635 ;
        RECT 114.415 157.590 114.705 157.635 ;
        RECT 115.320 157.590 115.640 157.650 ;
        RECT 114.415 157.450 115.640 157.590 ;
        RECT 114.415 157.405 114.705 157.450 ;
        RECT 115.320 157.390 115.640 157.450 ;
        RECT 64.720 157.250 65.040 157.310 ;
        RECT 51.930 157.110 53.080 157.250 ;
        RECT 51.930 156.910 52.070 157.110 ;
        RECT 52.760 157.050 53.080 157.110 ;
        RECT 54.690 157.110 58.050 157.250 ;
        RECT 59.750 157.110 62.190 157.250 ;
        RECT 62.510 157.110 65.040 157.250 ;
        RECT 47.330 156.770 52.070 156.910 ;
        RECT 53.235 156.910 53.525 156.955 ;
        RECT 54.690 156.910 54.830 157.110 ;
        RECT 53.235 156.770 54.830 156.910 ;
        RECT 34.860 156.725 35.150 156.770 ;
        RECT 36.960 156.725 37.250 156.770 ;
        RECT 38.530 156.725 38.820 156.770 ;
        RECT 53.235 156.725 53.525 156.770 ;
        RECT 55.060 156.710 55.380 156.970 ;
        RECT 59.750 156.955 59.890 157.110 ;
        RECT 59.675 156.725 59.965 156.955 ;
        RECT 60.580 156.910 60.900 156.970 ;
        RECT 62.510 156.910 62.650 157.110 ;
        RECT 64.720 157.050 65.040 157.110 ;
        RECT 70.675 157.250 70.965 157.295 ;
        RECT 71.865 157.250 72.155 157.295 ;
        RECT 74.385 157.250 74.675 157.295 ;
        RECT 70.675 157.110 74.675 157.250 ;
        RECT 70.675 157.065 70.965 157.110 ;
        RECT 71.865 157.065 72.155 157.110 ;
        RECT 74.385 157.065 74.675 157.110 ;
        RECT 87.260 157.250 87.580 157.310 ;
        RECT 89.575 157.250 89.865 157.295 ;
        RECT 87.260 157.110 89.865 157.250 ;
        RECT 87.260 157.050 87.580 157.110 ;
        RECT 89.575 157.065 89.865 157.110 ;
        RECT 97.380 157.050 97.700 157.310 ;
        RECT 97.840 157.250 98.160 157.310 ;
        RECT 101.995 157.250 102.285 157.295 ;
        RECT 97.840 157.110 102.285 157.250 ;
        RECT 97.840 157.050 98.160 157.110 ;
        RECT 101.995 157.065 102.285 157.110 ;
        RECT 107.055 157.065 107.345 157.295 ;
        RECT 107.975 157.250 108.265 157.295 ;
        RECT 108.420 157.250 108.740 157.310 ;
        RECT 107.975 157.110 108.740 157.250 ;
        RECT 107.975 157.065 108.265 157.110 ;
        RECT 60.580 156.770 62.650 156.910 ;
        RECT 63.815 156.910 64.105 156.955 ;
        RECT 67.480 156.910 67.800 156.970 ;
        RECT 63.815 156.770 67.800 156.910 ;
        RECT 60.580 156.710 60.900 156.770 ;
        RECT 63.815 156.725 64.105 156.770 ;
        RECT 67.480 156.710 67.800 156.770 ;
        RECT 70.280 156.910 70.570 156.955 ;
        RECT 72.380 156.910 72.670 156.955 ;
        RECT 73.950 156.910 74.240 156.955 ;
        RECT 70.280 156.770 74.240 156.910 ;
        RECT 70.280 156.725 70.570 156.770 ;
        RECT 72.380 156.725 72.670 156.770 ;
        RECT 73.950 156.725 74.240 156.770 ;
        RECT 95.095 156.910 95.385 156.955 ;
        RECT 96.460 156.910 96.780 156.970 ;
        RECT 95.095 156.770 96.780 156.910 ;
        RECT 107.130 156.910 107.270 157.065 ;
        RECT 108.420 157.050 108.740 157.110 ;
        RECT 114.860 157.050 115.180 157.310 ;
        RECT 115.795 157.065 116.085 157.295 ;
        RECT 116.255 157.250 116.545 157.295 ;
        RECT 116.790 157.250 116.930 157.790 ;
        RECT 117.250 157.790 121.070 157.930 ;
        RECT 117.250 157.650 117.390 157.790 ;
        RECT 117.160 157.390 117.480 157.650 ;
        RECT 117.635 157.590 117.925 157.635 ;
        RECT 118.080 157.590 118.400 157.650 ;
        RECT 117.635 157.450 118.400 157.590 ;
        RECT 117.635 157.405 117.925 157.450 ;
        RECT 118.080 157.390 118.400 157.450 ;
        RECT 118.540 157.590 118.860 157.650 ;
        RECT 120.380 157.590 120.700 157.650 ;
        RECT 118.540 157.450 120.700 157.590 ;
        RECT 120.930 157.590 121.070 157.790 ;
        RECT 126.835 157.745 127.125 157.975 ;
        RECT 130.515 157.930 130.805 157.975 ;
        RECT 131.420 157.930 131.740 157.990 ;
        RECT 130.515 157.790 131.740 157.930 ;
        RECT 130.515 157.745 130.805 157.790 ;
        RECT 131.420 157.730 131.740 157.790 ;
        RECT 135.530 157.930 135.820 157.975 ;
        RECT 141.080 157.930 141.400 157.990 ;
        RECT 135.530 157.790 141.400 157.930 ;
        RECT 135.530 157.745 135.820 157.790 ;
        RECT 141.080 157.730 141.400 157.790 ;
        RECT 120.930 157.580 121.990 157.590 ;
        RECT 122.695 157.580 122.985 157.635 ;
        RECT 120.930 157.450 122.985 157.580 ;
        RECT 118.540 157.390 118.860 157.450 ;
        RECT 120.380 157.390 120.700 157.450 ;
        RECT 121.850 157.440 122.985 157.450 ;
        RECT 122.695 157.405 122.985 157.440 ;
        RECT 123.155 157.580 123.445 157.635 ;
        RECT 124.060 157.590 124.380 157.650 ;
        RECT 124.535 157.590 124.825 157.635 ;
        RECT 123.690 157.580 124.825 157.590 ;
        RECT 123.155 157.450 124.825 157.580 ;
        RECT 123.155 157.440 123.830 157.450 ;
        RECT 123.155 157.405 123.445 157.440 ;
        RECT 124.060 157.390 124.380 157.450 ;
        RECT 124.535 157.405 124.825 157.450 ;
        RECT 125.440 157.390 125.760 157.650 ;
        RECT 127.755 157.590 128.045 157.635 ;
        RECT 128.200 157.590 128.520 157.650 ;
        RECT 127.755 157.450 128.520 157.590 ;
        RECT 127.755 157.405 128.045 157.450 ;
        RECT 128.200 157.390 128.520 157.450 ;
        RECT 129.135 157.590 129.425 157.635 ;
        RECT 129.580 157.590 129.900 157.650 ;
        RECT 129.135 157.450 129.900 157.590 ;
        RECT 129.135 157.405 129.425 157.450 ;
        RECT 129.580 157.390 129.900 157.450 ;
        RECT 130.040 157.390 130.360 157.650 ;
        RECT 130.975 157.590 131.265 157.635 ;
        RECT 133.260 157.590 133.580 157.650 ;
        RECT 130.975 157.450 133.580 157.590 ;
        RECT 130.975 157.405 131.265 157.450 ;
        RECT 133.260 157.390 133.580 157.450 ;
        RECT 133.720 157.590 134.040 157.650 ;
        RECT 134.195 157.590 134.485 157.635 ;
        RECT 143.395 157.590 143.685 157.635 ;
        RECT 133.720 157.450 134.485 157.590 ;
        RECT 133.720 157.390 134.040 157.450 ;
        RECT 134.195 157.405 134.485 157.450 ;
        RECT 134.685 157.450 143.685 157.590 ;
        RECT 116.255 157.110 116.930 157.250 ;
        RECT 116.255 157.065 116.545 157.110 ;
        RECT 115.870 156.910 116.010 157.065 ;
        RECT 119.460 157.050 119.780 157.310 ;
        RECT 121.775 157.065 122.065 157.295 ;
        RECT 122.235 157.250 122.525 157.295 ;
        RECT 125.900 157.250 126.220 157.310 ;
        RECT 122.235 157.110 126.220 157.250 ;
        RECT 122.235 157.065 122.525 157.110 ;
        RECT 116.715 156.910 117.005 156.955 ;
        RECT 107.130 156.770 115.090 156.910 ;
        RECT 115.870 156.770 117.005 156.910 ;
        RECT 95.095 156.725 95.385 156.770 ;
        RECT 96.460 156.710 96.780 156.770 ;
        RECT 114.950 156.630 115.090 156.770 ;
        RECT 116.715 156.725 117.005 156.770 ;
        RECT 117.160 156.910 117.480 156.970 ;
        RECT 119.015 156.910 119.305 156.955 ;
        RECT 117.160 156.770 119.305 156.910 ;
        RECT 121.850 156.910 121.990 157.065 ;
        RECT 125.900 157.050 126.220 157.110 ;
        RECT 127.280 157.250 127.600 157.310 ;
        RECT 134.685 157.250 134.825 157.450 ;
        RECT 143.395 157.405 143.685 157.450 ;
        RECT 127.280 157.110 134.825 157.250 ;
        RECT 135.075 157.250 135.365 157.295 ;
        RECT 136.265 157.250 136.555 157.295 ;
        RECT 138.785 157.250 139.075 157.295 ;
        RECT 135.075 157.110 139.075 157.250 ;
        RECT 127.280 157.050 127.600 157.110 ;
        RECT 135.075 157.065 135.365 157.110 ;
        RECT 136.265 157.065 136.555 157.110 ;
        RECT 138.785 157.065 139.075 157.110 ;
        RECT 143.840 157.050 144.160 157.310 ;
        RECT 144.760 157.050 145.080 157.310 ;
        RECT 122.680 156.910 123.000 156.970 ;
        RECT 124.995 156.910 125.285 156.955 ;
        RECT 121.850 156.770 122.450 156.910 ;
        RECT 117.160 156.710 117.480 156.770 ;
        RECT 119.015 156.725 119.305 156.770 ;
        RECT 122.310 156.630 122.450 156.770 ;
        RECT 122.680 156.770 125.285 156.910 ;
        RECT 122.680 156.710 123.000 156.770 ;
        RECT 124.995 156.725 125.285 156.770 ;
        RECT 134.680 156.910 134.970 156.955 ;
        RECT 136.780 156.910 137.070 156.955 ;
        RECT 138.350 156.910 138.640 156.955 ;
        RECT 134.680 156.770 138.640 156.910 ;
        RECT 134.680 156.725 134.970 156.770 ;
        RECT 136.780 156.725 137.070 156.770 ;
        RECT 138.350 156.725 138.640 156.770 ;
        RECT 32.995 156.385 33.285 156.615 ;
        RECT 33.915 156.570 34.205 156.615 ;
        RECT 36.200 156.570 36.520 156.630 ;
        RECT 33.915 156.430 36.520 156.570 ;
        RECT 33.915 156.385 34.205 156.430 ;
        RECT 36.200 156.370 36.520 156.430 ;
        RECT 39.880 156.570 40.200 156.630 ;
        RECT 41.275 156.570 41.565 156.615 ;
        RECT 39.880 156.430 41.565 156.570 ;
        RECT 39.880 156.370 40.200 156.430 ;
        RECT 41.275 156.385 41.565 156.430 ;
        RECT 50.000 156.570 50.320 156.630 ;
        RECT 54.600 156.570 54.920 156.630 ;
        RECT 50.000 156.430 54.920 156.570 ;
        RECT 50.000 156.370 50.320 156.430 ;
        RECT 54.600 156.370 54.920 156.430 ;
        RECT 58.740 156.570 59.060 156.630 ;
        RECT 69.320 156.570 69.640 156.630 ;
        RECT 58.740 156.430 69.640 156.570 ;
        RECT 58.740 156.370 59.060 156.430 ;
        RECT 69.320 156.370 69.640 156.430 ;
        RECT 86.800 156.370 87.120 156.630 ;
        RECT 103.820 156.370 104.140 156.630 ;
        RECT 114.860 156.370 115.180 156.630 ;
        RECT 115.320 156.370 115.640 156.630 ;
        RECT 115.780 156.570 116.100 156.630 ;
        RECT 118.080 156.570 118.400 156.630 ;
        RECT 115.780 156.430 118.400 156.570 ;
        RECT 115.780 156.370 116.100 156.430 ;
        RECT 118.080 156.370 118.400 156.430 ;
        RECT 122.220 156.370 122.540 156.630 ;
        RECT 124.060 156.370 124.380 156.630 ;
        RECT 128.675 156.570 128.965 156.615 ;
        RECT 130.040 156.570 130.360 156.630 ;
        RECT 128.675 156.430 130.360 156.570 ;
        RECT 128.675 156.385 128.965 156.430 ;
        RECT 130.040 156.370 130.360 156.430 ;
        RECT 137.400 156.570 137.720 156.630 ;
        RECT 141.095 156.570 141.385 156.615 ;
        RECT 137.400 156.430 141.385 156.570 ;
        RECT 137.400 156.370 137.720 156.430 ;
        RECT 141.095 156.385 141.385 156.430 ;
        RECT 141.540 156.370 141.860 156.630 ;
        RECT 17.270 155.750 146.990 156.230 ;
        RECT 31.155 155.550 31.445 155.595 ;
        RECT 32.060 155.550 32.380 155.610 ;
        RECT 31.155 155.410 32.380 155.550 ;
        RECT 31.155 155.365 31.445 155.410 ;
        RECT 32.060 155.350 32.380 155.410 ;
        RECT 44.955 155.550 45.245 155.595 ;
        RECT 51.380 155.550 51.700 155.610 ;
        RECT 44.955 155.410 51.700 155.550 ;
        RECT 44.955 155.365 45.245 155.410 ;
        RECT 51.380 155.350 51.700 155.410 ;
        RECT 61.515 155.550 61.805 155.595 ;
        RECT 62.895 155.550 63.185 155.595 ;
        RECT 61.515 155.410 63.185 155.550 ;
        RECT 61.515 155.365 61.805 155.410 ;
        RECT 62.895 155.365 63.185 155.410 ;
        RECT 87.260 155.350 87.580 155.610 ;
        RECT 106.120 155.350 106.440 155.610 ;
        RECT 107.960 155.350 108.280 155.610 ;
        RECT 111.640 155.550 111.960 155.610 ;
        RECT 115.335 155.550 115.625 155.595 ;
        RECT 111.640 155.410 115.625 155.550 ;
        RECT 111.640 155.350 111.960 155.410 ;
        RECT 115.335 155.365 115.625 155.410 ;
        RECT 119.460 155.550 119.780 155.610 ;
        RECT 123.615 155.550 123.905 155.595 ;
        RECT 142.920 155.550 143.240 155.610 ;
        RECT 145.235 155.550 145.525 155.595 ;
        RECT 119.460 155.410 123.905 155.550 ;
        RECT 119.460 155.350 119.780 155.410 ;
        RECT 123.615 155.365 123.905 155.410 ;
        RECT 132.430 155.410 139.010 155.550 ;
        RECT 33.900 155.210 34.190 155.255 ;
        RECT 35.470 155.210 35.760 155.255 ;
        RECT 37.570 155.210 37.860 155.255 ;
        RECT 33.900 155.070 37.860 155.210 ;
        RECT 33.900 155.025 34.190 155.070 ;
        RECT 35.470 155.025 35.760 155.070 ;
        RECT 37.570 155.025 37.860 155.070 ;
        RECT 38.040 155.010 38.360 155.270 ;
        RECT 47.700 155.010 48.020 155.270 ;
        RECT 58.280 155.210 58.600 155.270 ;
        RECT 57.910 155.070 58.600 155.210 ;
        RECT 33.465 154.870 33.755 154.915 ;
        RECT 35.985 154.870 36.275 154.915 ;
        RECT 37.175 154.870 37.465 154.915 ;
        RECT 33.465 154.730 37.465 154.870 ;
        RECT 38.130 154.870 38.270 155.010 ;
        RECT 38.130 154.730 44.250 154.870 ;
        RECT 33.465 154.685 33.755 154.730 ;
        RECT 35.985 154.685 36.275 154.730 ;
        RECT 37.175 154.685 37.465 154.730 ;
        RECT 34.820 154.530 35.140 154.590 ;
        RECT 38.055 154.530 38.345 154.575 ;
        RECT 34.820 154.390 38.345 154.530 ;
        RECT 34.820 154.330 35.140 154.390 ;
        RECT 38.055 154.345 38.345 154.390 ;
        RECT 38.500 154.330 38.820 154.590 ;
        RECT 38.960 154.530 39.280 154.590 ;
        RECT 39.435 154.530 39.725 154.575 ;
        RECT 38.960 154.390 39.725 154.530 ;
        RECT 38.960 154.330 39.280 154.390 ;
        RECT 39.435 154.345 39.725 154.390 ;
        RECT 39.880 154.330 40.200 154.590 ;
        RECT 40.355 154.345 40.645 154.575 ;
        RECT 40.800 154.530 41.120 154.590 ;
        RECT 40.800 154.390 41.950 154.530 ;
        RECT 36.200 154.190 36.520 154.250 ;
        RECT 36.720 154.190 37.010 154.235 ;
        RECT 36.200 154.050 37.010 154.190 ;
        RECT 38.590 154.190 38.730 154.330 ;
        RECT 40.430 154.190 40.570 154.345 ;
        RECT 40.800 154.330 41.120 154.390 ;
        RECT 38.590 154.050 40.570 154.190 ;
        RECT 41.810 154.190 41.950 154.390 ;
        RECT 42.180 154.330 42.500 154.590 ;
        RECT 42.640 154.330 42.960 154.590 ;
        RECT 44.110 154.575 44.250 154.730 ;
        RECT 43.575 154.345 43.865 154.575 ;
        RECT 44.035 154.345 44.325 154.575 ;
        RECT 45.415 154.345 45.705 154.575 ;
        RECT 43.650 154.190 43.790 154.345 ;
        RECT 45.490 154.190 45.630 154.345 ;
        RECT 46.780 154.330 47.100 154.590 ;
        RECT 57.910 154.575 58.050 155.070 ;
        RECT 58.280 155.010 58.600 155.070 ;
        RECT 59.215 155.210 59.505 155.255 ;
        RECT 59.675 155.210 59.965 155.255 ;
        RECT 66.560 155.210 66.880 155.270 ;
        RECT 59.215 155.070 66.880 155.210 ;
        RECT 59.215 155.025 59.505 155.070 ;
        RECT 59.675 155.025 59.965 155.070 ;
        RECT 66.560 155.010 66.880 155.070 ;
        RECT 90.020 155.210 90.310 155.255 ;
        RECT 91.590 155.210 91.880 155.255 ;
        RECT 93.690 155.210 93.980 155.255 ;
        RECT 90.020 155.070 93.980 155.210 ;
        RECT 90.020 155.025 90.310 155.070 ;
        RECT 91.590 155.025 91.880 155.070 ;
        RECT 93.690 155.025 93.980 155.070 ;
        RECT 95.120 155.210 95.410 155.255 ;
        RECT 97.220 155.210 97.510 155.255 ;
        RECT 98.790 155.210 99.080 155.255 ;
        RECT 95.120 155.070 99.080 155.210 ;
        RECT 95.120 155.025 95.410 155.070 ;
        RECT 97.220 155.025 97.510 155.070 ;
        RECT 98.790 155.025 99.080 155.070 ;
        RECT 110.720 155.210 111.010 155.255 ;
        RECT 112.290 155.210 112.580 155.255 ;
        RECT 114.390 155.210 114.680 155.255 ;
        RECT 110.720 155.070 114.680 155.210 ;
        RECT 110.720 155.025 111.010 155.070 ;
        RECT 112.290 155.025 112.580 155.070 ;
        RECT 114.390 155.025 114.680 155.070 ;
        RECT 114.860 155.210 115.180 155.270 ;
        RECT 120.840 155.210 121.160 155.270 ;
        RECT 114.860 155.070 121.160 155.210 ;
        RECT 114.860 155.010 115.180 155.070 ;
        RECT 120.840 155.010 121.160 155.070 ;
        RECT 124.060 155.210 124.380 155.270 ;
        RECT 124.060 155.070 127.970 155.210 ;
        RECT 124.060 155.010 124.380 155.070 ;
        RECT 60.580 154.870 60.900 154.930 ;
        RECT 89.585 154.870 89.875 154.915 ;
        RECT 92.105 154.870 92.395 154.915 ;
        RECT 93.295 154.870 93.585 154.915 ;
        RECT 58.370 154.730 64.950 154.870 ;
        RECT 58.370 154.575 58.510 154.730 ;
        RECT 60.580 154.670 60.900 154.730 ;
        RECT 57.835 154.345 58.125 154.575 ;
        RECT 58.295 154.345 58.585 154.575 ;
        RECT 41.810 154.050 45.630 154.190 ;
        RECT 57.910 154.190 58.050 154.345 ;
        RECT 64.810 154.250 64.950 154.730 ;
        RECT 89.585 154.730 93.585 154.870 ;
        RECT 89.585 154.685 89.875 154.730 ;
        RECT 92.105 154.685 92.395 154.730 ;
        RECT 93.295 154.685 93.585 154.730 ;
        RECT 94.160 154.870 94.480 154.930 ;
        RECT 94.635 154.870 94.925 154.915 ;
        RECT 94.160 154.730 94.925 154.870 ;
        RECT 94.160 154.670 94.480 154.730 ;
        RECT 94.635 154.685 94.925 154.730 ;
        RECT 95.515 154.870 95.805 154.915 ;
        RECT 96.705 154.870 96.995 154.915 ;
        RECT 99.225 154.870 99.515 154.915 ;
        RECT 95.515 154.730 99.515 154.870 ;
        RECT 95.515 154.685 95.805 154.730 ;
        RECT 96.705 154.685 96.995 154.730 ;
        RECT 99.225 154.685 99.515 154.730 ;
        RECT 110.285 154.870 110.575 154.915 ;
        RECT 112.805 154.870 113.095 154.915 ;
        RECT 113.995 154.870 114.285 154.915 ;
        RECT 110.285 154.730 114.285 154.870 ;
        RECT 110.285 154.685 110.575 154.730 ;
        RECT 112.805 154.685 113.095 154.730 ;
        RECT 113.995 154.685 114.285 154.730 ;
        RECT 116.700 154.870 117.020 154.930 ;
        RECT 118.095 154.870 118.385 154.915 ;
        RECT 116.700 154.730 118.385 154.870 ;
        RECT 116.700 154.670 117.020 154.730 ;
        RECT 118.095 154.685 118.385 154.730 ;
        RECT 122.695 154.870 122.985 154.915 ;
        RECT 123.155 154.870 123.445 154.915 ;
        RECT 126.360 154.870 126.680 154.930 ;
        RECT 127.830 154.915 127.970 155.070 ;
        RECT 122.695 154.730 123.445 154.870 ;
        RECT 122.695 154.685 122.985 154.730 ;
        RECT 123.155 154.685 123.445 154.730 ;
        RECT 124.150 154.730 126.680 154.870 ;
        RECT 73.920 154.530 74.240 154.590 ;
        RECT 78.535 154.530 78.825 154.575 ;
        RECT 78.980 154.530 79.300 154.590 ;
        RECT 73.920 154.390 79.300 154.530 ;
        RECT 73.920 154.330 74.240 154.390 ;
        RECT 78.535 154.345 78.825 154.390 ;
        RECT 78.980 154.330 79.300 154.390 ;
        RECT 79.900 154.330 80.220 154.590 ;
        RECT 97.380 154.530 97.700 154.590 ;
        RECT 102.915 154.530 103.205 154.575 ;
        RECT 97.380 154.390 103.205 154.530 ;
        RECT 97.380 154.330 97.700 154.390 ;
        RECT 102.915 154.345 103.205 154.390 ;
        RECT 112.100 154.530 112.420 154.590 ;
        RECT 114.875 154.530 115.165 154.575 ;
        RECT 112.100 154.390 115.165 154.530 ;
        RECT 112.100 154.330 112.420 154.390 ;
        RECT 114.875 154.345 115.165 154.390 ;
        RECT 115.320 154.330 115.640 154.590 ;
        RECT 117.635 154.530 117.925 154.575 ;
        RECT 119.000 154.530 119.320 154.590 ;
        RECT 124.150 154.575 124.290 154.730 ;
        RECT 126.360 154.670 126.680 154.730 ;
        RECT 127.755 154.685 128.045 154.915 ;
        RECT 130.960 154.870 131.280 154.930 ;
        RECT 132.430 154.915 132.570 155.410 ;
        RECT 134.680 155.210 134.970 155.255 ;
        RECT 136.780 155.210 137.070 155.255 ;
        RECT 138.350 155.210 138.640 155.255 ;
        RECT 134.680 155.070 138.640 155.210 ;
        RECT 138.870 155.210 139.010 155.410 ;
        RECT 142.920 155.410 145.525 155.550 ;
        RECT 142.920 155.350 143.240 155.410 ;
        RECT 145.235 155.365 145.525 155.410 ;
        RECT 143.380 155.210 143.700 155.270 ;
        RECT 138.870 155.070 143.700 155.210 ;
        RECT 134.680 155.025 134.970 155.070 ;
        RECT 136.780 155.025 137.070 155.070 ;
        RECT 138.350 155.025 138.640 155.070 ;
        RECT 143.380 155.010 143.700 155.070 ;
        RECT 132.355 154.870 132.645 154.915 ;
        RECT 130.960 154.730 132.645 154.870 ;
        RECT 130.960 154.670 131.280 154.730 ;
        RECT 132.355 154.685 132.645 154.730 ;
        RECT 133.720 154.870 134.040 154.930 ;
        RECT 134.195 154.870 134.485 154.915 ;
        RECT 133.720 154.730 134.485 154.870 ;
        RECT 133.720 154.670 134.040 154.730 ;
        RECT 134.195 154.685 134.485 154.730 ;
        RECT 135.075 154.870 135.365 154.915 ;
        RECT 136.265 154.870 136.555 154.915 ;
        RECT 138.785 154.870 139.075 154.915 ;
        RECT 135.075 154.730 139.075 154.870 ;
        RECT 135.075 154.685 135.365 154.730 ;
        RECT 136.265 154.685 136.555 154.730 ;
        RECT 138.785 154.685 139.075 154.730 ;
        RECT 119.475 154.530 119.765 154.575 ;
        RECT 117.635 154.390 119.765 154.530 ;
        RECT 117.635 154.345 117.925 154.390 ;
        RECT 119.000 154.330 119.320 154.390 ;
        RECT 119.475 154.345 119.765 154.390 ;
        RECT 124.075 154.345 124.365 154.575 ;
        RECT 124.535 154.345 124.825 154.575 ;
        RECT 135.530 154.530 135.820 154.575 ;
        RECT 141.540 154.530 141.860 154.590 ;
        RECT 135.530 154.390 141.860 154.530 ;
        RECT 135.530 154.345 135.820 154.390 ;
        RECT 63.815 154.190 64.105 154.235 ;
        RECT 57.910 154.050 64.105 154.190 ;
        RECT 36.200 153.990 36.520 154.050 ;
        RECT 36.720 154.005 37.010 154.050 ;
        RECT 63.815 154.005 64.105 154.050 ;
        RECT 35.740 153.850 36.060 153.910 ;
        RECT 38.515 153.850 38.805 153.895 ;
        RECT 35.740 153.710 38.805 153.850 ;
        RECT 35.740 153.650 36.060 153.710 ;
        RECT 38.515 153.665 38.805 153.710 ;
        RECT 42.180 153.850 42.500 153.910 ;
        RECT 45.860 153.850 46.180 153.910 ;
        RECT 42.180 153.710 46.180 153.850 ;
        RECT 42.180 153.650 42.500 153.710 ;
        RECT 45.860 153.650 46.180 153.710 ;
        RECT 57.360 153.850 57.680 153.910 ;
        RECT 61.515 153.850 61.805 153.895 ;
        RECT 57.360 153.710 61.805 153.850 ;
        RECT 57.360 153.650 57.680 153.710 ;
        RECT 61.515 153.665 61.805 153.710 ;
        RECT 62.420 153.650 62.740 153.910 ;
        RECT 63.890 153.850 64.030 154.005 ;
        RECT 64.720 153.990 65.040 154.250 ;
        RECT 77.615 154.190 77.905 154.235 ;
        RECT 79.990 154.190 80.130 154.330 ;
        RECT 77.615 154.050 80.130 154.190 ;
        RECT 92.950 154.190 93.240 154.235 ;
        RECT 93.700 154.190 94.020 154.250 ;
        RECT 92.950 154.050 94.020 154.190 ;
        RECT 77.615 154.005 77.905 154.050 ;
        RECT 92.950 154.005 93.240 154.050 ;
        RECT 93.700 153.990 94.020 154.050 ;
        RECT 94.620 154.190 94.940 154.250 ;
        RECT 95.860 154.190 96.150 154.235 ;
        RECT 113.650 154.190 113.940 154.235 ;
        RECT 115.410 154.190 115.550 154.330 ;
        RECT 94.620 154.050 96.150 154.190 ;
        RECT 94.620 153.990 94.940 154.050 ;
        RECT 95.860 154.005 96.150 154.050 ;
        RECT 96.550 154.050 102.210 154.190 ;
        RECT 68.400 153.850 68.720 153.910 ;
        RECT 63.890 153.710 68.720 153.850 ;
        RECT 68.400 153.650 68.720 153.710 ;
        RECT 74.840 153.850 75.160 153.910 ;
        RECT 76.220 153.850 76.540 153.910 ;
        RECT 76.695 153.850 76.985 153.895 ;
        RECT 74.840 153.710 76.985 153.850 ;
        RECT 74.840 153.650 75.160 153.710 ;
        RECT 76.220 153.650 76.540 153.710 ;
        RECT 76.695 153.665 76.985 153.710 ;
        RECT 79.440 153.650 79.760 153.910 ;
        RECT 83.580 153.850 83.900 153.910 ;
        RECT 96.550 153.850 96.690 154.050 ;
        RECT 83.580 153.710 96.690 153.850 ;
        RECT 98.300 153.850 98.620 153.910 ;
        RECT 101.535 153.850 101.825 153.895 ;
        RECT 98.300 153.710 101.825 153.850 ;
        RECT 102.070 153.850 102.210 154.050 ;
        RECT 113.650 154.050 115.550 154.190 ;
        RECT 118.080 154.190 118.400 154.250 ;
        RECT 124.610 154.190 124.750 154.345 ;
        RECT 141.540 154.330 141.860 154.390 ;
        RECT 142.015 154.345 142.305 154.575 ;
        RECT 118.080 154.050 124.750 154.190 ;
        RECT 137.400 154.190 137.720 154.250 ;
        RECT 142.090 154.190 142.230 154.345 ;
        RECT 137.400 154.050 142.230 154.190 ;
        RECT 113.650 154.005 113.940 154.050 ;
        RECT 118.080 153.990 118.400 154.050 ;
        RECT 137.400 153.990 137.720 154.050 ;
        RECT 115.780 153.850 116.100 153.910 ;
        RECT 102.070 153.710 116.100 153.850 ;
        RECT 83.580 153.650 83.900 153.710 ;
        RECT 98.300 153.650 98.620 153.710 ;
        RECT 101.535 153.665 101.825 153.710 ;
        RECT 115.780 153.650 116.100 153.710 ;
        RECT 117.175 153.850 117.465 153.895 ;
        RECT 120.840 153.850 121.160 153.910 ;
        RECT 117.175 153.710 121.160 153.850 ;
        RECT 117.175 153.665 117.465 153.710 ;
        RECT 120.840 153.650 121.160 153.710 ;
        RECT 124.995 153.850 125.285 153.895 ;
        RECT 125.440 153.850 125.760 153.910 ;
        RECT 124.995 153.710 125.760 153.850 ;
        RECT 124.995 153.665 125.285 153.710 ;
        RECT 125.440 153.650 125.760 153.710 ;
        RECT 126.820 153.650 127.140 153.910 ;
        RECT 127.295 153.850 127.585 153.895 ;
        RECT 129.135 153.850 129.425 153.895 ;
        RECT 127.295 153.710 129.425 153.850 ;
        RECT 127.295 153.665 127.585 153.710 ;
        RECT 129.135 153.665 129.425 153.710 ;
        RECT 141.095 153.850 141.385 153.895 ;
        RECT 142.000 153.850 142.320 153.910 ;
        RECT 141.095 153.710 142.320 153.850 ;
        RECT 141.095 153.665 141.385 153.710 ;
        RECT 142.000 153.650 142.320 153.710 ;
        RECT 17.270 153.030 146.990 153.510 ;
        RECT 38.040 152.630 38.360 152.890 ;
        RECT 38.960 152.830 39.280 152.890 ;
        RECT 39.435 152.830 39.725 152.875 ;
        RECT 38.960 152.690 39.725 152.830 ;
        RECT 38.960 152.630 39.280 152.690 ;
        RECT 39.435 152.645 39.725 152.690 ;
        RECT 40.355 152.830 40.645 152.875 ;
        RECT 40.800 152.830 41.120 152.890 ;
        RECT 40.355 152.690 41.120 152.830 ;
        RECT 40.355 152.645 40.645 152.690 ;
        RECT 40.800 152.630 41.120 152.690 ;
        RECT 59.215 152.830 59.505 152.875 ;
        RECT 61.040 152.830 61.360 152.890 ;
        RECT 59.215 152.690 61.360 152.830 ;
        RECT 59.215 152.645 59.505 152.690 ;
        RECT 61.040 152.630 61.360 152.690 ;
        RECT 67.035 152.830 67.325 152.875 ;
        RECT 68.400 152.830 68.720 152.890 ;
        RECT 78.520 152.830 78.840 152.890 ;
        RECT 80.360 152.830 80.680 152.890 ;
        RECT 67.035 152.690 68.720 152.830 ;
        RECT 67.035 152.645 67.325 152.690 ;
        RECT 68.400 152.630 68.720 152.690 ;
        RECT 72.170 152.690 80.680 152.830 ;
        RECT 36.215 152.490 36.505 152.535 ;
        RECT 39.880 152.490 40.200 152.550 ;
        RECT 32.150 152.350 36.505 152.490 ;
        RECT 29.300 151.810 29.620 151.870 ;
        RECT 32.150 151.855 32.290 152.350 ;
        RECT 36.215 152.305 36.505 152.350 ;
        RECT 37.210 152.350 40.200 152.490 ;
        RECT 37.210 152.195 37.350 152.350 ;
        RECT 39.880 152.290 40.200 152.350 ;
        RECT 54.140 152.490 54.460 152.550 ;
        RECT 58.295 152.490 58.585 152.535 ;
        RECT 58.740 152.490 59.060 152.550 ;
        RECT 60.580 152.490 60.900 152.550 ;
        RECT 54.140 152.350 59.060 152.490 ;
        RECT 54.140 152.290 54.460 152.350 ;
        RECT 58.295 152.305 58.585 152.350 ;
        RECT 58.740 152.290 59.060 152.350 ;
        RECT 59.750 152.350 60.900 152.490 ;
        RECT 35.755 151.965 36.045 152.195 ;
        RECT 37.135 151.965 37.425 152.195 ;
        RECT 38.500 152.150 38.820 152.210 ;
        RECT 41.275 152.150 41.565 152.195 ;
        RECT 38.500 152.010 41.565 152.150 ;
        RECT 32.075 151.810 32.365 151.855 ;
        RECT 35.280 151.810 35.600 151.870 ;
        RECT 29.300 151.670 32.365 151.810 ;
        RECT 29.300 151.610 29.620 151.670 ;
        RECT 32.075 151.625 32.365 151.670 ;
        RECT 33.990 151.670 35.600 151.810 ;
        RECT 35.830 151.810 35.970 151.965 ;
        RECT 38.500 151.950 38.820 152.010 ;
        RECT 41.275 151.965 41.565 152.010 ;
        RECT 53.680 152.150 54.000 152.210 ;
        RECT 54.600 152.150 54.920 152.210 ;
        RECT 53.680 152.010 54.920 152.150 ;
        RECT 53.680 151.950 54.000 152.010 ;
        RECT 54.600 151.950 54.920 152.010 ;
        RECT 55.520 151.950 55.840 152.210 ;
        RECT 56.455 152.150 56.745 152.195 ;
        RECT 59.750 152.150 59.890 152.350 ;
        RECT 60.580 152.290 60.900 152.350 ;
        RECT 61.470 152.490 61.760 152.535 ;
        RECT 62.420 152.490 62.740 152.550 ;
        RECT 61.470 152.350 62.740 152.490 ;
        RECT 61.470 152.305 61.760 152.350 ;
        RECT 62.420 152.290 62.740 152.350 ;
        RECT 56.455 152.010 59.890 152.150 ;
        RECT 56.455 151.965 56.745 152.010 ;
        RECT 60.120 151.950 60.440 152.210 ;
        RECT 72.170 152.195 72.310 152.690 ;
        RECT 78.520 152.630 78.840 152.690 ;
        RECT 80.360 152.630 80.680 152.690 ;
        RECT 93.700 152.830 94.020 152.890 ;
        RECT 93.700 152.690 104.050 152.830 ;
        RECT 93.700 152.630 94.020 152.690 ;
        RECT 103.910 152.550 104.050 152.690 ;
        RECT 119.000 152.630 119.320 152.890 ;
        RECT 123.615 152.830 123.905 152.875 ;
        RECT 127.280 152.830 127.600 152.890 ;
        RECT 123.615 152.690 127.600 152.830 ;
        RECT 123.615 152.645 123.905 152.690 ;
        RECT 127.280 152.630 127.600 152.690 ;
        RECT 130.960 152.630 131.280 152.890 ;
        RECT 138.780 152.630 139.100 152.890 ;
        RECT 141.095 152.830 141.385 152.875 ;
        RECT 142.920 152.830 143.240 152.890 ;
        RECT 141.095 152.690 143.240 152.830 ;
        RECT 141.095 152.645 141.385 152.690 ;
        RECT 142.920 152.630 143.240 152.690 ;
        RECT 143.840 152.830 144.160 152.890 ;
        RECT 145.235 152.830 145.525 152.875 ;
        RECT 143.840 152.690 145.525 152.830 ;
        RECT 143.840 152.630 144.160 152.690 ;
        RECT 145.235 152.645 145.525 152.690 ;
        RECT 86.340 152.490 86.660 152.550 ;
        RECT 90.480 152.490 90.800 152.550 ;
        RECT 94.160 152.490 94.480 152.550 ;
        RECT 74.470 152.350 86.660 152.490 ;
        RECT 72.095 151.965 72.385 152.195 ;
        RECT 73.015 152.150 73.305 152.195 ;
        RECT 73.920 152.150 74.240 152.210 ;
        RECT 74.470 152.195 74.610 152.350 ;
        RECT 86.340 152.290 86.660 152.350 ;
        RECT 88.730 152.350 94.480 152.490 ;
        RECT 73.015 152.010 74.240 152.150 ;
        RECT 73.015 151.965 73.305 152.010 ;
        RECT 73.920 151.950 74.240 152.010 ;
        RECT 74.395 151.965 74.685 152.195 ;
        RECT 85.880 152.150 86.200 152.210 ;
        RECT 88.730 152.195 88.870 152.350 ;
        RECT 90.480 152.290 90.800 152.350 ;
        RECT 94.160 152.290 94.480 152.350 ;
        RECT 103.820 152.490 104.140 152.550 ;
        RECT 112.100 152.490 112.420 152.550 ;
        RECT 133.720 152.490 134.040 152.550 ;
        RECT 103.820 152.350 105.890 152.490 ;
        RECT 103.820 152.290 104.140 152.350 ;
        RECT 87.320 152.150 87.610 152.195 ;
        RECT 85.880 152.010 87.610 152.150 ;
        RECT 85.880 151.950 86.200 152.010 ;
        RECT 87.320 151.965 87.610 152.010 ;
        RECT 88.655 151.965 88.945 152.195 ;
        RECT 92.795 152.150 93.085 152.195 ;
        RECT 96.920 152.150 97.240 152.210 ;
        RECT 92.795 152.010 97.240 152.150 ;
        RECT 92.795 151.965 93.085 152.010 ;
        RECT 96.920 151.950 97.240 152.010 ;
        RECT 98.300 151.950 98.620 152.210 ;
        RECT 100.615 152.150 100.905 152.195 ;
        RECT 101.060 152.150 101.380 152.210 ;
        RECT 100.615 152.010 101.380 152.150 ;
        RECT 100.615 151.965 100.905 152.010 ;
        RECT 101.060 151.950 101.380 152.010 ;
        RECT 104.740 151.950 105.060 152.210 ;
        RECT 105.750 152.195 105.890 152.350 ;
        RECT 112.100 152.350 134.040 152.490 ;
        RECT 112.100 152.290 112.420 152.350 ;
        RECT 105.675 151.965 105.965 152.195 ;
        RECT 113.450 152.150 113.740 152.195 ;
        RECT 117.160 152.150 117.480 152.210 ;
        RECT 113.450 152.010 117.480 152.150 ;
        RECT 113.450 151.965 113.740 152.010 ;
        RECT 117.160 151.950 117.480 152.010 ;
        RECT 120.855 152.150 121.145 152.195 ;
        RECT 121.300 152.150 121.620 152.210 ;
        RECT 120.855 152.010 121.620 152.150 ;
        RECT 120.855 151.965 121.145 152.010 ;
        RECT 121.300 151.950 121.620 152.010 ;
        RECT 121.775 151.965 122.065 152.195 ;
        RECT 38.960 151.810 39.280 151.870 ;
        RECT 35.830 151.670 39.280 151.810 ;
        RECT 33.990 151.515 34.130 151.670 ;
        RECT 35.280 151.610 35.600 151.670 ;
        RECT 38.960 151.610 39.280 151.670 ;
        RECT 61.015 151.810 61.305 151.855 ;
        RECT 62.205 151.810 62.495 151.855 ;
        RECT 64.725 151.810 65.015 151.855 ;
        RECT 61.015 151.670 65.015 151.810 ;
        RECT 61.015 151.625 61.305 151.670 ;
        RECT 62.205 151.625 62.495 151.670 ;
        RECT 64.725 151.625 65.015 151.670 ;
        RECT 72.555 151.810 72.845 151.855 ;
        RECT 75.300 151.810 75.620 151.870 ;
        RECT 72.555 151.670 75.620 151.810 ;
        RECT 72.555 151.625 72.845 151.670 ;
        RECT 75.300 151.610 75.620 151.670 ;
        RECT 75.775 151.625 76.065 151.855 ;
        RECT 78.060 151.810 78.380 151.870 ;
        RECT 78.995 151.810 79.285 151.855 ;
        RECT 78.060 151.670 79.285 151.810 ;
        RECT 33.915 151.285 34.205 151.515 ;
        RECT 60.620 151.470 60.910 151.515 ;
        RECT 62.720 151.470 63.010 151.515 ;
        RECT 64.290 151.470 64.580 151.515 ;
        RECT 60.620 151.330 64.580 151.470 ;
        RECT 75.850 151.470 75.990 151.625 ;
        RECT 78.060 151.610 78.380 151.670 ;
        RECT 78.995 151.625 79.285 151.670 ;
        RECT 79.440 151.610 79.760 151.870 ;
        RECT 84.065 151.810 84.355 151.855 ;
        RECT 86.585 151.810 86.875 151.855 ;
        RECT 87.775 151.810 88.065 151.855 ;
        RECT 84.065 151.670 88.065 151.810 ;
        RECT 84.065 151.625 84.355 151.670 ;
        RECT 86.585 151.625 86.875 151.670 ;
        RECT 87.775 151.625 88.065 151.670 ;
        RECT 93.700 151.610 94.020 151.870 ;
        RECT 94.175 151.810 94.465 151.855 ;
        RECT 95.095 151.810 95.385 151.855 ;
        RECT 94.175 151.670 95.385 151.810 ;
        RECT 94.175 151.625 94.465 151.670 ;
        RECT 95.095 151.625 95.385 151.670 ;
        RECT 103.375 151.810 103.665 151.855 ;
        RECT 106.135 151.810 106.425 151.855 ;
        RECT 103.375 151.670 106.425 151.810 ;
        RECT 103.375 151.625 103.665 151.670 ;
        RECT 106.135 151.625 106.425 151.670 ;
        RECT 109.340 151.810 109.660 151.870 ;
        RECT 112.100 151.810 112.420 151.870 ;
        RECT 109.340 151.670 112.420 151.810 ;
        RECT 109.340 151.610 109.660 151.670 ;
        RECT 112.100 151.610 112.420 151.670 ;
        RECT 112.995 151.810 113.285 151.855 ;
        RECT 114.185 151.810 114.475 151.855 ;
        RECT 116.705 151.810 116.995 151.855 ;
        RECT 112.995 151.670 116.995 151.810 ;
        RECT 112.995 151.625 113.285 151.670 ;
        RECT 114.185 151.625 114.475 151.670 ;
        RECT 116.705 151.625 116.995 151.670 ;
        RECT 120.380 151.810 120.700 151.870 ;
        RECT 121.850 151.810 121.990 151.965 ;
        RECT 122.220 151.950 122.540 152.210 ;
        RECT 122.695 152.150 122.985 152.195 ;
        RECT 123.600 152.150 123.920 152.210 ;
        RECT 124.150 152.195 124.290 152.350 ;
        RECT 133.720 152.290 134.040 152.350 ;
        RECT 139.790 152.350 142.230 152.490 ;
        RECT 125.440 152.195 125.760 152.210 ;
        RECT 122.695 152.010 123.920 152.150 ;
        RECT 122.695 151.965 122.985 152.010 ;
        RECT 123.600 151.950 123.920 152.010 ;
        RECT 124.075 151.965 124.365 152.195 ;
        RECT 125.410 152.150 125.760 152.195 ;
        RECT 125.245 152.010 125.760 152.150 ;
        RECT 125.410 151.965 125.760 152.010 ;
        RECT 125.440 151.950 125.760 151.965 ;
        RECT 137.400 151.950 137.720 152.210 ;
        RECT 139.790 152.195 139.930 152.350 ;
        RECT 142.090 152.210 142.230 152.350 ;
        RECT 139.715 151.965 140.005 152.195 ;
        RECT 140.160 151.950 140.480 152.210 ;
        RECT 142.000 151.950 142.320 152.210 ;
        RECT 120.380 151.670 121.990 151.810 ;
        RECT 124.955 151.810 125.245 151.855 ;
        RECT 126.145 151.810 126.435 151.855 ;
        RECT 128.665 151.810 128.955 151.855 ;
        RECT 143.840 151.810 144.160 151.870 ;
        RECT 124.955 151.670 128.955 151.810 ;
        RECT 120.380 151.610 120.700 151.670 ;
        RECT 124.955 151.625 125.245 151.670 ;
        RECT 126.145 151.625 126.435 151.670 ;
        RECT 128.665 151.625 128.955 151.670 ;
        RECT 138.410 151.670 144.160 151.810 ;
        RECT 79.530 151.470 79.670 151.610 ;
        RECT 75.850 151.330 79.670 151.470 ;
        RECT 84.500 151.470 84.790 151.515 ;
        RECT 86.070 151.470 86.360 151.515 ;
        RECT 88.170 151.470 88.460 151.515 ;
        RECT 84.500 151.330 88.460 151.470 ;
        RECT 60.620 151.285 60.910 151.330 ;
        RECT 62.720 151.285 63.010 151.330 ;
        RECT 64.290 151.285 64.580 151.330 ;
        RECT 84.500 151.285 84.790 151.330 ;
        RECT 86.070 151.285 86.360 151.330 ;
        RECT 88.170 151.285 88.460 151.330 ;
        RECT 91.875 151.470 92.165 151.515 ;
        RECT 94.620 151.470 94.940 151.530 ;
        RECT 138.410 151.515 138.550 151.670 ;
        RECT 143.840 151.610 144.160 151.670 ;
        RECT 91.875 151.330 94.940 151.470 ;
        RECT 91.875 151.285 92.165 151.330 ;
        RECT 32.060 151.130 32.380 151.190 ;
        RECT 33.990 151.130 34.130 151.285 ;
        RECT 94.620 151.270 94.940 151.330 ;
        RECT 112.600 151.470 112.890 151.515 ;
        RECT 114.700 151.470 114.990 151.515 ;
        RECT 116.270 151.470 116.560 151.515 ;
        RECT 112.600 151.330 116.560 151.470 ;
        RECT 112.600 151.285 112.890 151.330 ;
        RECT 114.700 151.285 114.990 151.330 ;
        RECT 116.270 151.285 116.560 151.330 ;
        RECT 124.560 151.470 124.850 151.515 ;
        RECT 126.660 151.470 126.950 151.515 ;
        RECT 128.230 151.470 128.520 151.515 ;
        RECT 124.560 151.330 128.520 151.470 ;
        RECT 124.560 151.285 124.850 151.330 ;
        RECT 126.660 151.285 126.950 151.330 ;
        RECT 128.230 151.285 128.520 151.330 ;
        RECT 138.335 151.285 138.625 151.515 ;
        RECT 32.060 150.990 34.130 151.130 ;
        RECT 34.375 151.130 34.665 151.175 ;
        RECT 35.280 151.130 35.600 151.190 ;
        RECT 34.375 150.990 35.600 151.130 ;
        RECT 32.060 150.930 32.380 150.990 ;
        RECT 34.375 150.945 34.665 150.990 ;
        RECT 35.280 150.930 35.600 150.990 ;
        RECT 38.500 150.930 38.820 151.190 ;
        RECT 54.600 151.130 54.920 151.190 ;
        RECT 55.075 151.130 55.365 151.175 ;
        RECT 54.600 150.990 55.365 151.130 ;
        RECT 54.600 150.930 54.920 150.990 ;
        RECT 55.075 150.945 55.365 150.990 ;
        RECT 58.280 150.930 58.600 151.190 ;
        RECT 73.460 150.930 73.780 151.190 ;
        RECT 76.680 150.930 77.000 151.190 ;
        RECT 81.755 151.130 82.045 151.175 ;
        RECT 83.580 151.130 83.900 151.190 ;
        RECT 81.755 150.990 83.900 151.130 ;
        RECT 81.755 150.945 82.045 150.990 ;
        RECT 83.580 150.930 83.900 150.990 ;
        RECT 94.160 151.130 94.480 151.190 ;
        RECT 103.835 151.130 104.125 151.175 ;
        RECT 94.160 150.990 104.125 151.130 ;
        RECT 94.160 150.930 94.480 150.990 ;
        RECT 103.835 150.945 104.125 150.990 ;
        RECT 17.270 150.310 146.990 150.790 ;
        RECT 34.375 150.110 34.665 150.155 ;
        RECT 35.740 150.110 36.060 150.170 ;
        RECT 34.375 149.970 36.060 150.110 ;
        RECT 34.375 149.925 34.665 149.970 ;
        RECT 35.740 149.910 36.060 149.970 ;
        RECT 40.800 150.110 41.120 150.170 ;
        RECT 42.655 150.110 42.945 150.155 ;
        RECT 40.800 149.970 42.945 150.110 ;
        RECT 40.800 149.910 41.120 149.970 ;
        RECT 42.655 149.925 42.945 149.970 ;
        RECT 52.775 150.110 53.065 150.155 ;
        RECT 58.280 150.110 58.600 150.170 ;
        RECT 52.775 149.970 58.600 150.110 ;
        RECT 52.775 149.925 53.065 149.970 ;
        RECT 58.280 149.910 58.600 149.970 ;
        RECT 64.720 150.110 65.040 150.170 ;
        RECT 67.035 150.110 67.325 150.155 ;
        RECT 64.720 149.970 67.325 150.110 ;
        RECT 64.720 149.910 65.040 149.970 ;
        RECT 67.035 149.925 67.325 149.970 ;
        RECT 67.955 149.925 68.245 150.155 ;
        RECT 76.680 150.110 77.000 150.170 ;
        RECT 70.790 149.970 77.000 150.110 ;
        RECT 36.240 149.770 36.530 149.815 ;
        RECT 38.340 149.770 38.630 149.815 ;
        RECT 39.910 149.770 40.200 149.815 ;
        RECT 36.240 149.630 40.200 149.770 ;
        RECT 36.240 149.585 36.530 149.630 ;
        RECT 38.340 149.585 38.630 149.630 ;
        RECT 39.910 149.585 40.200 149.630 ;
        RECT 53.680 149.770 54.000 149.830 ;
        RECT 56.440 149.770 56.760 149.830 ;
        RECT 66.100 149.770 66.420 149.830 ;
        RECT 68.030 149.770 68.170 149.925 ;
        RECT 53.680 149.630 54.830 149.770 ;
        RECT 53.680 149.570 54.000 149.630 ;
        RECT 34.820 149.430 35.140 149.490 ;
        RECT 35.740 149.430 36.060 149.490 ;
        RECT 34.820 149.290 36.060 149.430 ;
        RECT 34.820 149.230 35.140 149.290 ;
        RECT 35.740 149.230 36.060 149.290 ;
        RECT 36.635 149.430 36.925 149.475 ;
        RECT 37.825 149.430 38.115 149.475 ;
        RECT 40.345 149.430 40.635 149.475 ;
        RECT 36.635 149.290 40.635 149.430 ;
        RECT 36.635 149.245 36.925 149.290 ;
        RECT 37.825 149.245 38.115 149.290 ;
        RECT 40.345 149.245 40.635 149.290 ;
        RECT 52.760 149.430 53.080 149.490 ;
        RECT 54.690 149.475 54.830 149.630 ;
        RECT 55.150 149.630 64.030 149.770 ;
        RECT 55.150 149.490 55.290 149.630 ;
        RECT 56.440 149.570 56.760 149.630 ;
        RECT 54.155 149.430 54.445 149.475 ;
        RECT 52.760 149.290 54.445 149.430 ;
        RECT 52.760 149.230 53.080 149.290 ;
        RECT 54.155 149.245 54.445 149.290 ;
        RECT 54.615 149.245 54.905 149.475 ;
        RECT 32.535 149.090 32.825 149.135 ;
        RECT 38.500 149.090 38.820 149.150 ;
        RECT 32.535 148.950 38.820 149.090 ;
        RECT 32.535 148.905 32.825 148.950 ;
        RECT 38.500 148.890 38.820 148.950 ;
        RECT 50.000 149.090 50.320 149.150 ;
        RECT 53.695 149.090 53.985 149.135 ;
        RECT 50.000 148.950 53.985 149.090 ;
        RECT 54.690 149.090 54.830 149.245 ;
        RECT 55.060 149.230 55.380 149.490 ;
        RECT 60.120 149.430 60.440 149.490 ;
        RECT 61.515 149.430 61.805 149.475 ;
        RECT 62.420 149.430 62.740 149.490 ;
        RECT 60.120 149.290 63.570 149.430 ;
        RECT 60.120 149.230 60.440 149.290 ;
        RECT 61.515 149.245 61.805 149.290 ;
        RECT 62.420 149.230 62.740 149.290 ;
        RECT 62.880 149.090 63.200 149.150 ;
        RECT 63.430 149.135 63.570 149.290 ;
        RECT 54.690 148.950 63.200 149.090 ;
        RECT 50.000 148.890 50.320 148.950 ;
        RECT 53.695 148.905 53.985 148.950 ;
        RECT 62.880 148.890 63.200 148.950 ;
        RECT 63.355 148.905 63.645 149.135 ;
        RECT 63.890 149.090 64.030 149.630 ;
        RECT 66.100 149.630 68.170 149.770 ;
        RECT 66.100 149.570 66.420 149.630 ;
        RECT 68.860 149.430 69.180 149.490 ;
        RECT 70.790 149.475 70.930 149.970 ;
        RECT 76.680 149.910 77.000 149.970 ;
        RECT 85.880 149.910 86.200 150.170 ;
        RECT 86.340 150.110 86.660 150.170 ;
        RECT 88.655 150.110 88.945 150.155 ;
        RECT 86.340 149.970 88.945 150.110 ;
        RECT 86.340 149.910 86.660 149.970 ;
        RECT 88.655 149.925 88.945 149.970 ;
        RECT 97.395 150.110 97.685 150.155 ;
        RECT 101.060 150.110 101.380 150.170 ;
        RECT 97.395 149.970 101.380 150.110 ;
        RECT 97.395 149.925 97.685 149.970 ;
        RECT 101.060 149.910 101.380 149.970 ;
        RECT 123.155 150.110 123.445 150.155 ;
        RECT 126.820 150.110 127.140 150.170 ;
        RECT 123.155 149.970 127.140 150.110 ;
        RECT 123.155 149.925 123.445 149.970 ;
        RECT 126.820 149.910 127.140 149.970 ;
        RECT 134.180 150.110 134.500 150.170 ;
        RECT 142.475 150.110 142.765 150.155 ;
        RECT 134.180 149.970 142.765 150.110 ;
        RECT 134.180 149.910 134.500 149.970 ;
        RECT 142.475 149.925 142.765 149.970 ;
        RECT 144.760 149.910 145.080 150.170 ;
        RECT 71.660 149.770 71.950 149.815 ;
        RECT 73.760 149.770 74.050 149.815 ;
        RECT 75.330 149.770 75.620 149.815 ;
        RECT 71.660 149.630 75.620 149.770 ;
        RECT 71.660 149.585 71.950 149.630 ;
        RECT 73.760 149.585 74.050 149.630 ;
        RECT 75.330 149.585 75.620 149.630 ;
        RECT 78.060 149.770 78.380 149.830 ;
        RECT 90.980 149.770 91.270 149.815 ;
        RECT 93.080 149.770 93.370 149.815 ;
        RECT 94.650 149.770 94.940 149.815 ;
        RECT 78.060 149.630 82.890 149.770 ;
        RECT 78.060 149.570 78.380 149.630 ;
        RECT 68.860 149.290 69.550 149.430 ;
        RECT 68.860 149.230 69.180 149.290 ;
        RECT 69.410 149.135 69.550 149.290 ;
        RECT 70.715 149.245 71.005 149.475 ;
        RECT 72.055 149.430 72.345 149.475 ;
        RECT 73.245 149.430 73.535 149.475 ;
        RECT 75.765 149.430 76.055 149.475 ;
        RECT 72.055 149.290 76.055 149.430 ;
        RECT 72.055 149.245 72.345 149.290 ;
        RECT 73.245 149.245 73.535 149.290 ;
        RECT 75.765 149.245 76.055 149.290 ;
        RECT 77.140 149.430 77.460 149.490 ;
        RECT 82.750 149.475 82.890 149.630 ;
        RECT 90.980 149.630 94.940 149.770 ;
        RECT 90.980 149.585 91.270 149.630 ;
        RECT 93.080 149.585 93.370 149.630 ;
        RECT 94.650 149.585 94.940 149.630 ;
        RECT 102.440 149.570 102.760 149.830 ;
        RECT 106.120 149.570 106.440 149.830 ;
        RECT 118.540 149.770 118.860 149.830 ;
        RECT 124.075 149.770 124.365 149.815 ;
        RECT 129.580 149.770 129.900 149.830 ;
        RECT 118.540 149.630 123.370 149.770 ;
        RECT 118.540 149.570 118.860 149.630 ;
        RECT 81.295 149.430 81.585 149.475 ;
        RECT 77.140 149.290 81.585 149.430 ;
        RECT 77.140 149.230 77.460 149.290 ;
        RECT 81.295 149.245 81.585 149.290 ;
        RECT 82.675 149.245 82.965 149.475 ;
        RECT 83.580 149.230 83.900 149.490 ;
        RECT 90.480 149.230 90.800 149.490 ;
        RECT 91.375 149.430 91.665 149.475 ;
        RECT 92.565 149.430 92.855 149.475 ;
        RECT 95.085 149.430 95.375 149.475 ;
        RECT 122.680 149.430 123.000 149.490 ;
        RECT 91.375 149.290 95.375 149.430 ;
        RECT 91.375 149.245 91.665 149.290 ;
        RECT 92.565 149.245 92.855 149.290 ;
        RECT 95.085 149.245 95.375 149.290 ;
        RECT 120.470 149.290 123.000 149.430 ;
        RECT 123.230 149.430 123.370 149.630 ;
        RECT 124.075 149.630 129.900 149.770 ;
        RECT 124.075 149.585 124.365 149.630 ;
        RECT 129.580 149.570 129.900 149.630 ;
        RECT 128.660 149.430 128.980 149.490 ;
        RECT 136.020 149.430 136.340 149.490 ;
        RECT 137.415 149.430 137.705 149.475 ;
        RECT 123.230 149.290 123.830 149.430 ;
        RECT 63.890 148.950 69.090 149.090 ;
        RECT 32.060 148.750 32.380 148.810 ;
        RECT 34.375 148.750 34.665 148.795 ;
        RECT 34.820 148.750 35.140 148.810 ;
        RECT 36.980 148.750 37.270 148.795 ;
        RECT 32.060 148.610 35.140 148.750 ;
        RECT 32.060 148.550 32.380 148.610 ;
        RECT 34.375 148.565 34.665 148.610 ;
        RECT 34.820 148.550 35.140 148.610 ;
        RECT 35.370 148.610 37.270 148.750 ;
        RECT 35.370 148.455 35.510 148.610 ;
        RECT 36.980 148.565 37.270 148.610 ;
        RECT 44.940 148.550 45.260 148.810 ;
        RECT 49.095 148.750 49.385 148.795 ;
        RECT 57.835 148.750 58.125 148.795 ;
        RECT 66.560 148.750 66.880 148.810 ;
        RECT 68.950 148.795 69.090 148.950 ;
        RECT 69.335 148.905 69.625 149.135 ;
        RECT 69.795 148.905 70.085 149.135 ;
        RECT 70.240 149.090 70.560 149.150 ;
        RECT 71.175 149.090 71.465 149.135 ;
        RECT 70.240 148.950 71.465 149.090 ;
        RECT 49.095 148.610 66.880 148.750 ;
        RECT 49.095 148.565 49.385 148.610 ;
        RECT 57.835 148.565 58.125 148.610 ;
        RECT 66.560 148.550 66.880 148.610 ;
        RECT 68.875 148.565 69.165 148.795 ;
        RECT 35.295 148.225 35.585 148.455 ;
        RECT 55.520 148.410 55.840 148.470 ;
        RECT 64.720 148.410 65.040 148.470 ;
        RECT 67.825 148.410 68.115 148.455 ;
        RECT 55.520 148.270 68.115 148.410 ;
        RECT 69.870 148.410 70.010 148.905 ;
        RECT 70.240 148.890 70.560 148.950 ;
        RECT 71.175 148.905 71.465 148.950 ;
        RECT 79.440 148.890 79.760 149.150 ;
        RECT 80.360 149.090 80.680 149.150 ;
        RECT 86.355 149.090 86.645 149.135 ;
        RECT 80.360 148.950 86.645 149.090 ;
        RECT 80.360 148.890 80.680 148.950 ;
        RECT 86.355 148.905 86.645 148.950 ;
        RECT 87.720 148.890 88.040 149.150 ;
        RECT 91.830 149.090 92.120 149.135 ;
        RECT 94.160 149.090 94.480 149.150 ;
        RECT 91.830 148.950 94.480 149.090 ;
        RECT 91.830 148.905 92.120 148.950 ;
        RECT 94.160 148.890 94.480 148.950 ;
        RECT 98.760 149.090 99.080 149.150 ;
        RECT 100.155 149.090 100.445 149.135 ;
        RECT 102.900 149.090 103.220 149.150 ;
        RECT 119.460 149.090 119.780 149.150 ;
        RECT 120.470 149.135 120.610 149.290 ;
        RECT 122.680 149.230 123.000 149.290 ;
        RECT 98.760 148.950 103.220 149.090 ;
        RECT 98.760 148.890 99.080 148.950 ;
        RECT 100.155 148.905 100.445 148.950 ;
        RECT 102.900 148.890 103.220 148.950 ;
        RECT 103.450 148.950 119.780 149.090 ;
        RECT 70.715 148.750 71.005 148.795 ;
        RECT 72.400 148.750 72.690 148.795 ;
        RECT 70.715 148.610 72.690 148.750 ;
        RECT 70.715 148.565 71.005 148.610 ;
        RECT 72.400 148.565 72.690 148.610 ;
        RECT 78.520 148.550 78.840 148.810 ;
        RECT 78.980 148.750 79.300 148.810 ;
        RECT 79.915 148.750 80.205 148.795 ;
        RECT 78.980 148.610 80.205 148.750 ;
        RECT 78.980 148.550 79.300 148.610 ;
        RECT 79.915 148.565 80.205 148.610 ;
        RECT 81.740 148.750 82.060 148.810 ;
        RECT 84.055 148.750 84.345 148.795 ;
        RECT 81.740 148.610 84.345 148.750 ;
        RECT 81.740 148.550 82.060 148.610 ;
        RECT 84.055 148.565 84.345 148.610 ;
        RECT 88.180 148.750 88.500 148.810 ;
        RECT 98.315 148.750 98.605 148.795 ;
        RECT 103.450 148.750 103.590 148.950 ;
        RECT 119.460 148.890 119.780 148.950 ;
        RECT 120.395 148.905 120.685 149.135 ;
        RECT 121.300 148.890 121.620 149.150 ;
        RECT 121.760 148.890 122.080 149.150 ;
        RECT 122.235 149.090 122.525 149.135 ;
        RECT 123.140 149.090 123.460 149.150 ;
        RECT 123.690 149.135 123.830 149.290 ;
        RECT 124.150 149.290 132.110 149.430 ;
        RECT 124.150 149.150 124.290 149.290 ;
        RECT 128.660 149.230 128.980 149.290 ;
        RECT 122.235 148.950 123.460 149.090 ;
        RECT 122.235 148.905 122.525 148.950 ;
        RECT 123.140 148.890 123.460 148.950 ;
        RECT 123.615 148.905 123.905 149.135 ;
        RECT 124.060 148.890 124.380 149.150 ;
        RECT 124.535 149.090 124.825 149.135 ;
        RECT 125.900 149.090 126.220 149.150 ;
        RECT 124.535 148.950 126.220 149.090 ;
        RECT 124.535 148.905 124.825 148.950 ;
        RECT 125.900 148.890 126.220 148.950 ;
        RECT 130.040 148.890 130.360 149.150 ;
        RECT 130.500 149.090 130.820 149.150 ;
        RECT 131.970 149.135 132.110 149.290 ;
        RECT 136.020 149.290 137.705 149.430 ;
        RECT 136.020 149.230 136.340 149.290 ;
        RECT 137.415 149.245 137.705 149.290 ;
        RECT 130.975 149.090 131.265 149.135 ;
        RECT 130.500 148.950 131.265 149.090 ;
        RECT 130.500 148.890 130.820 148.950 ;
        RECT 130.975 148.905 131.265 148.950 ;
        RECT 131.895 148.905 132.185 149.135 ;
        RECT 140.160 149.090 140.480 149.150 ;
        RECT 141.555 149.090 141.845 149.135 ;
        RECT 140.160 148.950 141.845 149.090 ;
        RECT 140.160 148.890 140.480 148.950 ;
        RECT 141.555 148.905 141.845 148.950 ;
        RECT 143.380 148.890 143.700 149.150 ;
        RECT 143.840 148.890 144.160 149.150 ;
        RECT 88.180 148.610 103.590 148.750 ;
        RECT 103.835 148.750 104.125 148.795 ;
        RECT 104.295 148.750 104.585 148.795 ;
        RECT 131.435 148.750 131.725 148.795 ;
        RECT 136.495 148.750 136.785 148.795 ;
        RECT 103.835 148.610 130.270 148.750 ;
        RECT 88.180 148.550 88.500 148.610 ;
        RECT 98.315 148.565 98.605 148.610 ;
        RECT 103.835 148.565 104.125 148.610 ;
        RECT 104.295 148.565 104.585 148.610 ;
        RECT 130.130 148.470 130.270 148.610 ;
        RECT 131.435 148.610 132.110 148.750 ;
        RECT 131.435 148.565 131.725 148.610 ;
        RECT 131.970 148.470 132.110 148.610 ;
        RECT 132.890 148.610 136.785 148.750 ;
        RECT 76.220 148.410 76.540 148.470 ;
        RECT 69.870 148.270 76.540 148.410 ;
        RECT 55.520 148.210 55.840 148.270 ;
        RECT 64.720 148.210 65.040 148.270 ;
        RECT 67.825 148.225 68.115 148.270 ;
        RECT 76.220 148.210 76.540 148.270 ;
        RECT 78.075 148.410 78.365 148.455 ;
        RECT 79.440 148.410 79.760 148.470 ;
        RECT 78.075 148.270 79.760 148.410 ;
        RECT 78.075 148.225 78.365 148.270 ;
        RECT 79.440 148.210 79.760 148.270 ;
        RECT 86.340 148.410 86.660 148.470 ;
        RECT 86.815 148.410 87.105 148.455 ;
        RECT 86.340 148.270 87.105 148.410 ;
        RECT 86.340 148.210 86.660 148.270 ;
        RECT 86.815 148.225 87.105 148.270 ;
        RECT 101.520 148.210 101.840 148.470 ;
        RECT 106.580 148.210 106.900 148.470 ;
        RECT 130.040 148.210 130.360 148.470 ;
        RECT 131.880 148.210 132.200 148.470 ;
        RECT 132.890 148.455 133.030 148.610 ;
        RECT 136.495 148.565 136.785 148.610 ;
        RECT 132.815 148.225 133.105 148.455 ;
        RECT 134.640 148.210 134.960 148.470 ;
        RECT 136.955 148.410 137.245 148.455 ;
        RECT 138.795 148.410 139.085 148.455 ;
        RECT 136.955 148.270 139.085 148.410 ;
        RECT 136.955 148.225 137.245 148.270 ;
        RECT 138.795 148.225 139.085 148.270 ;
        RECT 17.270 147.590 146.990 148.070 ;
        RECT 29.300 147.190 29.620 147.450 ;
        RECT 35.280 147.390 35.600 147.450 ;
        RECT 34.910 147.250 35.600 147.390 ;
        RECT 34.910 147.095 35.050 147.250 ;
        RECT 35.280 147.190 35.600 147.250 ;
        RECT 39.420 147.390 39.740 147.450 ;
        RECT 42.180 147.390 42.500 147.450 ;
        RECT 39.420 147.250 42.500 147.390 ;
        RECT 39.420 147.190 39.740 147.250 ;
        RECT 42.180 147.190 42.500 147.250 ;
        RECT 55.060 147.390 55.380 147.450 ;
        RECT 55.535 147.390 55.825 147.435 ;
        RECT 66.100 147.390 66.420 147.450 ;
        RECT 55.060 147.250 55.825 147.390 ;
        RECT 55.060 147.190 55.380 147.250 ;
        RECT 55.535 147.205 55.825 147.250 ;
        RECT 63.890 147.250 66.420 147.390 ;
        RECT 34.880 146.865 35.170 147.095 ;
        RECT 44.940 147.050 45.260 147.110 ;
        RECT 53.235 147.050 53.525 147.095 ;
        RECT 57.360 147.050 57.680 147.110 ;
        RECT 36.290 146.910 45.630 147.050 ;
        RECT 20.115 146.710 20.405 146.755 ;
        RECT 22.860 146.710 23.180 146.770 ;
        RECT 20.115 146.570 23.180 146.710 ;
        RECT 20.115 146.525 20.405 146.570 ;
        RECT 22.860 146.510 23.180 146.570 ;
        RECT 35.740 146.710 36.060 146.770 ;
        RECT 36.290 146.755 36.430 146.910 ;
        RECT 44.940 146.850 45.260 146.910 ;
        RECT 36.215 146.710 36.505 146.755 ;
        RECT 35.740 146.570 36.505 146.710 ;
        RECT 35.740 146.510 36.060 146.570 ;
        RECT 36.215 146.525 36.505 146.570 ;
        RECT 38.975 146.710 39.265 146.755 ;
        RECT 39.420 146.710 39.740 146.770 ;
        RECT 38.975 146.570 39.740 146.710 ;
        RECT 38.975 146.525 39.265 146.570 ;
        RECT 39.420 146.510 39.740 146.570 ;
        RECT 39.895 146.525 40.185 146.755 ;
        RECT 41.275 146.525 41.565 146.755 ;
        RECT 31.625 146.370 31.915 146.415 ;
        RECT 34.145 146.370 34.435 146.415 ;
        RECT 35.335 146.370 35.625 146.415 ;
        RECT 31.625 146.230 35.625 146.370 ;
        RECT 31.625 146.185 31.915 146.230 ;
        RECT 34.145 146.185 34.435 146.230 ;
        RECT 35.335 146.185 35.625 146.230 ;
        RECT 38.500 146.370 38.820 146.430 ;
        RECT 39.970 146.370 40.110 146.525 ;
        RECT 38.500 146.230 40.110 146.370 ;
        RECT 41.350 146.370 41.490 146.525 ;
        RECT 42.180 146.510 42.500 146.770 ;
        RECT 42.640 146.510 42.960 146.770 ;
        RECT 45.490 146.755 45.630 146.910 ;
        RECT 53.235 146.910 57.680 147.050 ;
        RECT 53.235 146.865 53.525 146.910 ;
        RECT 57.360 146.850 57.680 146.910 ;
        RECT 61.040 147.095 61.360 147.110 ;
        RECT 61.040 147.050 61.390 147.095 ;
        RECT 62.880 147.050 63.200 147.110 ;
        RECT 63.890 147.095 64.030 147.250 ;
        RECT 66.100 147.190 66.420 147.250 ;
        RECT 77.155 147.390 77.445 147.435 ;
        RECT 78.980 147.390 79.300 147.450 ;
        RECT 77.155 147.250 79.300 147.390 ;
        RECT 77.155 147.205 77.445 147.250 ;
        RECT 78.980 147.190 79.300 147.250 ;
        RECT 81.755 147.390 82.045 147.435 ;
        RECT 87.720 147.390 88.040 147.450 ;
        RECT 81.755 147.250 88.040 147.390 ;
        RECT 81.755 147.205 82.045 147.250 ;
        RECT 87.720 147.190 88.040 147.250 ;
        RECT 100.615 147.390 100.905 147.435 ;
        RECT 104.740 147.390 105.060 147.450 ;
        RECT 100.615 147.250 105.060 147.390 ;
        RECT 100.615 147.205 100.905 147.250 ;
        RECT 104.740 147.190 105.060 147.250 ;
        RECT 105.660 147.390 105.980 147.450 ;
        RECT 108.895 147.390 109.185 147.435 ;
        RECT 139.700 147.390 140.020 147.450 ;
        RECT 105.660 147.250 140.020 147.390 ;
        RECT 105.660 147.190 105.980 147.250 ;
        RECT 108.895 147.205 109.185 147.250 ;
        RECT 139.700 147.190 140.020 147.250 ;
        RECT 140.160 147.190 140.480 147.450 ;
        RECT 141.555 147.205 141.845 147.435 ;
        RECT 63.815 147.050 64.105 147.095 ;
        RECT 61.040 146.910 61.555 147.050 ;
        RECT 62.880 146.910 64.105 147.050 ;
        RECT 61.040 146.865 61.390 146.910 ;
        RECT 61.040 146.850 61.360 146.865 ;
        RECT 62.880 146.850 63.200 146.910 ;
        RECT 63.815 146.865 64.105 146.910 ;
        RECT 64.720 146.850 65.040 147.110 ;
        RECT 71.590 147.050 71.880 147.095 ;
        RECT 73.460 147.050 73.780 147.110 ;
        RECT 71.590 146.910 73.780 147.050 ;
        RECT 71.590 146.865 71.880 146.910 ;
        RECT 73.460 146.850 73.780 146.910 ;
        RECT 78.520 147.050 78.840 147.110 ;
        RECT 101.520 147.050 101.840 147.110 ;
        RECT 103.220 147.050 103.510 147.095 ;
        RECT 78.520 146.910 86.570 147.050 ;
        RECT 78.520 146.850 78.840 146.910 ;
        RECT 45.415 146.525 45.705 146.755 ;
        RECT 50.000 146.510 50.320 146.770 ;
        RECT 50.935 146.710 51.225 146.755 ;
        RECT 51.395 146.710 51.685 146.755 ;
        RECT 55.520 146.710 55.840 146.770 ;
        RECT 50.935 146.570 55.840 146.710 ;
        RECT 50.935 146.525 51.225 146.570 ;
        RECT 51.395 146.525 51.685 146.570 ;
        RECT 55.520 146.510 55.840 146.570 ;
        RECT 62.420 146.510 62.740 146.770 ;
        RECT 68.860 146.710 69.180 146.770 ;
        RECT 79.900 146.710 80.220 146.770 ;
        RECT 86.430 146.755 86.570 146.910 ;
        RECT 99.310 146.910 100.370 147.050 ;
        RECT 85.895 146.710 86.185 146.755 ;
        RECT 68.860 146.570 79.670 146.710 ;
        RECT 68.860 146.510 69.180 146.570 ;
        RECT 46.780 146.370 47.100 146.430 ;
        RECT 41.350 146.230 47.100 146.370 ;
        RECT 38.500 146.170 38.820 146.230 ;
        RECT 32.060 146.030 32.350 146.075 ;
        RECT 33.630 146.030 33.920 146.075 ;
        RECT 35.730 146.030 36.020 146.075 ;
        RECT 32.060 145.890 36.020 146.030 ;
        RECT 39.970 146.030 40.110 146.230 ;
        RECT 46.780 146.170 47.100 146.230 ;
        RECT 49.095 146.370 49.385 146.415 ;
        RECT 52.760 146.370 53.080 146.430 ;
        RECT 49.095 146.230 53.080 146.370 ;
        RECT 49.095 146.185 49.385 146.230 ;
        RECT 52.760 146.170 53.080 146.230 ;
        RECT 57.845 146.370 58.135 146.415 ;
        RECT 60.365 146.370 60.655 146.415 ;
        RECT 61.555 146.370 61.845 146.415 ;
        RECT 57.845 146.230 61.845 146.370 ;
        RECT 57.845 146.185 58.135 146.230 ;
        RECT 60.365 146.185 60.655 146.230 ;
        RECT 61.555 146.185 61.845 146.230 ;
        RECT 70.240 146.170 70.560 146.430 ;
        RECT 71.135 146.370 71.425 146.415 ;
        RECT 72.325 146.370 72.615 146.415 ;
        RECT 74.845 146.370 75.135 146.415 ;
        RECT 71.135 146.230 75.135 146.370 ;
        RECT 71.135 146.185 71.425 146.230 ;
        RECT 72.325 146.185 72.615 146.230 ;
        RECT 74.845 146.185 75.135 146.230 ;
        RECT 78.980 146.170 79.300 146.430 ;
        RECT 79.530 146.370 79.670 146.570 ;
        RECT 79.900 146.570 86.185 146.710 ;
        RECT 79.900 146.510 80.220 146.570 ;
        RECT 85.895 146.525 86.185 146.570 ;
        RECT 86.355 146.525 86.645 146.755 ;
        RECT 97.380 146.710 97.700 146.770 ;
        RECT 97.855 146.710 98.145 146.755 ;
        RECT 97.380 146.570 98.145 146.710 ;
        RECT 97.380 146.510 97.700 146.570 ;
        RECT 97.855 146.525 98.145 146.570 ;
        RECT 98.315 146.710 98.605 146.755 ;
        RECT 98.760 146.710 99.080 146.770 ;
        RECT 99.310 146.755 99.450 146.910 ;
        RECT 98.315 146.570 99.080 146.710 ;
        RECT 98.315 146.525 98.605 146.570 ;
        RECT 98.760 146.510 99.080 146.570 ;
        RECT 99.235 146.525 99.525 146.755 ;
        RECT 99.680 146.510 100.000 146.770 ;
        RECT 100.230 146.710 100.370 146.910 ;
        RECT 101.520 146.910 103.510 147.050 ;
        RECT 101.520 146.850 101.840 146.910 ;
        RECT 103.220 146.865 103.510 146.910 ;
        RECT 106.580 147.050 106.900 147.110 ;
        RECT 110.580 147.050 110.870 147.095 ;
        RECT 106.580 146.910 110.870 147.050 ;
        RECT 106.580 146.850 106.900 146.910 ;
        RECT 110.580 146.865 110.870 146.910 ;
        RECT 128.660 147.050 128.980 147.110 ;
        RECT 128.660 146.910 130.270 147.050 ;
        RECT 128.660 146.850 128.980 146.910 ;
        RECT 105.660 146.710 105.980 146.770 ;
        RECT 100.230 146.570 105.980 146.710 ;
        RECT 105.660 146.510 105.980 146.570 ;
        RECT 109.340 146.510 109.660 146.770 ;
        RECT 117.620 146.710 117.940 146.770 ;
        RECT 120.380 146.710 120.700 146.770 ;
        RECT 123.615 146.710 123.905 146.755 ;
        RECT 117.620 146.570 123.905 146.710 ;
        RECT 117.620 146.510 117.940 146.570 ;
        RECT 120.380 146.510 120.700 146.570 ;
        RECT 123.615 146.525 123.905 146.570 ;
        RECT 129.120 146.710 129.440 146.770 ;
        RECT 129.595 146.710 129.885 146.755 ;
        RECT 129.120 146.570 129.885 146.710 ;
        RECT 130.130 146.710 130.270 146.910 ;
        RECT 130.500 146.850 130.820 147.110 ;
        RECT 130.975 147.050 131.265 147.095 ;
        RECT 132.800 147.050 133.120 147.110 ;
        RECT 134.640 147.095 134.960 147.110 ;
        RECT 134.610 147.050 134.960 147.095 ;
        RECT 130.975 146.910 133.120 147.050 ;
        RECT 134.445 146.910 134.960 147.050 ;
        RECT 130.975 146.865 131.265 146.910 ;
        RECT 132.800 146.850 133.120 146.910 ;
        RECT 134.610 146.865 134.960 146.910 ;
        RECT 134.640 146.850 134.960 146.865 ;
        RECT 131.435 146.710 131.725 146.755 ;
        RECT 130.130 146.570 131.725 146.710 ;
        RECT 129.120 146.510 129.440 146.570 ;
        RECT 129.595 146.525 129.885 146.570 ;
        RECT 131.435 146.525 131.725 146.570 ;
        RECT 133.275 146.710 133.565 146.755 ;
        RECT 133.720 146.710 134.040 146.770 ;
        RECT 133.275 146.570 134.040 146.710 ;
        RECT 140.250 146.710 140.390 147.190 ;
        RECT 140.635 146.710 140.925 146.755 ;
        RECT 140.250 146.570 140.925 146.710 ;
        RECT 141.630 146.710 141.770 147.205 ;
        RECT 144.760 147.190 145.080 147.450 ;
        RECT 142.015 146.710 142.305 146.755 ;
        RECT 141.630 146.570 142.305 146.710 ;
        RECT 133.275 146.525 133.565 146.570 ;
        RECT 133.720 146.510 134.040 146.570 ;
        RECT 140.635 146.525 140.925 146.570 ;
        RECT 142.015 146.525 142.305 146.570 ;
        RECT 143.855 146.525 144.145 146.755 ;
        RECT 81.740 146.370 82.060 146.430 ;
        RECT 79.530 146.230 82.060 146.370 ;
        RECT 81.740 146.170 82.060 146.230 ;
        RECT 82.200 146.170 82.520 146.430 ;
        RECT 87.720 146.370 88.040 146.430 ;
        RECT 101.995 146.370 102.285 146.415 ;
        RECT 87.720 146.230 102.285 146.370 ;
        RECT 87.720 146.170 88.040 146.230 ;
        RECT 101.995 146.185 102.285 146.230 ;
        RECT 102.875 146.370 103.165 146.415 ;
        RECT 104.065 146.370 104.355 146.415 ;
        RECT 106.585 146.370 106.875 146.415 ;
        RECT 102.875 146.230 106.875 146.370 ;
        RECT 102.875 146.185 103.165 146.230 ;
        RECT 104.065 146.185 104.355 146.230 ;
        RECT 106.585 146.185 106.875 146.230 ;
        RECT 110.235 146.370 110.525 146.415 ;
        RECT 111.425 146.370 111.715 146.415 ;
        RECT 113.945 146.370 114.235 146.415 ;
        RECT 110.235 146.230 114.235 146.370 ;
        RECT 110.235 146.185 110.525 146.230 ;
        RECT 111.425 146.185 111.715 146.230 ;
        RECT 113.945 146.185 114.235 146.230 ;
        RECT 134.155 146.370 134.445 146.415 ;
        RECT 135.345 146.370 135.635 146.415 ;
        RECT 137.865 146.370 138.155 146.415 ;
        RECT 134.155 146.230 138.155 146.370 ;
        RECT 134.155 146.185 134.445 146.230 ;
        RECT 135.345 146.185 135.635 146.230 ;
        RECT 137.865 146.185 138.155 146.230 ;
        RECT 41.720 146.030 42.040 146.090 ;
        RECT 42.640 146.030 42.960 146.090 ;
        RECT 39.970 145.890 42.960 146.030 ;
        RECT 32.060 145.845 32.350 145.890 ;
        RECT 33.630 145.845 33.920 145.890 ;
        RECT 35.730 145.845 36.020 145.890 ;
        RECT 41.720 145.830 42.040 145.890 ;
        RECT 42.640 145.830 42.960 145.890 ;
        RECT 58.280 146.030 58.570 146.075 ;
        RECT 59.850 146.030 60.140 146.075 ;
        RECT 61.950 146.030 62.240 146.075 ;
        RECT 58.280 145.890 62.240 146.030 ;
        RECT 58.280 145.845 58.570 145.890 ;
        RECT 59.850 145.845 60.140 145.890 ;
        RECT 61.950 145.845 62.240 145.890 ;
        RECT 70.740 146.030 71.030 146.075 ;
        RECT 72.840 146.030 73.130 146.075 ;
        RECT 74.410 146.030 74.700 146.075 ;
        RECT 70.740 145.890 74.700 146.030 ;
        RECT 70.740 145.845 71.030 145.890 ;
        RECT 72.840 145.845 73.130 145.890 ;
        RECT 74.410 145.845 74.700 145.890 ;
        RECT 79.440 146.030 79.760 146.090 ;
        RECT 102.480 146.030 102.770 146.075 ;
        RECT 104.580 146.030 104.870 146.075 ;
        RECT 106.150 146.030 106.440 146.075 ;
        RECT 79.440 145.890 86.570 146.030 ;
        RECT 79.440 145.830 79.760 145.890 ;
        RECT 86.430 145.750 86.570 145.890 ;
        RECT 102.480 145.890 106.440 146.030 ;
        RECT 102.480 145.845 102.770 145.890 ;
        RECT 104.580 145.845 104.870 145.890 ;
        RECT 106.150 145.845 106.440 145.890 ;
        RECT 109.840 146.030 110.130 146.075 ;
        RECT 111.940 146.030 112.230 146.075 ;
        RECT 113.510 146.030 113.800 146.075 ;
        RECT 133.760 146.030 134.050 146.075 ;
        RECT 135.860 146.030 136.150 146.075 ;
        RECT 137.430 146.030 137.720 146.075 ;
        RECT 143.930 146.030 144.070 146.525 ;
        RECT 109.840 145.890 113.800 146.030 ;
        RECT 109.840 145.845 110.130 145.890 ;
        RECT 111.940 145.845 112.230 145.890 ;
        RECT 113.510 145.845 113.800 145.890 ;
        RECT 116.330 145.890 133.030 146.030 ;
        RECT 116.330 145.750 116.470 145.890 ;
        RECT 19.180 145.490 19.500 145.750 ;
        RECT 36.660 145.690 36.980 145.750 ;
        RECT 38.055 145.690 38.345 145.735 ;
        RECT 36.660 145.550 38.345 145.690 ;
        RECT 36.660 145.490 36.980 145.550 ;
        RECT 38.055 145.505 38.345 145.550 ;
        RECT 39.420 145.690 39.740 145.750 ;
        RECT 40.355 145.690 40.645 145.735 ;
        RECT 39.420 145.550 40.645 145.690 ;
        RECT 39.420 145.490 39.740 145.550 ;
        RECT 40.355 145.505 40.645 145.550 ;
        RECT 42.180 145.690 42.500 145.750 ;
        RECT 45.860 145.690 46.180 145.750 ;
        RECT 49.080 145.690 49.400 145.750 ;
        RECT 42.180 145.550 49.400 145.690 ;
        RECT 42.180 145.490 42.500 145.550 ;
        RECT 45.860 145.490 46.180 145.550 ;
        RECT 49.080 145.490 49.400 145.550 ;
        RECT 53.220 145.490 53.540 145.750 ;
        RECT 54.140 145.490 54.460 145.750 ;
        RECT 62.880 145.490 63.200 145.750 ;
        RECT 85.420 145.490 85.740 145.750 ;
        RECT 86.340 145.490 86.660 145.750 ;
        RECT 87.260 145.690 87.580 145.750 ;
        RECT 87.735 145.690 88.025 145.735 ;
        RECT 87.260 145.550 88.025 145.690 ;
        RECT 87.260 145.490 87.580 145.550 ;
        RECT 87.735 145.505 88.025 145.550 ;
        RECT 116.240 145.490 116.560 145.750 ;
        RECT 117.620 145.690 117.940 145.750 ;
        RECT 120.855 145.690 121.145 145.735 ;
        RECT 117.620 145.550 121.145 145.690 ;
        RECT 117.620 145.490 117.940 145.550 ;
        RECT 120.855 145.505 121.145 145.550 ;
        RECT 132.340 145.490 132.660 145.750 ;
        RECT 132.890 145.690 133.030 145.890 ;
        RECT 133.760 145.890 137.720 146.030 ;
        RECT 133.760 145.845 134.050 145.890 ;
        RECT 135.860 145.845 136.150 145.890 ;
        RECT 137.430 145.845 137.720 145.890 ;
        RECT 137.950 145.890 144.070 146.030 ;
        RECT 137.950 145.690 138.090 145.890 ;
        RECT 132.890 145.550 138.090 145.690 ;
        RECT 142.920 145.490 143.240 145.750 ;
        RECT 17.270 144.870 146.990 145.350 ;
        RECT 36.215 144.485 36.505 144.715 ;
        RECT 36.290 144.330 36.430 144.485 ;
        RECT 39.420 144.470 39.740 144.730 ;
        RECT 44.020 144.670 44.340 144.730 ;
        RECT 40.890 144.530 44.340 144.670 ;
        RECT 40.890 144.330 41.030 144.530 ;
        RECT 44.020 144.470 44.340 144.530 ;
        RECT 46.780 144.670 47.100 144.730 ;
        RECT 47.715 144.670 48.005 144.715 ;
        RECT 46.780 144.530 48.005 144.670 ;
        RECT 46.780 144.470 47.100 144.530 ;
        RECT 47.715 144.485 48.005 144.530 ;
        RECT 36.290 144.190 41.030 144.330 ;
        RECT 41.300 144.330 41.590 144.375 ;
        RECT 43.400 144.330 43.690 144.375 ;
        RECT 44.970 144.330 45.260 144.375 ;
        RECT 41.300 144.190 45.260 144.330 ;
        RECT 41.300 144.145 41.590 144.190 ;
        RECT 43.400 144.145 43.690 144.190 ;
        RECT 44.970 144.145 45.260 144.190 ;
        RECT 35.740 143.990 36.060 144.050 ;
        RECT 40.815 143.990 41.105 144.035 ;
        RECT 35.740 143.850 41.105 143.990 ;
        RECT 35.740 143.790 36.060 143.850 ;
        RECT 40.815 143.805 41.105 143.850 ;
        RECT 41.695 143.990 41.985 144.035 ;
        RECT 42.885 143.990 43.175 144.035 ;
        RECT 45.405 143.990 45.695 144.035 ;
        RECT 41.695 143.850 45.695 143.990 ;
        RECT 41.695 143.805 41.985 143.850 ;
        RECT 42.885 143.805 43.175 143.850 ;
        RECT 45.405 143.805 45.695 143.850 ;
        RECT 20.115 143.650 20.405 143.695 ;
        RECT 20.560 143.650 20.880 143.710 ;
        RECT 37.595 143.650 37.885 143.695 ;
        RECT 47.240 143.650 47.560 143.710 ;
        RECT 20.115 143.510 20.880 143.650 ;
        RECT 20.115 143.465 20.405 143.510 ;
        RECT 20.560 143.450 20.880 143.510 ;
        RECT 35.370 143.510 37.365 143.650 ;
        RECT 34.820 143.310 35.140 143.370 ;
        RECT 35.370 143.355 35.510 143.510 ;
        RECT 36.200 143.355 36.520 143.370 ;
        RECT 35.295 143.310 35.585 143.355 ;
        RECT 34.820 143.170 35.585 143.310 ;
        RECT 34.820 143.110 35.140 143.170 ;
        RECT 35.295 143.125 35.585 143.170 ;
        RECT 36.200 143.125 36.585 143.355 ;
        RECT 37.225 143.310 37.365 143.510 ;
        RECT 37.595 143.510 47.560 143.650 ;
        RECT 37.595 143.465 37.885 143.510 ;
        RECT 47.240 143.450 47.560 143.510 ;
        RECT 39.435 143.310 39.725 143.355 ;
        RECT 42.040 143.310 42.330 143.355 ;
        RECT 37.225 143.170 39.725 143.310 ;
        RECT 39.435 143.125 39.725 143.170 ;
        RECT 40.430 143.170 42.330 143.310 ;
        RECT 47.790 143.310 47.930 144.485 ;
        RECT 49.080 144.470 49.400 144.730 ;
        RECT 53.220 144.470 53.540 144.730 ;
        RECT 54.600 144.470 54.920 144.730 ;
        RECT 62.880 144.670 63.200 144.730 ;
        RECT 56.530 144.530 63.200 144.670 ;
        RECT 48.160 144.330 48.480 144.390 ;
        RECT 50.000 144.330 50.320 144.390 ;
        RECT 56.530 144.330 56.670 144.530 ;
        RECT 62.880 144.470 63.200 144.530 ;
        RECT 63.340 144.470 63.660 144.730 ;
        RECT 75.300 144.670 75.620 144.730 ;
        RECT 79.900 144.670 80.220 144.730 ;
        RECT 75.300 144.530 80.220 144.670 ;
        RECT 75.300 144.470 75.620 144.530 ;
        RECT 79.900 144.470 80.220 144.530 ;
        RECT 80.375 144.670 80.665 144.715 ;
        RECT 82.200 144.670 82.520 144.730 ;
        RECT 80.375 144.530 82.520 144.670 ;
        RECT 80.375 144.485 80.665 144.530 ;
        RECT 82.200 144.470 82.520 144.530 ;
        RECT 96.920 144.470 97.240 144.730 ;
        RECT 102.440 144.670 102.760 144.730 ;
        RECT 103.375 144.670 103.665 144.715 ;
        RECT 102.440 144.530 103.665 144.670 ;
        RECT 102.440 144.470 102.760 144.530 ;
        RECT 103.375 144.485 103.665 144.530 ;
        RECT 106.120 144.670 106.440 144.730 ;
        RECT 107.975 144.670 108.265 144.715 ;
        RECT 106.120 144.530 108.265 144.670 ;
        RECT 106.120 144.470 106.440 144.530 ;
        RECT 107.975 144.485 108.265 144.530 ;
        RECT 118.555 144.670 118.845 144.715 ;
        RECT 124.520 144.670 124.840 144.730 ;
        RECT 118.555 144.530 124.840 144.670 ;
        RECT 118.555 144.485 118.845 144.530 ;
        RECT 124.520 144.470 124.840 144.530 ;
        RECT 48.160 144.190 50.320 144.330 ;
        RECT 48.160 144.130 48.480 144.190 ;
        RECT 50.000 144.130 50.320 144.190 ;
        RECT 54.690 144.190 56.670 144.330 ;
        RECT 56.940 144.330 57.230 144.375 ;
        RECT 59.040 144.330 59.330 144.375 ;
        RECT 60.610 144.330 60.900 144.375 ;
        RECT 56.940 144.190 60.900 144.330 ;
        RECT 50.090 143.650 50.230 144.130 ;
        RECT 51.395 143.650 51.685 143.695 ;
        RECT 50.090 143.510 51.685 143.650 ;
        RECT 51.395 143.465 51.685 143.510 ;
        RECT 52.315 143.650 52.605 143.695 ;
        RECT 52.760 143.650 53.080 143.710 ;
        RECT 52.315 143.510 53.080 143.650 ;
        RECT 52.315 143.465 52.605 143.510 ;
        RECT 52.760 143.450 53.080 143.510 ;
        RECT 48.175 143.310 48.465 143.355 ;
        RECT 47.790 143.170 48.465 143.310 ;
        RECT 36.200 143.110 36.520 143.125 ;
        RECT 15.960 142.970 16.280 143.030 ;
        RECT 19.195 142.970 19.485 143.015 ;
        RECT 15.960 142.830 19.485 142.970 ;
        RECT 15.960 142.770 16.280 142.830 ;
        RECT 19.195 142.785 19.485 142.830 ;
        RECT 37.135 142.970 37.425 143.015 ;
        RECT 38.040 142.970 38.360 143.030 ;
        RECT 40.430 143.015 40.570 143.170 ;
        RECT 42.040 143.125 42.330 143.170 ;
        RECT 48.175 143.125 48.465 143.170 ;
        RECT 53.680 143.110 54.000 143.370 ;
        RECT 54.690 143.355 54.830 144.190 ;
        RECT 56.940 144.145 57.230 144.190 ;
        RECT 59.040 144.145 59.330 144.190 ;
        RECT 60.610 144.145 60.900 144.190 ;
        RECT 72.580 144.330 72.870 144.375 ;
        RECT 74.680 144.330 74.970 144.375 ;
        RECT 76.250 144.330 76.540 144.375 ;
        RECT 72.580 144.190 76.540 144.330 ;
        RECT 72.580 144.145 72.870 144.190 ;
        RECT 74.680 144.145 74.970 144.190 ;
        RECT 76.250 144.145 76.540 144.190 ;
        RECT 78.520 144.330 78.840 144.390 ;
        RECT 78.995 144.330 79.285 144.375 ;
        RECT 88.680 144.330 88.970 144.375 ;
        RECT 90.780 144.330 91.070 144.375 ;
        RECT 92.350 144.330 92.640 144.375 ;
        RECT 78.520 144.190 85.190 144.330 ;
        RECT 78.520 144.130 78.840 144.190 ;
        RECT 78.995 144.145 79.285 144.190 ;
        RECT 85.050 144.035 85.190 144.190 ;
        RECT 88.680 144.190 92.640 144.330 ;
        RECT 88.680 144.145 88.970 144.190 ;
        RECT 90.780 144.145 91.070 144.190 ;
        RECT 92.350 144.145 92.640 144.190 ;
        RECT 99.680 144.130 100.000 144.390 ;
        RECT 121.300 144.330 121.590 144.375 ;
        RECT 122.870 144.330 123.160 144.375 ;
        RECT 124.970 144.330 125.260 144.375 ;
        RECT 121.300 144.190 125.260 144.330 ;
        RECT 121.300 144.145 121.590 144.190 ;
        RECT 122.870 144.145 123.160 144.190 ;
        RECT 124.970 144.145 125.260 144.190 ;
        RECT 134.220 144.330 134.510 144.375 ;
        RECT 136.320 144.330 136.610 144.375 ;
        RECT 137.890 144.330 138.180 144.375 ;
        RECT 134.220 144.190 138.180 144.330 ;
        RECT 134.220 144.145 134.510 144.190 ;
        RECT 136.320 144.145 136.610 144.190 ;
        RECT 137.890 144.145 138.180 144.190 ;
        RECT 140.635 144.145 140.925 144.375 ;
        RECT 57.335 143.990 57.625 144.035 ;
        RECT 58.525 143.990 58.815 144.035 ;
        RECT 61.045 143.990 61.335 144.035 ;
        RECT 57.335 143.850 61.335 143.990 ;
        RECT 57.335 143.805 57.625 143.850 ;
        RECT 58.525 143.805 58.815 143.850 ;
        RECT 61.045 143.805 61.335 143.850 ;
        RECT 72.975 143.990 73.265 144.035 ;
        RECT 74.165 143.990 74.455 144.035 ;
        RECT 76.685 143.990 76.975 144.035 ;
        RECT 72.975 143.850 76.975 143.990 ;
        RECT 72.975 143.805 73.265 143.850 ;
        RECT 74.165 143.805 74.455 143.850 ;
        RECT 76.685 143.805 76.975 143.850 ;
        RECT 80.835 143.990 81.125 144.035 ;
        RECT 82.215 143.990 82.505 144.035 ;
        RECT 80.835 143.850 82.505 143.990 ;
        RECT 80.835 143.805 81.125 143.850 ;
        RECT 82.215 143.805 82.505 143.850 ;
        RECT 84.975 143.805 85.265 144.035 ;
        RECT 87.720 143.990 88.040 144.050 ;
        RECT 88.195 143.990 88.485 144.035 ;
        RECT 87.720 143.850 88.485 143.990 ;
        RECT 87.720 143.790 88.040 143.850 ;
        RECT 88.195 143.805 88.485 143.850 ;
        RECT 89.075 143.990 89.365 144.035 ;
        RECT 90.265 143.990 90.555 144.035 ;
        RECT 92.785 143.990 93.075 144.035 ;
        RECT 99.770 143.990 99.910 144.130 ;
        RECT 89.075 143.850 93.075 143.990 ;
        RECT 89.075 143.805 89.365 143.850 ;
        RECT 90.265 143.805 90.555 143.850 ;
        RECT 92.785 143.805 93.075 143.850 ;
        RECT 97.930 143.850 99.910 143.990 ;
        RECT 56.455 143.650 56.745 143.695 ;
        RECT 62.420 143.650 62.740 143.710 ;
        RECT 56.455 143.510 62.740 143.650 ;
        RECT 56.455 143.465 56.745 143.510 ;
        RECT 62.420 143.450 62.740 143.510 ;
        RECT 72.080 143.450 72.400 143.710 ;
        RECT 79.440 143.450 79.760 143.710 ;
        RECT 85.420 143.650 85.740 143.710 ;
        RECT 85.895 143.650 86.185 143.695 ;
        RECT 85.420 143.510 86.185 143.650 ;
        RECT 85.420 143.450 85.740 143.510 ;
        RECT 85.895 143.465 86.185 143.510 ;
        RECT 86.815 143.650 87.105 143.695 ;
        RECT 87.260 143.650 87.580 143.710 ;
        RECT 97.930 143.695 98.070 143.850 ;
        RECT 105.660 143.790 105.980 144.050 ;
        RECT 106.595 143.990 106.885 144.035 ;
        RECT 111.195 143.990 111.485 144.035 ;
        RECT 114.860 143.990 115.180 144.050 ;
        RECT 106.595 143.850 115.180 143.990 ;
        RECT 106.595 143.805 106.885 143.850 ;
        RECT 111.195 143.805 111.485 143.850 ;
        RECT 114.860 143.790 115.180 143.850 ;
        RECT 120.865 143.990 121.155 144.035 ;
        RECT 123.385 143.990 123.675 144.035 ;
        RECT 124.575 143.990 124.865 144.035 ;
        RECT 120.865 143.850 124.865 143.990 ;
        RECT 120.865 143.805 121.155 143.850 ;
        RECT 123.385 143.805 123.675 143.850 ;
        RECT 124.575 143.805 124.865 143.850 ;
        RECT 125.455 143.990 125.745 144.035 ;
        RECT 134.615 143.990 134.905 144.035 ;
        RECT 135.805 143.990 136.095 144.035 ;
        RECT 138.325 143.990 138.615 144.035 ;
        RECT 125.455 143.850 133.950 143.990 ;
        RECT 125.455 143.805 125.745 143.850 ;
        RECT 86.815 143.510 87.580 143.650 ;
        RECT 86.815 143.465 87.105 143.510 ;
        RECT 87.260 143.450 87.580 143.510 ;
        RECT 97.855 143.465 98.145 143.695 ;
        RECT 98.315 143.465 98.605 143.695 ;
        RECT 98.760 143.650 99.080 143.710 ;
        RECT 99.235 143.650 99.525 143.695 ;
        RECT 98.760 143.510 99.525 143.650 ;
        RECT 89.560 143.355 89.880 143.370 ;
        RECT 54.690 143.170 54.985 143.355 ;
        RECT 57.680 143.310 57.970 143.355 ;
        RECT 54.695 143.125 54.985 143.170 ;
        RECT 55.610 143.170 57.970 143.310 ;
        RECT 37.135 142.830 38.360 142.970 ;
        RECT 37.135 142.785 37.425 142.830 ;
        RECT 38.040 142.770 38.360 142.830 ;
        RECT 40.355 142.785 40.645 143.015 ;
        RECT 44.480 142.970 44.800 143.030 ;
        RECT 55.610 143.015 55.750 143.170 ;
        RECT 57.680 143.125 57.970 143.170 ;
        RECT 73.430 143.310 73.720 143.355 ;
        RECT 86.355 143.310 86.645 143.355 ;
        RECT 73.430 143.170 86.645 143.310 ;
        RECT 73.430 143.125 73.720 143.170 ;
        RECT 86.355 143.125 86.645 143.170 ;
        RECT 89.530 143.125 89.880 143.355 ;
        RECT 98.390 143.310 98.530 143.465 ;
        RECT 98.760 143.450 99.080 143.510 ;
        RECT 99.235 143.465 99.525 143.510 ;
        RECT 99.680 143.450 100.000 143.710 ;
        RECT 101.520 143.650 101.840 143.710 ;
        RECT 105.215 143.650 105.505 143.695 ;
        RECT 121.760 143.650 122.080 143.710 ;
        RECT 101.520 143.510 122.080 143.650 ;
        RECT 101.520 143.450 101.840 143.510 ;
        RECT 105.215 143.465 105.505 143.510 ;
        RECT 121.760 143.450 122.080 143.510 ;
        RECT 124.980 143.650 125.300 143.710 ;
        RECT 133.810 143.695 133.950 143.850 ;
        RECT 134.615 143.850 138.615 143.990 ;
        RECT 140.710 143.990 140.850 144.145 ;
        RECT 142.000 143.990 142.320 144.050 ;
        RECT 143.855 143.990 144.145 144.035 ;
        RECT 140.710 143.850 144.145 143.990 ;
        RECT 134.615 143.805 134.905 143.850 ;
        RECT 135.805 143.805 136.095 143.850 ;
        RECT 138.325 143.805 138.615 143.850 ;
        RECT 142.000 143.790 142.320 143.850 ;
        RECT 143.855 143.805 144.145 143.850 ;
        RECT 125.915 143.650 126.205 143.695 ;
        RECT 124.980 143.510 126.205 143.650 ;
        RECT 124.980 143.450 125.300 143.510 ;
        RECT 125.915 143.465 126.205 143.510 ;
        RECT 133.735 143.650 134.025 143.695 ;
        RECT 133.735 143.510 136.250 143.650 ;
        RECT 133.735 143.465 134.025 143.510 ;
        RECT 136.110 143.370 136.250 143.510 ;
        RECT 110.275 143.310 110.565 143.355 ;
        RECT 116.240 143.310 116.560 143.370 ;
        RECT 98.390 143.170 116.560 143.310 ;
        RECT 110.275 143.125 110.565 143.170 ;
        RECT 89.560 143.110 89.880 143.125 ;
        RECT 116.240 143.110 116.560 143.170 ;
        RECT 124.230 143.310 124.520 143.355 ;
        RECT 128.200 143.310 128.520 143.370 ;
        RECT 124.230 143.170 128.520 143.310 ;
        RECT 124.230 143.125 124.520 143.170 ;
        RECT 128.200 143.110 128.520 143.170 ;
        RECT 134.180 143.310 134.500 143.370 ;
        RECT 134.960 143.310 135.250 143.355 ;
        RECT 134.180 143.170 135.250 143.310 ;
        RECT 134.180 143.110 134.500 143.170 ;
        RECT 134.960 143.125 135.250 143.170 ;
        RECT 136.020 143.110 136.340 143.370 ;
        RECT 49.175 142.970 49.465 143.015 ;
        RECT 44.480 142.830 49.465 142.970 ;
        RECT 44.480 142.770 44.800 142.830 ;
        RECT 49.175 142.785 49.465 142.830 ;
        RECT 55.535 142.785 55.825 143.015 ;
        RECT 95.080 142.770 95.400 143.030 ;
        RECT 109.815 142.970 110.105 143.015 ;
        RECT 113.940 142.970 114.260 143.030 ;
        RECT 122.220 142.970 122.540 143.030 ;
        RECT 109.815 142.830 122.540 142.970 ;
        RECT 109.815 142.785 110.105 142.830 ;
        RECT 113.940 142.770 114.260 142.830 ;
        RECT 122.220 142.770 122.540 142.830 ;
        RECT 129.135 142.970 129.425 143.015 ;
        RECT 130.500 142.970 130.820 143.030 ;
        RECT 129.135 142.830 130.820 142.970 ;
        RECT 129.135 142.785 129.425 142.830 ;
        RECT 130.500 142.770 130.820 142.830 ;
        RECT 141.080 142.770 141.400 143.030 ;
        RECT 17.270 142.150 146.990 142.630 ;
        RECT 42.180 141.950 42.500 142.010 ;
        RECT 42.655 141.950 42.945 141.995 ;
        RECT 42.180 141.810 42.945 141.950 ;
        RECT 42.180 141.750 42.500 141.810 ;
        RECT 42.655 141.765 42.945 141.810 ;
        RECT 22.860 141.610 23.180 141.670 ;
        RECT 28.395 141.610 28.685 141.655 ;
        RECT 22.860 141.470 28.685 141.610 ;
        RECT 22.860 141.410 23.180 141.470 ;
        RECT 28.395 141.425 28.685 141.470 ;
        RECT 37.090 141.610 37.380 141.655 ;
        RECT 38.040 141.610 38.360 141.670 ;
        RECT 37.090 141.470 38.360 141.610 ;
        RECT 37.090 141.425 37.380 141.470 ;
        RECT 38.040 141.410 38.360 141.470 ;
        RECT 18.720 141.270 19.040 141.330 ;
        RECT 20.475 141.270 20.765 141.315 ;
        RECT 18.720 141.130 20.765 141.270 ;
        RECT 18.720 141.070 19.040 141.130 ;
        RECT 20.475 141.085 20.765 141.130 ;
        RECT 27.475 141.270 27.765 141.315 ;
        RECT 27.920 141.270 28.240 141.330 ;
        RECT 27.475 141.130 28.240 141.270 ;
        RECT 27.475 141.085 27.765 141.130 ;
        RECT 27.920 141.070 28.240 141.130 ;
        RECT 35.740 141.070 36.060 141.330 ;
        RECT 42.730 141.270 42.870 141.765 ;
        RECT 44.020 141.750 44.340 142.010 ;
        RECT 51.395 141.950 51.685 141.995 ;
        RECT 52.760 141.950 53.080 142.010 ;
        RECT 51.395 141.810 53.080 141.950 ;
        RECT 51.395 141.765 51.685 141.810 ;
        RECT 52.760 141.750 53.080 141.810 ;
        RECT 78.060 141.750 78.380 142.010 ;
        RECT 85.435 141.950 85.725 141.995 ;
        RECT 87.355 141.950 87.645 141.995 ;
        RECT 85.435 141.810 87.645 141.950 ;
        RECT 85.435 141.765 85.725 141.810 ;
        RECT 87.355 141.765 87.645 141.810 ;
        RECT 89.115 141.950 89.405 141.995 ;
        RECT 89.560 141.950 89.880 142.010 ;
        RECT 89.115 141.810 89.880 141.950 ;
        RECT 89.115 141.765 89.405 141.810 ;
        RECT 89.560 141.750 89.880 141.810 ;
        RECT 90.955 141.950 91.245 141.995 ;
        RECT 95.080 141.950 95.400 142.010 ;
        RECT 105.200 141.950 105.520 142.010 ;
        RECT 90.955 141.810 105.520 141.950 ;
        RECT 90.955 141.765 91.245 141.810 ;
        RECT 95.080 141.750 95.400 141.810 ;
        RECT 105.200 141.750 105.520 141.810 ;
        RECT 120.380 141.950 120.700 142.010 ;
        RECT 120.855 141.950 121.145 141.995 ;
        RECT 120.380 141.810 121.145 141.950 ;
        RECT 120.380 141.750 120.700 141.810 ;
        RECT 120.855 141.765 121.145 141.810 ;
        RECT 128.200 141.750 128.520 142.010 ;
        RECT 133.735 141.950 134.025 141.995 ;
        RECT 134.180 141.950 134.500 142.010 ;
        RECT 133.735 141.810 134.500 141.950 ;
        RECT 133.735 141.765 134.025 141.810 ;
        RECT 134.180 141.750 134.500 141.810 ;
        RECT 135.575 141.950 135.865 141.995 ;
        RECT 141.080 141.950 141.400 142.010 ;
        RECT 135.575 141.810 141.400 141.950 ;
        RECT 135.575 141.765 135.865 141.810 ;
        RECT 141.080 141.750 141.400 141.810 ;
        RECT 142.935 141.765 143.225 141.995 ;
        RECT 54.140 141.610 54.460 141.670 ;
        RECT 56.960 141.610 57.250 141.655 ;
        RECT 54.140 141.470 57.250 141.610 ;
        RECT 54.140 141.410 54.460 141.470 ;
        RECT 56.960 141.425 57.250 141.470 ;
        RECT 77.140 141.410 77.460 141.670 ;
        RECT 85.880 141.610 86.200 141.670 ;
        RECT 86.355 141.610 86.645 141.655 ;
        RECT 78.610 141.470 86.645 141.610 ;
        RECT 43.575 141.270 43.865 141.315 ;
        RECT 42.730 141.130 43.865 141.270 ;
        RECT 43.575 141.085 43.865 141.130 ;
        RECT 44.480 141.070 44.800 141.330 ;
        RECT 58.295 141.270 58.585 141.315 ;
        RECT 65.655 141.270 65.945 141.315 ;
        RECT 58.295 141.130 65.945 141.270 ;
        RECT 58.295 141.085 58.585 141.130 ;
        RECT 65.655 141.085 65.945 141.130 ;
        RECT 66.560 141.270 66.880 141.330 ;
        RECT 78.610 141.315 78.750 141.470 ;
        RECT 85.880 141.410 86.200 141.470 ;
        RECT 86.355 141.425 86.645 141.470 ;
        RECT 104.280 141.610 104.600 141.670 ;
        RECT 110.735 141.610 111.025 141.655 ;
        RECT 136.020 141.610 136.340 141.670 ;
        RECT 104.280 141.470 111.025 141.610 ;
        RECT 104.280 141.410 104.600 141.470 ;
        RECT 110.735 141.425 111.025 141.470 ;
        RECT 127.830 141.470 136.340 141.610 ;
        RECT 69.335 141.270 69.625 141.315 ;
        RECT 66.560 141.130 69.625 141.270 ;
        RECT 19.180 140.730 19.500 140.990 ;
        RECT 20.075 140.930 20.365 140.975 ;
        RECT 21.265 140.930 21.555 140.975 ;
        RECT 23.785 140.930 24.075 140.975 ;
        RECT 20.075 140.790 24.075 140.930 ;
        RECT 20.075 140.745 20.365 140.790 ;
        RECT 21.265 140.745 21.555 140.790 ;
        RECT 23.785 140.745 24.075 140.790 ;
        RECT 36.635 140.930 36.925 140.975 ;
        RECT 37.825 140.930 38.115 140.975 ;
        RECT 40.345 140.930 40.635 140.975 ;
        RECT 36.635 140.790 40.635 140.930 ;
        RECT 36.635 140.745 36.925 140.790 ;
        RECT 37.825 140.745 38.115 140.790 ;
        RECT 40.345 140.745 40.635 140.790 ;
        RECT 41.720 140.930 42.040 140.990 ;
        RECT 44.570 140.930 44.710 141.070 ;
        RECT 41.720 140.790 44.710 140.930 ;
        RECT 53.705 140.930 53.995 140.975 ;
        RECT 56.225 140.930 56.515 140.975 ;
        RECT 57.415 140.930 57.705 140.975 ;
        RECT 53.705 140.790 57.705 140.930 ;
        RECT 65.730 140.930 65.870 141.085 ;
        RECT 66.560 141.070 66.880 141.130 ;
        RECT 69.335 141.085 69.625 141.130 ;
        RECT 78.075 141.085 78.365 141.315 ;
        RECT 78.535 141.085 78.825 141.315 ;
        RECT 82.660 141.270 82.980 141.330 ;
        RECT 84.975 141.270 85.265 141.315 ;
        RECT 85.420 141.270 85.740 141.330 ;
        RECT 87.260 141.270 87.580 141.330 ;
        RECT 82.660 141.130 87.580 141.270 ;
        RECT 69.780 140.930 70.100 140.990 ;
        RECT 73.015 140.930 73.305 140.975 ;
        RECT 65.730 140.790 73.305 140.930 ;
        RECT 41.720 140.730 42.040 140.790 ;
        RECT 53.705 140.745 53.995 140.790 ;
        RECT 56.225 140.745 56.515 140.790 ;
        RECT 57.415 140.745 57.705 140.790 ;
        RECT 69.780 140.730 70.100 140.790 ;
        RECT 73.015 140.745 73.305 140.790 ;
        RECT 76.220 140.930 76.540 140.990 ;
        RECT 78.150 140.930 78.290 141.085 ;
        RECT 82.660 141.070 82.980 141.130 ;
        RECT 84.975 141.085 85.265 141.130 ;
        RECT 85.420 141.070 85.740 141.130 ;
        RECT 87.260 141.070 87.580 141.130 ;
        RECT 108.895 141.270 109.185 141.315 ;
        RECT 109.340 141.270 109.660 141.330 ;
        RECT 108.895 141.130 109.660 141.270 ;
        RECT 108.895 141.085 109.185 141.130 ;
        RECT 109.340 141.070 109.660 141.130 ;
        RECT 112.575 141.270 112.865 141.315 ;
        RECT 113.480 141.270 113.800 141.330 ;
        RECT 112.575 141.130 113.800 141.270 ;
        RECT 112.575 141.085 112.865 141.130 ;
        RECT 113.480 141.070 113.800 141.130 ;
        RECT 117.620 141.070 117.940 141.330 ;
        RECT 127.830 141.315 127.970 141.470 ;
        RECT 136.020 141.410 136.340 141.470 ;
        RECT 139.240 141.610 139.560 141.670 ;
        RECT 139.715 141.610 140.005 141.655 ;
        RECT 139.240 141.470 140.005 141.610 ;
        RECT 139.240 141.410 139.560 141.470 ;
        RECT 139.715 141.425 140.005 141.470 ;
        RECT 119.015 141.085 119.305 141.315 ;
        RECT 119.935 141.270 120.225 141.315 ;
        RECT 126.420 141.270 126.710 141.315 ;
        RECT 119.935 141.130 126.710 141.270 ;
        RECT 119.935 141.085 120.225 141.130 ;
        RECT 126.420 141.085 126.710 141.130 ;
        RECT 127.755 141.085 128.045 141.315 ;
        RECT 76.220 140.790 78.290 140.930 ;
        RECT 81.740 140.930 82.060 140.990 ;
        RECT 86.340 140.930 86.660 140.990 ;
        RECT 90.020 140.930 90.340 140.990 ;
        RECT 91.415 140.930 91.705 140.975 ;
        RECT 81.740 140.790 91.705 140.930 ;
        RECT 76.220 140.730 76.540 140.790 ;
        RECT 81.740 140.730 82.060 140.790 ;
        RECT 86.340 140.730 86.660 140.790 ;
        RECT 90.020 140.730 90.340 140.790 ;
        RECT 91.415 140.745 91.705 140.790 ;
        RECT 91.875 140.745 92.165 140.975 ;
        RECT 19.680 140.590 19.970 140.635 ;
        RECT 21.780 140.590 22.070 140.635 ;
        RECT 23.350 140.590 23.640 140.635 ;
        RECT 19.680 140.450 23.640 140.590 ;
        RECT 19.680 140.405 19.970 140.450 ;
        RECT 21.780 140.405 22.070 140.450 ;
        RECT 23.350 140.405 23.640 140.450 ;
        RECT 36.240 140.590 36.530 140.635 ;
        RECT 38.340 140.590 38.630 140.635 ;
        RECT 39.910 140.590 40.200 140.635 ;
        RECT 36.240 140.450 40.200 140.590 ;
        RECT 36.240 140.405 36.530 140.450 ;
        RECT 38.340 140.405 38.630 140.450 ;
        RECT 39.910 140.405 40.200 140.450 ;
        RECT 54.140 140.590 54.430 140.635 ;
        RECT 55.710 140.590 56.000 140.635 ;
        RECT 57.810 140.590 58.100 140.635 ;
        RECT 54.140 140.450 58.100 140.590 ;
        RECT 54.140 140.405 54.430 140.450 ;
        RECT 55.710 140.405 56.000 140.450 ;
        RECT 57.810 140.405 58.100 140.450 ;
        RECT 88.195 140.590 88.485 140.635 ;
        RECT 91.950 140.590 92.090 140.745 ;
        RECT 102.440 140.730 102.760 140.990 ;
        RECT 110.260 140.730 110.580 140.990 ;
        RECT 119.090 140.930 119.230 141.085 ;
        RECT 129.120 141.070 129.440 141.330 ;
        RECT 130.500 141.070 130.820 141.330 ;
        RECT 135.560 141.270 135.880 141.330 ;
        RECT 135.560 141.130 139.470 141.270 ;
        RECT 135.560 141.070 135.880 141.130 ;
        RECT 122.220 140.930 122.540 140.990 ;
        RECT 119.090 140.790 122.540 140.930 ;
        RECT 122.220 140.730 122.540 140.790 ;
        RECT 123.165 140.930 123.455 140.975 ;
        RECT 125.685 140.930 125.975 140.975 ;
        RECT 126.875 140.930 127.165 140.975 ;
        RECT 123.165 140.790 127.165 140.930 ;
        RECT 123.165 140.745 123.455 140.790 ;
        RECT 125.685 140.745 125.975 140.790 ;
        RECT 126.875 140.745 127.165 140.790 ;
        RECT 132.340 140.930 132.660 140.990 ;
        RECT 136.035 140.930 136.325 140.975 ;
        RECT 132.340 140.790 136.325 140.930 ;
        RECT 132.340 140.730 132.660 140.790 ;
        RECT 136.035 140.745 136.325 140.790 ;
        RECT 136.495 140.745 136.785 140.975 ;
        RECT 139.330 140.930 139.470 141.130 ;
        RECT 142.000 141.070 142.320 141.330 ;
        RECT 143.010 141.270 143.150 141.765 ;
        RECT 143.855 141.270 144.145 141.315 ;
        RECT 143.010 141.130 144.145 141.270 ;
        RECT 143.855 141.085 144.145 141.130 ;
        RECT 140.175 140.930 140.465 140.975 ;
        RECT 139.330 140.790 140.465 140.930 ;
        RECT 140.175 140.745 140.465 140.790 ;
        RECT 88.195 140.450 92.090 140.590 ;
        RECT 103.820 140.590 104.140 140.650 ;
        RECT 109.815 140.590 110.105 140.635 ;
        RECT 118.095 140.590 118.385 140.635 ;
        RECT 118.540 140.590 118.860 140.650 ;
        RECT 103.820 140.450 118.860 140.590 ;
        RECT 88.195 140.405 88.485 140.450 ;
        RECT 103.820 140.390 104.140 140.450 ;
        RECT 109.815 140.405 110.105 140.450 ;
        RECT 118.095 140.405 118.385 140.450 ;
        RECT 118.540 140.390 118.860 140.450 ;
        RECT 123.600 140.590 123.890 140.635 ;
        RECT 125.170 140.590 125.460 140.635 ;
        RECT 127.270 140.590 127.560 140.635 ;
        RECT 130.055 140.590 130.345 140.635 ;
        RECT 123.600 140.450 127.560 140.590 ;
        RECT 123.600 140.405 123.890 140.450 ;
        RECT 125.170 140.405 125.460 140.450 ;
        RECT 127.270 140.405 127.560 140.450 ;
        RECT 127.830 140.450 130.345 140.590 ;
        RECT 20.560 140.250 20.880 140.310 ;
        RECT 26.095 140.250 26.385 140.295 ;
        RECT 20.560 140.110 26.385 140.250 ;
        RECT 20.560 140.050 20.880 140.110 ;
        RECT 26.095 140.065 26.385 140.110 ;
        RECT 29.315 140.250 29.605 140.295 ;
        RECT 31.140 140.250 31.460 140.310 ;
        RECT 29.315 140.110 31.460 140.250 ;
        RECT 29.315 140.065 29.605 140.110 ;
        RECT 31.140 140.050 31.460 140.110 ;
        RECT 87.260 140.050 87.580 140.310 ;
        RECT 105.675 140.250 105.965 140.295 ;
        RECT 107.040 140.250 107.360 140.310 ;
        RECT 105.675 140.110 107.360 140.250 ;
        RECT 105.675 140.065 105.965 140.110 ;
        RECT 107.040 140.050 107.360 140.110 ;
        RECT 107.975 140.250 108.265 140.295 ;
        RECT 108.420 140.250 108.740 140.310 ;
        RECT 107.975 140.110 108.740 140.250 ;
        RECT 118.630 140.250 118.770 140.390 ;
        RECT 127.830 140.250 127.970 140.450 ;
        RECT 130.055 140.405 130.345 140.450 ;
        RECT 135.100 140.590 135.420 140.650 ;
        RECT 136.570 140.590 136.710 140.745 ;
        RECT 135.100 140.450 136.710 140.590 ;
        RECT 140.250 140.590 140.390 140.745 ;
        RECT 140.620 140.730 140.940 140.990 ;
        RECT 144.300 140.590 144.620 140.650 ;
        RECT 140.250 140.450 144.620 140.590 ;
        RECT 135.100 140.390 135.420 140.450 ;
        RECT 144.300 140.390 144.620 140.450 ;
        RECT 144.760 140.390 145.080 140.650 ;
        RECT 118.630 140.110 127.970 140.250 ;
        RECT 132.340 140.250 132.660 140.310 ;
        RECT 137.875 140.250 138.165 140.295 ;
        RECT 132.340 140.110 138.165 140.250 ;
        RECT 107.975 140.065 108.265 140.110 ;
        RECT 108.420 140.050 108.740 140.110 ;
        RECT 132.340 140.050 132.660 140.110 ;
        RECT 137.875 140.065 138.165 140.110 ;
        RECT 17.270 139.430 146.990 139.910 ;
        RECT 18.720 139.030 19.040 139.290 ;
        RECT 22.860 139.030 23.180 139.290 ;
        RECT 27.920 139.230 28.240 139.290 ;
        RECT 31.600 139.230 31.920 139.290 ;
        RECT 24.790 139.090 31.920 139.230 ;
        RECT 21.955 138.550 22.245 138.595 ;
        RECT 24.790 138.550 24.930 139.090 ;
        RECT 27.920 139.030 28.240 139.090 ;
        RECT 31.600 139.030 31.920 139.090 ;
        RECT 72.095 139.230 72.385 139.275 ;
        RECT 72.540 139.230 72.860 139.290 ;
        RECT 72.095 139.090 72.860 139.230 ;
        RECT 72.095 139.045 72.385 139.090 ;
        RECT 72.540 139.030 72.860 139.090 ;
        RECT 73.015 139.230 73.305 139.275 ;
        RECT 76.220 139.230 76.540 139.290 ;
        RECT 82.675 139.230 82.965 139.275 ;
        RECT 73.015 139.090 82.965 139.230 ;
        RECT 73.015 139.045 73.305 139.090 ;
        RECT 76.220 139.030 76.540 139.090 ;
        RECT 82.675 139.045 82.965 139.090 ;
        RECT 25.620 138.890 25.910 138.935 ;
        RECT 27.190 138.890 27.480 138.935 ;
        RECT 29.290 138.890 29.580 138.935 ;
        RECT 25.620 138.750 29.580 138.890 ;
        RECT 25.620 138.705 25.910 138.750 ;
        RECT 27.190 138.705 27.480 138.750 ;
        RECT 29.290 138.705 29.580 138.750 ;
        RECT 32.075 138.890 32.365 138.935 ;
        RECT 32.520 138.890 32.840 138.950 ;
        RECT 73.460 138.890 73.780 138.950 ;
        RECT 32.075 138.750 32.840 138.890 ;
        RECT 32.075 138.705 32.365 138.750 ;
        RECT 32.520 138.690 32.840 138.750 ;
        RECT 69.870 138.750 73.780 138.890 ;
        RECT 21.955 138.410 24.930 138.550 ;
        RECT 25.185 138.550 25.475 138.595 ;
        RECT 27.705 138.550 27.995 138.595 ;
        RECT 28.895 138.550 29.185 138.595 ;
        RECT 25.185 138.410 29.185 138.550 ;
        RECT 21.955 138.365 22.245 138.410 ;
        RECT 25.185 138.365 25.475 138.410 ;
        RECT 27.705 138.365 27.995 138.410 ;
        RECT 28.895 138.365 29.185 138.410 ;
        RECT 31.140 138.550 31.460 138.610 ;
        RECT 31.140 138.410 33.210 138.550 ;
        RECT 31.140 138.350 31.460 138.410 ;
        RECT 20.560 138.010 20.880 138.270 ;
        RECT 24.700 138.210 25.020 138.270 ;
        RECT 29.775 138.210 30.065 138.255 ;
        RECT 24.700 138.070 30.065 138.210 ;
        RECT 24.700 138.010 25.020 138.070 ;
        RECT 29.775 138.025 30.065 138.070 ;
        RECT 30.220 138.210 30.540 138.270 ;
        RECT 33.070 138.255 33.210 138.410 ;
        RECT 69.870 138.255 70.010 138.750 ;
        RECT 73.460 138.690 73.780 138.750 ;
        RECT 70.240 138.350 70.560 138.610 ;
        RECT 71.635 138.550 71.925 138.595 ;
        RECT 73.920 138.550 74.240 138.610 ;
        RECT 71.635 138.410 74.240 138.550 ;
        RECT 82.750 138.550 82.890 139.045 ;
        RECT 85.420 139.030 85.740 139.290 ;
        RECT 103.820 139.230 104.140 139.290 ;
        RECT 106.595 139.230 106.885 139.275 ;
        RECT 87.350 139.090 91.630 139.230 ;
        RECT 84.515 138.890 84.805 138.935 ;
        RECT 87.350 138.890 87.490 139.090 ;
        RECT 84.515 138.750 87.490 138.890 ;
        RECT 87.735 138.890 88.025 138.935 ;
        RECT 87.735 138.750 91.170 138.890 ;
        RECT 84.515 138.705 84.805 138.750 ;
        RECT 87.735 138.705 88.025 138.750 ;
        RECT 86.355 138.550 86.645 138.595 ;
        RECT 87.260 138.550 87.580 138.610 ;
        RECT 91.030 138.595 91.170 138.750 ;
        RECT 82.750 138.410 87.580 138.550 ;
        RECT 71.635 138.365 71.925 138.410 ;
        RECT 73.920 138.350 74.240 138.410 ;
        RECT 86.355 138.365 86.645 138.410 ;
        RECT 87.260 138.350 87.580 138.410 ;
        RECT 90.955 138.365 91.245 138.595 ;
        RECT 91.490 138.550 91.630 139.090 ;
        RECT 103.820 139.090 106.885 139.230 ;
        RECT 103.820 139.030 104.140 139.090 ;
        RECT 106.595 139.045 106.885 139.090 ;
        RECT 110.260 139.030 110.580 139.290 ;
        RECT 119.920 139.230 120.240 139.290 ;
        RECT 127.280 139.230 127.600 139.290 ;
        RECT 128.215 139.230 128.505 139.275 ;
        RECT 119.920 139.090 128.505 139.230 ;
        RECT 119.920 139.030 120.240 139.090 ;
        RECT 127.280 139.030 127.600 139.090 ;
        RECT 128.215 139.045 128.505 139.090 ;
        RECT 129.120 139.230 129.440 139.290 ;
        RECT 133.735 139.230 134.025 139.275 ;
        RECT 129.120 139.090 134.025 139.230 ;
        RECT 129.120 139.030 129.440 139.090 ;
        RECT 133.735 139.045 134.025 139.090 ;
        RECT 135.650 139.090 137.630 139.230 ;
        RECT 98.760 138.890 99.080 138.950 ;
        RECT 103.360 138.890 103.680 138.950 ;
        RECT 98.760 138.750 103.680 138.890 ;
        RECT 98.760 138.690 99.080 138.750 ;
        RECT 103.360 138.690 103.680 138.750 ;
        RECT 114.440 138.890 114.730 138.935 ;
        RECT 116.540 138.890 116.830 138.935 ;
        RECT 118.110 138.890 118.400 138.935 ;
        RECT 114.440 138.750 118.400 138.890 ;
        RECT 114.440 138.705 114.730 138.750 ;
        RECT 116.540 138.705 116.830 138.750 ;
        RECT 118.110 138.705 118.400 138.750 ;
        RECT 120.840 138.690 121.160 138.950 ;
        RECT 121.800 138.890 122.090 138.935 ;
        RECT 123.900 138.890 124.190 138.935 ;
        RECT 125.470 138.890 125.760 138.935 ;
        RECT 121.800 138.750 125.760 138.890 ;
        RECT 121.800 138.705 122.090 138.750 ;
        RECT 123.900 138.705 124.190 138.750 ;
        RECT 125.470 138.705 125.760 138.750 ;
        RECT 132.340 138.690 132.660 138.950 ;
        RECT 132.815 138.890 133.105 138.935 ;
        RECT 135.650 138.890 135.790 139.090 ;
        RECT 132.815 138.750 135.790 138.890 ;
        RECT 132.815 138.705 133.105 138.750 ;
        RECT 136.480 138.690 136.800 138.950 ;
        RECT 95.095 138.550 95.385 138.595 ;
        RECT 91.490 138.410 95.385 138.550 ;
        RECT 95.095 138.365 95.385 138.410 ;
        RECT 100.140 138.550 100.460 138.610 ;
        RECT 100.140 138.410 103.590 138.550 ;
        RECT 100.140 138.350 100.460 138.410 ;
        RECT 31.615 138.210 31.905 138.255 ;
        RECT 30.220 138.070 31.905 138.210 ;
        RECT 30.220 138.010 30.540 138.070 ;
        RECT 31.615 138.025 31.905 138.070 ;
        RECT 32.535 138.025 32.825 138.255 ;
        RECT 32.995 138.025 33.285 138.255 ;
        RECT 69.795 138.025 70.085 138.255 ;
        RECT 74.855 138.210 75.145 138.255 ;
        RECT 77.140 138.210 77.460 138.270 ;
        RECT 74.855 138.070 77.460 138.210 ;
        RECT 74.855 138.025 75.145 138.070 ;
        RECT 21.035 137.870 21.325 137.915 ;
        RECT 24.240 137.870 24.560 137.930 ;
        RECT 21.035 137.730 24.560 137.870 ;
        RECT 21.035 137.685 21.325 137.730 ;
        RECT 24.240 137.670 24.560 137.730 ;
        RECT 28.550 137.870 28.840 137.915 ;
        RECT 30.695 137.870 30.985 137.915 ;
        RECT 28.550 137.730 30.985 137.870 ;
        RECT 28.550 137.685 28.840 137.730 ;
        RECT 30.695 137.685 30.985 137.730 ;
        RECT 31.140 137.870 31.460 137.930 ;
        RECT 32.610 137.870 32.750 138.025 ;
        RECT 77.140 138.010 77.460 138.070 ;
        RECT 82.660 138.010 82.980 138.270 ;
        RECT 83.595 138.210 83.885 138.255 ;
        RECT 84.975 138.210 85.265 138.255 ;
        RECT 85.880 138.210 86.200 138.270 ;
        RECT 83.595 138.070 86.200 138.210 ;
        RECT 83.595 138.025 83.885 138.070 ;
        RECT 84.975 138.025 85.265 138.070 ;
        RECT 85.880 138.010 86.200 138.070 ;
        RECT 90.020 138.010 90.340 138.270 ;
        RECT 93.240 138.210 93.560 138.270 ;
        RECT 103.450 138.255 103.590 138.410 ;
        RECT 107.040 138.350 107.360 138.610 ;
        RECT 112.560 138.550 112.880 138.610 ;
        RECT 113.035 138.550 113.325 138.595 ;
        RECT 112.560 138.410 113.325 138.550 ;
        RECT 112.560 138.350 112.880 138.410 ;
        RECT 113.035 138.365 113.325 138.410 ;
        RECT 114.835 138.550 115.125 138.595 ;
        RECT 116.025 138.550 116.315 138.595 ;
        RECT 118.545 138.550 118.835 138.595 ;
        RECT 114.835 138.410 118.835 138.550 ;
        RECT 114.835 138.365 115.125 138.410 ;
        RECT 116.025 138.365 116.315 138.410 ;
        RECT 118.545 138.365 118.835 138.410 ;
        RECT 122.195 138.550 122.485 138.595 ;
        RECT 123.385 138.550 123.675 138.595 ;
        RECT 125.905 138.550 126.195 138.595 ;
        RECT 122.195 138.410 126.195 138.550 ;
        RECT 122.195 138.365 122.485 138.410 ;
        RECT 123.385 138.365 123.675 138.410 ;
        RECT 125.905 138.365 126.195 138.410 ;
        RECT 130.040 138.550 130.360 138.610 ;
        RECT 130.515 138.550 130.805 138.595 ;
        RECT 136.570 138.550 136.710 138.690 ;
        RECT 130.040 138.410 130.805 138.550 ;
        RECT 130.040 138.350 130.360 138.410 ;
        RECT 130.515 138.365 130.805 138.410 ;
        RECT 136.110 138.410 136.710 138.550 ;
        RECT 137.490 138.550 137.630 139.090 ;
        RECT 144.300 139.030 144.620 139.290 ;
        RECT 137.900 138.890 138.190 138.935 ;
        RECT 140.000 138.890 140.290 138.935 ;
        RECT 141.570 138.890 141.860 138.935 ;
        RECT 137.900 138.750 141.860 138.890 ;
        RECT 137.900 138.705 138.190 138.750 ;
        RECT 140.000 138.705 140.290 138.750 ;
        RECT 141.570 138.705 141.860 138.750 ;
        RECT 138.295 138.550 138.585 138.595 ;
        RECT 139.485 138.550 139.775 138.595 ;
        RECT 142.005 138.550 142.295 138.595 ;
        RECT 137.490 138.410 138.090 138.550 ;
        RECT 101.535 138.210 101.825 138.255 ;
        RECT 93.240 138.070 101.825 138.210 ;
        RECT 93.240 138.010 93.560 138.070 ;
        RECT 101.535 138.025 101.825 138.070 ;
        RECT 102.455 138.025 102.745 138.255 ;
        RECT 103.375 138.210 103.665 138.255 ;
        RECT 104.280 138.210 104.600 138.270 ;
        RECT 103.375 138.070 104.600 138.210 ;
        RECT 103.375 138.025 103.665 138.070 ;
        RECT 31.140 137.730 32.750 137.870 ;
        RECT 66.560 137.870 66.880 137.930 ;
        RECT 86.800 137.870 87.120 137.930 ;
        RECT 89.560 137.870 89.880 137.930 ;
        RECT 66.560 137.730 89.880 137.870 ;
        RECT 90.110 137.870 90.250 138.010 ;
        RECT 94.175 137.870 94.465 137.915 ;
        RECT 90.110 137.730 94.465 137.870 ;
        RECT 102.530 137.870 102.670 138.025 ;
        RECT 104.280 138.010 104.600 138.070 ;
        RECT 105.660 138.010 105.980 138.270 ;
        RECT 111.640 138.210 111.960 138.270 ;
        RECT 113.955 138.210 114.245 138.255 ;
        RECT 120.840 138.210 121.160 138.270 ;
        RECT 121.315 138.210 121.605 138.255 ;
        RECT 111.640 138.070 131.650 138.210 ;
        RECT 111.640 138.010 111.960 138.070 ;
        RECT 113.955 138.025 114.245 138.070 ;
        RECT 120.840 138.010 121.160 138.070 ;
        RECT 121.315 138.025 121.605 138.070 ;
        RECT 114.400 137.870 114.720 137.930 ;
        RECT 102.530 137.730 114.720 137.870 ;
        RECT 31.140 137.670 31.460 137.730 ;
        RECT 66.560 137.670 66.880 137.730 ;
        RECT 86.800 137.670 87.120 137.730 ;
        RECT 89.560 137.670 89.880 137.730 ;
        RECT 94.175 137.685 94.465 137.730 ;
        RECT 114.400 137.670 114.720 137.730 ;
        RECT 115.290 137.870 115.580 137.915 ;
        RECT 116.700 137.870 117.020 137.930 ;
        RECT 122.680 137.915 123.000 137.930 ;
        RECT 115.290 137.730 117.020 137.870 ;
        RECT 115.290 137.685 115.580 137.730 ;
        RECT 116.700 137.670 117.020 137.730 ;
        RECT 122.650 137.685 123.000 137.915 ;
        RECT 131.510 137.870 131.650 138.070 ;
        RECT 134.640 138.010 134.960 138.270 ;
        RECT 135.115 138.210 135.405 138.255 ;
        RECT 135.560 138.210 135.880 138.270 ;
        RECT 136.110 138.255 136.250 138.410 ;
        RECT 135.115 138.070 135.880 138.210 ;
        RECT 135.115 138.025 135.405 138.070 ;
        RECT 135.560 138.010 135.880 138.070 ;
        RECT 136.035 138.025 136.325 138.255 ;
        RECT 136.495 138.210 136.785 138.255 ;
        RECT 136.940 138.210 137.260 138.270 ;
        RECT 136.495 138.070 137.260 138.210 ;
        RECT 136.495 138.025 136.785 138.070 ;
        RECT 136.940 138.010 137.260 138.070 ;
        RECT 137.415 138.025 137.705 138.255 ;
        RECT 137.950 138.210 138.090 138.410 ;
        RECT 138.295 138.410 142.295 138.550 ;
        RECT 138.295 138.365 138.585 138.410 ;
        RECT 139.485 138.365 139.775 138.410 ;
        RECT 142.005 138.365 142.295 138.410 ;
        RECT 138.695 138.210 138.985 138.255 ;
        RECT 137.950 138.070 138.985 138.210 ;
        RECT 138.695 138.025 138.985 138.070 ;
        RECT 137.490 137.870 137.630 138.025 ;
        RECT 131.510 137.730 137.630 137.870 ;
        RECT 122.680 137.670 123.000 137.685 ;
        RECT 136.110 137.590 136.250 137.730 ;
        RECT 70.240 137.530 70.560 137.590 ;
        RECT 73.015 137.530 73.305 137.575 ;
        RECT 77.600 137.530 77.920 137.590 ;
        RECT 70.240 137.390 77.920 137.530 ;
        RECT 70.240 137.330 70.560 137.390 ;
        RECT 73.015 137.345 73.305 137.390 ;
        RECT 77.600 137.330 77.920 137.390 ;
        RECT 88.180 137.330 88.500 137.590 ;
        RECT 90.480 137.330 90.800 137.590 ;
        RECT 90.940 137.530 91.260 137.590 ;
        RECT 92.335 137.530 92.625 137.575 ;
        RECT 90.940 137.390 92.625 137.530 ;
        RECT 90.940 137.330 91.260 137.390 ;
        RECT 92.335 137.345 92.625 137.390 ;
        RECT 94.620 137.330 94.940 137.590 ;
        RECT 104.740 137.330 105.060 137.590 ;
        RECT 136.020 137.330 136.340 137.590 ;
        RECT 17.270 136.710 146.990 137.190 ;
        RECT 21.495 136.510 21.785 136.555 ;
        RECT 30.220 136.510 30.540 136.570 ;
        RECT 21.495 136.370 30.540 136.510 ;
        RECT 21.495 136.325 21.785 136.370 ;
        RECT 30.220 136.310 30.540 136.370 ;
        RECT 32.520 136.310 32.840 136.570 ;
        RECT 73.460 136.510 73.780 136.570 ;
        RECT 99.695 136.510 99.985 136.555 ;
        RECT 102.440 136.510 102.760 136.570 ;
        RECT 73.460 136.370 76.910 136.510 ;
        RECT 73.460 136.310 73.780 136.370 ;
        RECT 16.420 136.170 16.740 136.230 ;
        RECT 66.575 136.170 66.865 136.215 ;
        RECT 70.560 136.170 70.850 136.215 ;
        RECT 16.420 136.030 20.790 136.170 ;
        RECT 16.420 135.970 16.740 136.030 ;
        RECT 20.650 135.875 20.790 136.030 ;
        RECT 66.575 136.030 70.850 136.170 ;
        RECT 66.575 135.985 66.865 136.030 ;
        RECT 70.560 135.985 70.850 136.030 ;
        RECT 26.080 135.875 26.400 135.890 ;
        RECT 20.115 135.645 20.405 135.875 ;
        RECT 20.575 135.645 20.865 135.875 ;
        RECT 26.050 135.645 26.400 135.875 ;
        RECT 20.190 135.150 20.330 135.645 ;
        RECT 26.080 135.630 26.400 135.645 ;
        RECT 32.060 135.630 32.380 135.890 ;
        RECT 65.180 135.630 65.500 135.890 ;
        RECT 66.115 135.830 66.405 135.875 ;
        RECT 67.020 135.830 67.340 135.890 ;
        RECT 66.115 135.690 67.340 135.830 ;
        RECT 66.115 135.645 66.405 135.690 ;
        RECT 67.020 135.630 67.340 135.690 ;
        RECT 67.495 135.645 67.785 135.875 ;
        RECT 21.020 135.490 21.340 135.550 ;
        RECT 24.700 135.490 25.020 135.550 ;
        RECT 21.020 135.350 25.020 135.490 ;
        RECT 21.020 135.290 21.340 135.350 ;
        RECT 24.700 135.290 25.020 135.350 ;
        RECT 25.595 135.490 25.885 135.535 ;
        RECT 26.785 135.490 27.075 135.535 ;
        RECT 29.305 135.490 29.595 135.535 ;
        RECT 67.570 135.490 67.710 135.645 ;
        RECT 68.400 135.630 68.720 135.890 ;
        RECT 69.335 135.830 69.625 135.875 ;
        RECT 69.780 135.830 70.100 135.890 ;
        RECT 76.770 135.875 76.910 136.370 ;
        RECT 99.695 136.370 102.760 136.510 ;
        RECT 99.695 136.325 99.985 136.370 ;
        RECT 102.440 136.310 102.760 136.370 ;
        RECT 112.560 136.510 112.880 136.570 ;
        RECT 113.955 136.510 114.245 136.555 ;
        RECT 112.560 136.370 114.245 136.510 ;
        RECT 112.560 136.310 112.880 136.370 ;
        RECT 113.955 136.325 114.245 136.370 ;
        RECT 116.700 136.310 117.020 136.570 ;
        RECT 122.220 136.510 122.540 136.570 ;
        RECT 128.675 136.510 128.965 136.555 ;
        RECT 134.640 136.510 134.960 136.570 ;
        RECT 122.220 136.370 128.965 136.510 ;
        RECT 122.220 136.310 122.540 136.370 ;
        RECT 128.675 136.325 128.965 136.370 ;
        RECT 129.670 136.370 134.960 136.510 ;
        RECT 88.180 136.215 88.500 136.230 ;
        RECT 88.150 136.170 88.500 136.215 ;
        RECT 78.970 136.030 82.890 136.170 ;
        RECT 87.985 136.030 88.500 136.170 ;
        RECT 69.335 135.690 70.100 135.830 ;
        RECT 69.335 135.645 69.625 135.690 ;
        RECT 69.780 135.630 70.100 135.690 ;
        RECT 76.695 135.830 76.985 135.875 ;
        RECT 77.140 135.830 77.460 135.890 ;
        RECT 76.695 135.690 77.460 135.830 ;
        RECT 76.695 135.645 76.985 135.690 ;
        RECT 77.140 135.630 77.460 135.690 ;
        RECT 77.600 135.875 77.920 135.890 ;
        RECT 77.600 135.830 77.955 135.875 ;
        RECT 78.970 135.830 79.110 136.030 ;
        RECT 77.600 135.690 79.110 135.830 ;
        RECT 77.600 135.645 77.955 135.690 ;
        RECT 79.455 135.645 79.745 135.875 ;
        RECT 81.295 135.830 81.585 135.875 ;
        RECT 82.200 135.830 82.520 135.890 ;
        RECT 82.750 135.875 82.890 136.030 ;
        RECT 88.150 135.985 88.500 136.030 ;
        RECT 88.180 135.970 88.500 135.985 ;
        RECT 104.740 136.170 105.060 136.230 ;
        RECT 108.420 136.215 108.740 136.230 ;
        RECT 105.260 136.170 105.550 136.215 ;
        RECT 108.390 136.170 108.740 136.215 ;
        RECT 104.740 136.030 105.550 136.170 ;
        RECT 108.225 136.030 108.740 136.170 ;
        RECT 104.740 135.970 105.060 136.030 ;
        RECT 105.260 135.985 105.550 136.030 ;
        RECT 108.390 135.985 108.740 136.030 ;
        RECT 108.420 135.970 108.740 135.985 ;
        RECT 111.640 135.970 111.960 136.230 ;
        RECT 121.300 136.170 121.620 136.230 ;
        RECT 121.300 136.030 123.830 136.170 ;
        RECT 121.300 135.970 121.620 136.030 ;
        RECT 81.295 135.690 82.520 135.830 ;
        RECT 81.295 135.645 81.585 135.690 ;
        RECT 77.600 135.630 77.920 135.645 ;
        RECT 25.595 135.350 29.595 135.490 ;
        RECT 25.595 135.305 25.885 135.350 ;
        RECT 26.785 135.305 27.075 135.350 ;
        RECT 29.305 135.305 29.595 135.350 ;
        RECT 66.190 135.350 67.710 135.490 ;
        RECT 70.215 135.490 70.505 135.535 ;
        RECT 71.405 135.490 71.695 135.535 ;
        RECT 73.925 135.490 74.215 135.535 ;
        RECT 70.215 135.350 74.215 135.490 ;
        RECT 25.200 135.150 25.490 135.195 ;
        RECT 27.300 135.150 27.590 135.195 ;
        RECT 28.870 135.150 29.160 135.195 ;
        RECT 20.190 135.010 24.930 135.150 ;
        RECT 15.960 134.810 16.280 134.870 ;
        RECT 19.195 134.810 19.485 134.855 ;
        RECT 15.960 134.670 19.485 134.810 ;
        RECT 24.790 134.810 24.930 135.010 ;
        RECT 25.200 135.010 29.160 135.150 ;
        RECT 25.200 134.965 25.490 135.010 ;
        RECT 27.300 134.965 27.590 135.010 ;
        RECT 28.870 134.965 29.160 135.010 ;
        RECT 66.190 134.870 66.330 135.350 ;
        RECT 70.215 135.305 70.505 135.350 ;
        RECT 71.405 135.305 71.695 135.350 ;
        RECT 73.925 135.305 74.215 135.350 ;
        RECT 79.530 135.490 79.670 135.645 ;
        RECT 82.200 135.630 82.520 135.690 ;
        RECT 82.675 135.645 82.965 135.875 ;
        RECT 84.515 135.830 84.805 135.875 ;
        RECT 85.880 135.830 86.200 135.890 ;
        RECT 84.515 135.690 86.200 135.830 ;
        RECT 84.515 135.645 84.805 135.690 ;
        RECT 80.360 135.490 80.680 135.550 ;
        RECT 84.590 135.490 84.730 135.645 ;
        RECT 85.880 135.630 86.200 135.690 ;
        RECT 86.815 135.830 87.105 135.875 ;
        RECT 87.260 135.830 87.580 135.890 ;
        RECT 86.815 135.690 87.580 135.830 ;
        RECT 86.815 135.645 87.105 135.690 ;
        RECT 87.260 135.630 87.580 135.690 ;
        RECT 106.595 135.830 106.885 135.875 ;
        RECT 107.055 135.830 107.345 135.875 ;
        RECT 111.730 135.830 111.870 135.970 ;
        RECT 106.595 135.690 111.870 135.830 ;
        RECT 106.595 135.645 106.885 135.690 ;
        RECT 107.055 135.645 107.345 135.690 ;
        RECT 117.620 135.630 117.940 135.890 ;
        RECT 118.540 135.630 118.860 135.890 ;
        RECT 123.690 135.875 123.830 136.030 ;
        RECT 123.615 135.645 123.905 135.875 ;
        RECT 127.280 135.630 127.600 135.890 ;
        RECT 129.670 135.875 129.810 136.370 ;
        RECT 134.640 136.310 134.960 136.370 ;
        RECT 144.760 136.310 145.080 136.570 ;
        RECT 133.275 136.170 133.565 136.215 ;
        RECT 130.130 136.030 140.850 136.170 ;
        RECT 130.130 135.875 130.270 136.030 ;
        RECT 133.275 135.985 133.565 136.030 ;
        RECT 129.595 135.645 129.885 135.875 ;
        RECT 130.055 135.645 130.345 135.875 ;
        RECT 130.975 135.645 131.265 135.875 ;
        RECT 79.530 135.350 80.680 135.490 ;
        RECT 69.820 135.150 70.110 135.195 ;
        RECT 71.920 135.150 72.210 135.195 ;
        RECT 73.490 135.150 73.780 135.195 ;
        RECT 77.155 135.150 77.445 135.195 ;
        RECT 69.820 135.010 73.780 135.150 ;
        RECT 69.820 134.965 70.110 135.010 ;
        RECT 71.920 134.965 72.210 135.010 ;
        RECT 73.490 134.965 73.780 135.010 ;
        RECT 75.390 135.010 77.445 135.150 ;
        RECT 31.600 134.810 31.920 134.870 ;
        RECT 24.790 134.670 31.920 134.810 ;
        RECT 15.960 134.610 16.280 134.670 ;
        RECT 19.195 134.625 19.485 134.670 ;
        RECT 31.600 134.610 31.920 134.670 ;
        RECT 66.100 134.610 66.420 134.870 ;
        RECT 67.020 134.810 67.340 134.870 ;
        RECT 75.390 134.810 75.530 135.010 ;
        RECT 77.155 134.965 77.445 135.010 ;
        RECT 67.020 134.670 75.530 134.810 ;
        RECT 76.220 134.810 76.540 134.870 ;
        RECT 79.530 134.810 79.670 135.350 ;
        RECT 80.360 135.290 80.680 135.350 ;
        RECT 81.370 135.350 84.730 135.490 ;
        RECT 87.695 135.490 87.985 135.535 ;
        RECT 88.885 135.490 89.175 135.535 ;
        RECT 91.405 135.490 91.695 135.535 ;
        RECT 87.695 135.350 91.695 135.490 ;
        RECT 76.220 134.670 79.670 134.810 ;
        RECT 79.900 134.810 80.220 134.870 ;
        RECT 81.370 134.855 81.510 135.350 ;
        RECT 87.695 135.305 87.985 135.350 ;
        RECT 88.885 135.305 89.175 135.350 ;
        RECT 91.405 135.305 91.695 135.350 ;
        RECT 102.005 135.490 102.295 135.535 ;
        RECT 104.525 135.490 104.815 135.535 ;
        RECT 105.715 135.490 106.005 135.535 ;
        RECT 102.005 135.350 106.005 135.490 ;
        RECT 102.005 135.305 102.295 135.350 ;
        RECT 104.525 135.305 104.815 135.350 ;
        RECT 105.715 135.305 106.005 135.350 ;
        RECT 107.935 135.490 108.225 135.535 ;
        RECT 109.125 135.490 109.415 135.535 ;
        RECT 111.645 135.490 111.935 135.535 ;
        RECT 107.935 135.350 111.935 135.490 ;
        RECT 107.935 135.305 108.225 135.350 ;
        RECT 109.125 135.305 109.415 135.350 ;
        RECT 111.645 135.305 111.935 135.350 ;
        RECT 119.015 135.490 119.305 135.535 ;
        RECT 120.855 135.490 121.145 135.535 ;
        RECT 129.670 135.490 129.810 135.645 ;
        RECT 119.015 135.350 121.145 135.490 ;
        RECT 119.015 135.305 119.305 135.350 ;
        RECT 120.855 135.305 121.145 135.350 ;
        RECT 122.310 135.350 129.810 135.490 ;
        RECT 81.740 135.150 82.060 135.210 ;
        RECT 87.300 135.150 87.590 135.195 ;
        RECT 89.400 135.150 89.690 135.195 ;
        RECT 90.970 135.150 91.260 135.195 ;
        RECT 81.740 135.010 83.350 135.150 ;
        RECT 81.740 134.950 82.060 135.010 ;
        RECT 81.295 134.810 81.585 134.855 ;
        RECT 79.900 134.670 81.585 134.810 ;
        RECT 67.020 134.610 67.340 134.670 ;
        RECT 76.220 134.610 76.540 134.670 ;
        RECT 79.900 134.610 80.220 134.670 ;
        RECT 81.295 134.625 81.585 134.670 ;
        RECT 82.200 134.610 82.520 134.870 ;
        RECT 83.210 134.855 83.350 135.010 ;
        RECT 87.300 135.010 91.260 135.150 ;
        RECT 87.300 134.965 87.590 135.010 ;
        RECT 89.400 134.965 89.690 135.010 ;
        RECT 90.970 134.965 91.260 135.010 ;
        RECT 102.440 135.150 102.730 135.195 ;
        RECT 104.010 135.150 104.300 135.195 ;
        RECT 106.110 135.150 106.400 135.195 ;
        RECT 102.440 135.010 106.400 135.150 ;
        RECT 102.440 134.965 102.730 135.010 ;
        RECT 104.010 134.965 104.300 135.010 ;
        RECT 106.110 134.965 106.400 135.010 ;
        RECT 107.540 135.150 107.830 135.195 ;
        RECT 109.640 135.150 109.930 135.195 ;
        RECT 111.210 135.150 111.500 135.195 ;
        RECT 107.540 135.010 111.500 135.150 ;
        RECT 107.540 134.965 107.830 135.010 ;
        RECT 109.640 134.965 109.930 135.010 ;
        RECT 111.210 134.965 111.500 135.010 ;
        RECT 115.320 135.150 115.640 135.210 ;
        RECT 122.310 135.150 122.450 135.350 ;
        RECT 131.050 135.150 131.190 135.645 ;
        RECT 131.420 135.630 131.740 135.890 ;
        RECT 133.720 135.630 134.040 135.890 ;
        RECT 136.480 135.830 136.800 135.890 ;
        RECT 137.315 135.830 137.605 135.875 ;
        RECT 136.480 135.690 137.605 135.830 ;
        RECT 140.710 135.830 140.850 136.030 ;
        RECT 143.855 135.830 144.145 135.875 ;
        RECT 144.300 135.830 144.620 135.890 ;
        RECT 140.710 135.690 143.150 135.830 ;
        RECT 136.480 135.630 136.800 135.690 ;
        RECT 137.315 135.645 137.605 135.690 ;
        RECT 132.815 135.305 133.105 135.535 ;
        RECT 115.320 135.010 122.450 135.150 ;
        RECT 122.770 135.010 131.190 135.150 ;
        RECT 132.890 135.150 133.030 135.305 ;
        RECT 136.020 135.290 136.340 135.550 ;
        RECT 136.915 135.490 137.205 135.535 ;
        RECT 138.105 135.490 138.395 135.535 ;
        RECT 140.625 135.490 140.915 135.535 ;
        RECT 136.915 135.350 140.915 135.490 ;
        RECT 136.915 135.305 137.205 135.350 ;
        RECT 138.105 135.305 138.395 135.350 ;
        RECT 140.625 135.305 140.915 135.350 ;
        RECT 143.010 135.195 143.150 135.690 ;
        RECT 143.855 135.690 144.620 135.830 ;
        RECT 143.855 135.645 144.145 135.690 ;
        RECT 144.300 135.630 144.620 135.690 ;
        RECT 136.520 135.150 136.810 135.195 ;
        RECT 138.620 135.150 138.910 135.195 ;
        RECT 140.190 135.150 140.480 135.195 ;
        RECT 132.890 135.010 136.250 135.150 ;
        RECT 115.320 134.950 115.640 135.010 ;
        RECT 83.135 134.625 83.425 134.855 ;
        RECT 84.500 134.810 84.820 134.870 ;
        RECT 85.435 134.810 85.725 134.855 ;
        RECT 84.500 134.670 85.725 134.810 ;
        RECT 84.500 134.610 84.820 134.670 ;
        RECT 85.435 134.625 85.725 134.670 ;
        RECT 90.480 134.810 90.800 134.870 ;
        RECT 93.700 134.810 94.020 134.870 ;
        RECT 90.480 134.670 94.020 134.810 ;
        RECT 90.480 134.610 90.800 134.670 ;
        RECT 93.700 134.610 94.020 134.670 ;
        RECT 119.460 134.810 119.780 134.870 ;
        RECT 122.770 134.810 122.910 135.010 ;
        RECT 119.460 134.670 122.910 134.810 ;
        RECT 123.140 134.810 123.460 134.870 ;
        RECT 124.535 134.810 124.825 134.855 ;
        RECT 123.140 134.670 124.825 134.810 ;
        RECT 119.460 134.610 119.780 134.670 ;
        RECT 123.140 134.610 123.460 134.670 ;
        RECT 124.535 134.625 124.825 134.670 ;
        RECT 135.560 134.610 135.880 134.870 ;
        RECT 136.110 134.810 136.250 135.010 ;
        RECT 136.520 135.010 140.480 135.150 ;
        RECT 136.520 134.965 136.810 135.010 ;
        RECT 138.620 134.965 138.910 135.010 ;
        RECT 140.190 134.965 140.480 135.010 ;
        RECT 142.935 135.150 143.225 135.195 ;
        RECT 143.840 135.150 144.160 135.210 ;
        RECT 142.935 135.010 144.160 135.150 ;
        RECT 142.935 134.965 143.225 135.010 ;
        RECT 143.840 134.950 144.160 135.010 ;
        RECT 140.620 134.810 140.940 134.870 ;
        RECT 136.110 134.670 140.940 134.810 ;
        RECT 140.620 134.610 140.940 134.670 ;
        RECT 17.270 133.990 146.990 134.470 ;
        RECT 26.080 133.790 26.400 133.850 ;
        RECT 27.015 133.790 27.305 133.835 ;
        RECT 26.080 133.650 27.305 133.790 ;
        RECT 26.080 133.590 26.400 133.650 ;
        RECT 27.015 133.605 27.305 133.650 ;
        RECT 65.180 133.790 65.500 133.850 ;
        RECT 68.400 133.790 68.720 133.850 ;
        RECT 69.795 133.790 70.085 133.835 ;
        RECT 76.220 133.790 76.540 133.850 ;
        RECT 65.180 133.650 68.170 133.790 ;
        RECT 65.180 133.590 65.500 133.650 ;
        RECT 19.680 133.450 19.970 133.495 ;
        RECT 21.780 133.450 22.070 133.495 ;
        RECT 23.350 133.450 23.640 133.495 ;
        RECT 19.680 133.310 23.640 133.450 ;
        RECT 19.680 133.265 19.970 133.310 ;
        RECT 21.780 133.265 22.070 133.310 ;
        RECT 23.350 133.265 23.640 133.310 ;
        RECT 28.395 133.450 28.685 133.495 ;
        RECT 31.140 133.450 31.460 133.510 ;
        RECT 28.395 133.310 31.460 133.450 ;
        RECT 28.395 133.265 28.685 133.310 ;
        RECT 31.140 133.250 31.460 133.310 ;
        RECT 62.460 133.450 62.750 133.495 ;
        RECT 64.560 133.450 64.850 133.495 ;
        RECT 66.130 133.450 66.420 133.495 ;
        RECT 62.460 133.310 66.420 133.450 ;
        RECT 62.460 133.265 62.750 133.310 ;
        RECT 64.560 133.265 64.850 133.310 ;
        RECT 66.130 133.265 66.420 133.310 ;
        RECT 20.075 133.110 20.365 133.155 ;
        RECT 21.265 133.110 21.555 133.155 ;
        RECT 23.785 133.110 24.075 133.155 ;
        RECT 20.075 132.970 24.075 133.110 ;
        RECT 20.075 132.925 20.365 132.970 ;
        RECT 21.265 132.925 21.555 132.970 ;
        RECT 23.785 132.925 24.075 132.970 ;
        RECT 28.855 133.110 29.145 133.155 ;
        RECT 33.455 133.110 33.745 133.155 ;
        RECT 28.855 132.970 33.745 133.110 ;
        RECT 28.855 132.925 29.145 132.970 ;
        RECT 33.455 132.925 33.745 132.970 ;
        RECT 62.855 133.110 63.145 133.155 ;
        RECT 64.045 133.110 64.335 133.155 ;
        RECT 66.565 133.110 66.855 133.155 ;
        RECT 62.855 132.970 66.855 133.110 ;
        RECT 68.030 133.110 68.170 133.650 ;
        RECT 68.400 133.650 70.085 133.790 ;
        RECT 68.400 133.590 68.720 133.650 ;
        RECT 69.795 133.605 70.085 133.650 ;
        RECT 71.710 133.650 76.540 133.790 ;
        RECT 71.710 133.155 71.850 133.650 ;
        RECT 76.220 133.590 76.540 133.650 ;
        RECT 77.140 133.790 77.460 133.850 ;
        RECT 79.455 133.790 79.745 133.835 ;
        RECT 79.900 133.790 80.220 133.850 ;
        RECT 113.480 133.790 113.800 133.850 ;
        RECT 114.875 133.790 115.165 133.835 ;
        RECT 115.320 133.790 115.640 133.850 ;
        RECT 77.140 133.650 80.220 133.790 ;
        RECT 77.140 133.590 77.460 133.650 ;
        RECT 79.455 133.605 79.745 133.650 ;
        RECT 79.900 133.590 80.220 133.650 ;
        RECT 101.610 133.650 112.790 133.790 ;
        RECT 73.040 133.450 73.330 133.495 ;
        RECT 75.140 133.450 75.430 133.495 ;
        RECT 76.710 133.450 77.000 133.495 ;
        RECT 73.040 133.310 77.000 133.450 ;
        RECT 73.040 133.265 73.330 133.310 ;
        RECT 75.140 133.265 75.430 133.310 ;
        RECT 76.710 133.265 77.000 133.310 ;
        RECT 88.220 133.450 88.510 133.495 ;
        RECT 90.320 133.450 90.610 133.495 ;
        RECT 91.890 133.450 92.180 133.495 ;
        RECT 88.220 133.310 92.180 133.450 ;
        RECT 88.220 133.265 88.510 133.310 ;
        RECT 90.320 133.265 90.610 133.310 ;
        RECT 91.890 133.265 92.180 133.310 ;
        RECT 71.635 133.110 71.925 133.155 ;
        RECT 68.030 132.970 71.925 133.110 ;
        RECT 62.855 132.925 63.145 132.970 ;
        RECT 64.045 132.925 64.335 132.970 ;
        RECT 66.565 132.925 66.855 132.970 ;
        RECT 71.635 132.925 71.925 132.970 ;
        RECT 72.080 133.110 72.400 133.170 ;
        RECT 72.555 133.110 72.845 133.155 ;
        RECT 72.080 132.970 72.845 133.110 ;
        RECT 72.080 132.910 72.400 132.970 ;
        RECT 72.555 132.925 72.845 132.970 ;
        RECT 73.435 133.110 73.725 133.155 ;
        RECT 74.625 133.110 74.915 133.155 ;
        RECT 77.145 133.110 77.435 133.155 ;
        RECT 73.435 132.970 77.435 133.110 ;
        RECT 73.435 132.925 73.725 132.970 ;
        RECT 74.625 132.925 74.915 132.970 ;
        RECT 77.145 132.925 77.435 132.970 ;
        RECT 84.500 132.910 84.820 133.170 ;
        RECT 87.720 132.910 88.040 133.170 ;
        RECT 88.615 133.110 88.905 133.155 ;
        RECT 89.805 133.110 90.095 133.155 ;
        RECT 92.325 133.110 92.615 133.155 ;
        RECT 88.615 132.970 92.615 133.110 ;
        RECT 88.615 132.925 88.905 132.970 ;
        RECT 89.805 132.925 90.095 132.970 ;
        RECT 92.325 132.925 92.615 132.970 ;
        RECT 93.700 133.110 94.020 133.170 ;
        RECT 100.155 133.110 100.445 133.155 ;
        RECT 101.610 133.110 101.750 133.650 ;
        RECT 107.055 133.265 107.345 133.495 ;
        RECT 108.460 133.450 108.750 133.495 ;
        RECT 110.560 133.450 110.850 133.495 ;
        RECT 112.130 133.450 112.420 133.495 ;
        RECT 108.460 133.310 112.420 133.450 ;
        RECT 112.650 133.450 112.790 133.650 ;
        RECT 113.480 133.650 115.640 133.790 ;
        RECT 113.480 133.590 113.800 133.650 ;
        RECT 114.875 133.605 115.165 133.650 ;
        RECT 115.320 133.590 115.640 133.650 ;
        RECT 120.855 133.790 121.145 133.835 ;
        RECT 122.680 133.790 123.000 133.850 ;
        RECT 120.855 133.650 123.000 133.790 ;
        RECT 120.855 133.605 121.145 133.650 ;
        RECT 122.680 133.590 123.000 133.650 ;
        RECT 136.035 133.790 136.325 133.835 ;
        RECT 136.480 133.790 136.800 133.850 ;
        RECT 136.035 133.650 136.800 133.790 ;
        RECT 136.035 133.605 136.325 133.650 ;
        RECT 136.480 133.590 136.800 133.650 ;
        RECT 144.760 133.590 145.080 133.850 ;
        RECT 128.200 133.450 128.520 133.510 ;
        RECT 130.960 133.450 131.280 133.510 ;
        RECT 112.650 133.310 131.280 133.450 ;
        RECT 108.460 133.265 108.750 133.310 ;
        RECT 110.560 133.265 110.850 133.310 ;
        RECT 112.130 133.265 112.420 133.310 ;
        RECT 93.700 132.970 101.750 133.110 ;
        RECT 103.360 133.110 103.680 133.170 ;
        RECT 103.835 133.110 104.125 133.155 ;
        RECT 103.360 132.970 104.125 133.110 ;
        RECT 93.700 132.910 94.020 132.970 ;
        RECT 100.155 132.925 100.445 132.970 ;
        RECT 103.360 132.910 103.680 132.970 ;
        RECT 103.835 132.925 104.125 132.970 ;
        RECT 104.280 133.110 104.600 133.170 ;
        RECT 104.755 133.110 105.045 133.155 ;
        RECT 104.280 132.970 105.045 133.110 ;
        RECT 104.280 132.910 104.600 132.970 ;
        RECT 104.755 132.925 105.045 132.970 ;
        RECT 19.195 132.770 19.485 132.815 ;
        RECT 19.640 132.770 19.960 132.830 ;
        RECT 19.195 132.630 19.960 132.770 ;
        RECT 19.195 132.585 19.485 132.630 ;
        RECT 19.640 132.570 19.960 132.630 ;
        RECT 27.935 132.585 28.225 132.815 ;
        RECT 29.315 132.770 29.605 132.815 ;
        RECT 30.695 132.770 30.985 132.815 ;
        RECT 29.315 132.630 30.985 132.770 ;
        RECT 29.315 132.585 29.605 132.630 ;
        RECT 30.695 132.585 30.985 132.630 ;
        RECT 20.530 132.430 20.820 132.475 ;
        RECT 21.940 132.430 22.260 132.490 ;
        RECT 20.530 132.290 22.260 132.430 ;
        RECT 20.530 132.245 20.820 132.290 ;
        RECT 21.940 132.230 22.260 132.290 ;
        RECT 26.080 131.890 26.400 132.150 ;
        RECT 28.010 132.090 28.150 132.585 ;
        RECT 31.600 132.570 31.920 132.830 ;
        RECT 33.915 132.770 34.205 132.815 ;
        RECT 33.915 132.630 34.315 132.770 ;
        RECT 33.915 132.585 34.205 132.630 ;
        RECT 32.520 132.430 32.840 132.490 ;
        RECT 33.990 132.430 34.130 132.585 ;
        RECT 61.960 132.570 62.280 132.830 ;
        RECT 67.020 132.770 67.340 132.830 ;
        RECT 73.920 132.815 74.240 132.830 ;
        RECT 70.715 132.770 71.005 132.815 ;
        RECT 67.020 132.630 71.005 132.770 ;
        RECT 67.020 132.570 67.340 132.630 ;
        RECT 70.715 132.585 71.005 132.630 ;
        RECT 73.890 132.585 74.240 132.815 ;
        RECT 85.435 132.770 85.725 132.815 ;
        RECT 86.340 132.770 86.660 132.830 ;
        RECT 85.435 132.630 86.660 132.770 ;
        RECT 85.435 132.585 85.725 132.630 ;
        RECT 73.920 132.570 74.240 132.585 ;
        RECT 86.340 132.570 86.660 132.630 ;
        RECT 89.070 132.770 89.360 132.815 ;
        RECT 90.940 132.770 91.260 132.830 ;
        RECT 89.070 132.630 91.260 132.770 ;
        RECT 89.070 132.585 89.360 132.630 ;
        RECT 90.940 132.570 91.260 132.630 ;
        RECT 98.760 132.570 99.080 132.830 ;
        RECT 107.130 132.770 107.270 133.265 ;
        RECT 128.200 133.250 128.520 133.310 ;
        RECT 130.960 133.250 131.280 133.310 ;
        RECT 135.560 133.250 135.880 133.510 ;
        RECT 108.855 133.110 109.145 133.155 ;
        RECT 110.045 133.110 110.335 133.155 ;
        RECT 112.565 133.110 112.855 133.155 ;
        RECT 108.855 132.970 112.855 133.110 ;
        RECT 108.855 132.925 109.145 132.970 ;
        RECT 110.045 132.925 110.335 132.970 ;
        RECT 112.565 132.925 112.855 132.970 ;
        RECT 118.540 133.110 118.860 133.170 ;
        RECT 122.695 133.110 122.985 133.155 ;
        RECT 118.540 132.970 122.985 133.110 ;
        RECT 118.540 132.910 118.860 132.970 ;
        RECT 122.695 132.925 122.985 132.970 ;
        RECT 123.140 132.910 123.460 133.170 ;
        RECT 107.975 132.770 108.265 132.815 ;
        RECT 111.640 132.770 111.960 132.830 ;
        RECT 107.130 132.630 107.730 132.770 ;
        RECT 35.740 132.430 36.060 132.490 ;
        RECT 32.520 132.290 36.060 132.430 ;
        RECT 32.520 132.230 32.840 132.290 ;
        RECT 35.740 132.230 36.060 132.290 ;
        RECT 63.310 132.430 63.600 132.475 ;
        RECT 64.720 132.430 65.040 132.490 ;
        RECT 63.310 132.290 65.040 132.430 ;
        RECT 63.310 132.245 63.600 132.290 ;
        RECT 64.720 132.230 65.040 132.290 ;
        RECT 84.975 132.430 85.265 132.475 ;
        RECT 95.555 132.430 95.845 132.475 ;
        RECT 84.975 132.290 95.845 132.430 ;
        RECT 84.975 132.245 85.265 132.290 ;
        RECT 95.555 132.245 95.845 132.290 ;
        RECT 102.915 132.430 103.205 132.475 ;
        RECT 105.215 132.430 105.505 132.475 ;
        RECT 102.915 132.290 105.505 132.430 ;
        RECT 107.590 132.430 107.730 132.630 ;
        RECT 107.975 132.630 111.960 132.770 ;
        RECT 107.975 132.585 108.265 132.630 ;
        RECT 111.640 132.570 111.960 132.630 ;
        RECT 121.775 132.770 122.065 132.815 ;
        RECT 128.660 132.770 128.980 132.830 ;
        RECT 121.775 132.630 128.980 132.770 ;
        RECT 121.775 132.585 122.065 132.630 ;
        RECT 128.660 132.570 128.980 132.630 ;
        RECT 142.000 132.570 142.320 132.830 ;
        RECT 143.840 132.570 144.160 132.830 ;
        RECT 109.200 132.430 109.490 132.475 ;
        RECT 107.590 132.290 109.490 132.430 ;
        RECT 102.915 132.245 103.205 132.290 ;
        RECT 105.215 132.245 105.505 132.290 ;
        RECT 109.200 132.245 109.490 132.290 ;
        RECT 130.500 132.430 130.820 132.490 ;
        RECT 133.735 132.430 134.025 132.475 ;
        RECT 130.500 132.290 134.025 132.430 ;
        RECT 130.500 132.230 130.820 132.290 ;
        RECT 133.735 132.245 134.025 132.290 ;
        RECT 30.220 132.090 30.540 132.150 ;
        RECT 34.820 132.090 35.140 132.150 ;
        RECT 28.010 131.950 35.140 132.090 ;
        RECT 30.220 131.890 30.540 131.950 ;
        RECT 34.820 131.890 35.140 131.950 ;
        RECT 68.400 132.090 68.720 132.150 ;
        RECT 68.875 132.090 69.165 132.135 ;
        RECT 68.400 131.950 69.165 132.090 ;
        RECT 68.400 131.890 68.720 131.950 ;
        RECT 68.875 131.905 69.165 131.950 ;
        RECT 86.800 132.090 87.120 132.150 ;
        RECT 87.275 132.090 87.565 132.135 ;
        RECT 86.800 131.950 87.565 132.090 ;
        RECT 86.800 131.890 87.120 131.950 ;
        RECT 87.275 131.905 87.565 131.950 ;
        RECT 94.620 132.090 94.940 132.150 ;
        RECT 98.300 132.090 98.620 132.150 ;
        RECT 136.480 132.090 136.800 132.150 ;
        RECT 139.240 132.090 139.560 132.150 ;
        RECT 94.620 131.950 139.560 132.090 ;
        RECT 94.620 131.890 94.940 131.950 ;
        RECT 98.300 131.890 98.620 131.950 ;
        RECT 136.480 131.890 136.800 131.950 ;
        RECT 139.240 131.890 139.560 131.950 ;
        RECT 142.920 131.890 143.240 132.150 ;
        RECT 17.270 131.270 146.990 131.750 ;
        RECT 21.940 130.870 22.260 131.130 ;
        RECT 72.080 131.070 72.400 131.130 ;
        RECT 103.360 131.070 103.680 131.130 ;
        RECT 107.040 131.070 107.360 131.130 ;
        RECT 72.080 130.930 84.270 131.070 ;
        RECT 72.080 130.870 72.400 130.930 ;
        RECT 23.795 130.730 24.085 130.775 ;
        RECT 26.080 130.730 26.400 130.790 ;
        RECT 20.190 130.590 26.400 130.730 ;
        RECT 20.190 130.435 20.330 130.590 ;
        RECT 23.795 130.545 24.085 130.590 ;
        RECT 26.080 130.530 26.400 130.590 ;
        RECT 63.815 130.730 64.105 130.775 ;
        RECT 66.560 130.730 66.880 130.790 ;
        RECT 63.815 130.590 66.880 130.730 ;
        RECT 63.815 130.545 64.105 130.590 ;
        RECT 66.560 130.530 66.880 130.590 ;
        RECT 20.115 130.205 20.405 130.435 ;
        RECT 24.240 130.190 24.560 130.450 ;
        RECT 61.960 130.390 62.280 130.450 ;
        RECT 70.700 130.435 71.020 130.450 ;
        RECT 62.895 130.390 63.185 130.435 ;
        RECT 61.960 130.250 63.185 130.390 ;
        RECT 61.960 130.190 62.280 130.250 ;
        RECT 62.895 130.205 63.185 130.250 ;
        RECT 70.670 130.205 71.020 130.435 ;
        RECT 25.175 130.050 25.465 130.095 ;
        RECT 32.520 130.050 32.840 130.110 ;
        RECT 25.175 129.910 32.840 130.050 ;
        RECT 62.970 130.050 63.110 130.205 ;
        RECT 70.700 130.190 71.020 130.205 ;
        RECT 82.660 130.435 82.980 130.450 ;
        RECT 84.130 130.435 84.270 130.930 ;
        RECT 103.360 130.930 107.360 131.070 ;
        RECT 103.360 130.870 103.680 130.930 ;
        RECT 107.040 130.870 107.360 130.930 ;
        RECT 129.120 131.070 129.440 131.130 ;
        RECT 131.880 131.070 132.200 131.130 ;
        RECT 137.400 131.070 137.720 131.130 ;
        RECT 129.120 130.930 137.720 131.070 ;
        RECT 129.120 130.870 129.440 130.930 ;
        RECT 131.880 130.870 132.200 130.930 ;
        RECT 137.400 130.870 137.720 130.930 ;
        RECT 87.720 130.730 88.040 130.790 ;
        RECT 85.510 130.590 88.040 130.730 ;
        RECT 85.510 130.435 85.650 130.590 ;
        RECT 87.720 130.530 88.040 130.590 ;
        RECT 104.280 130.730 104.600 130.790 ;
        RECT 104.280 130.590 108.650 130.730 ;
        RECT 104.280 130.530 104.600 130.590 ;
        RECT 86.800 130.435 87.120 130.450 ;
        RECT 82.660 130.205 83.010 130.435 ;
        RECT 84.055 130.390 84.345 130.435 ;
        RECT 85.435 130.390 85.725 130.435 ;
        RECT 86.770 130.390 87.120 130.435 ;
        RECT 84.055 130.250 85.725 130.390 ;
        RECT 86.605 130.250 87.120 130.390 ;
        RECT 84.055 130.205 84.345 130.250 ;
        RECT 85.435 130.205 85.725 130.250 ;
        RECT 86.770 130.205 87.120 130.250 ;
        RECT 82.660 130.190 82.980 130.205 ;
        RECT 86.800 130.190 87.120 130.205 ;
        RECT 106.580 130.190 106.900 130.450 ;
        RECT 107.040 130.190 107.360 130.450 ;
        RECT 107.960 130.190 108.280 130.450 ;
        RECT 108.510 130.435 108.650 130.590 ;
        RECT 109.340 130.530 109.660 130.790 ;
        RECT 142.000 130.730 142.320 130.790 ;
        RECT 121.390 130.590 142.320 130.730 ;
        RECT 108.435 130.205 108.725 130.435 ;
        RECT 111.640 130.190 111.960 130.450 ;
        RECT 112.100 130.390 112.420 130.450 ;
        RECT 112.935 130.390 113.225 130.435 ;
        RECT 112.100 130.250 113.225 130.390 ;
        RECT 112.100 130.190 112.420 130.250 ;
        RECT 112.935 130.205 113.225 130.250 ;
        RECT 66.560 130.050 66.880 130.110 ;
        RECT 67.955 130.050 68.245 130.095 ;
        RECT 69.335 130.050 69.625 130.095 ;
        RECT 62.970 129.910 69.625 130.050 ;
        RECT 25.175 129.865 25.465 129.910 ;
        RECT 32.520 129.850 32.840 129.910 ;
        RECT 66.560 129.850 66.880 129.910 ;
        RECT 67.955 129.865 68.245 129.910 ;
        RECT 69.335 129.865 69.625 129.910 ;
        RECT 70.215 130.050 70.505 130.095 ;
        RECT 71.405 130.050 71.695 130.095 ;
        RECT 73.925 130.050 74.215 130.095 ;
        RECT 70.215 129.910 74.215 130.050 ;
        RECT 70.215 129.865 70.505 129.910 ;
        RECT 71.405 129.865 71.695 129.910 ;
        RECT 73.925 129.865 74.215 129.910 ;
        RECT 79.465 130.050 79.755 130.095 ;
        RECT 81.985 130.050 82.275 130.095 ;
        RECT 83.175 130.050 83.465 130.095 ;
        RECT 79.465 129.910 83.465 130.050 ;
        RECT 79.465 129.865 79.755 129.910 ;
        RECT 81.985 129.865 82.275 129.910 ;
        RECT 83.175 129.865 83.465 129.910 ;
        RECT 86.315 130.050 86.605 130.095 ;
        RECT 87.505 130.050 87.795 130.095 ;
        RECT 90.025 130.050 90.315 130.095 ;
        RECT 98.315 130.050 98.605 130.095 ;
        RECT 98.760 130.050 99.080 130.110 ;
        RECT 111.180 130.050 111.500 130.110 ;
        RECT 86.315 129.910 90.315 130.050 ;
        RECT 86.315 129.865 86.605 129.910 ;
        RECT 87.505 129.865 87.795 129.910 ;
        RECT 90.025 129.865 90.315 129.910 ;
        RECT 92.410 129.910 111.500 130.050 ;
        RECT 15.960 129.710 16.280 129.770 ;
        RECT 92.410 129.755 92.550 129.910 ;
        RECT 98.315 129.865 98.605 129.910 ;
        RECT 98.760 129.850 99.080 129.910 ;
        RECT 111.180 129.850 111.500 129.910 ;
        RECT 112.535 130.050 112.825 130.095 ;
        RECT 113.725 130.050 114.015 130.095 ;
        RECT 116.245 130.050 116.535 130.095 ;
        RECT 112.535 129.910 116.535 130.050 ;
        RECT 112.535 129.865 112.825 129.910 ;
        RECT 113.725 129.865 114.015 129.910 ;
        RECT 116.245 129.865 116.535 129.910 ;
        RECT 19.195 129.710 19.485 129.755 ;
        RECT 15.960 129.570 19.485 129.710 ;
        RECT 15.960 129.510 16.280 129.570 ;
        RECT 19.195 129.525 19.485 129.570 ;
        RECT 69.820 129.710 70.110 129.755 ;
        RECT 71.920 129.710 72.210 129.755 ;
        RECT 73.490 129.710 73.780 129.755 ;
        RECT 69.820 129.570 73.780 129.710 ;
        RECT 69.820 129.525 70.110 129.570 ;
        RECT 71.920 129.525 72.210 129.570 ;
        RECT 73.490 129.525 73.780 129.570 ;
        RECT 79.900 129.710 80.190 129.755 ;
        RECT 81.470 129.710 81.760 129.755 ;
        RECT 83.570 129.710 83.860 129.755 ;
        RECT 79.900 129.570 83.860 129.710 ;
        RECT 79.900 129.525 80.190 129.570 ;
        RECT 81.470 129.525 81.760 129.570 ;
        RECT 83.570 129.525 83.860 129.570 ;
        RECT 85.920 129.710 86.210 129.755 ;
        RECT 88.020 129.710 88.310 129.755 ;
        RECT 89.590 129.710 89.880 129.755 ;
        RECT 85.920 129.570 89.880 129.710 ;
        RECT 85.920 129.525 86.210 129.570 ;
        RECT 88.020 129.525 88.310 129.570 ;
        RECT 89.590 129.525 89.880 129.570 ;
        RECT 92.335 129.525 92.625 129.755 ;
        RECT 112.140 129.710 112.430 129.755 ;
        RECT 114.240 129.710 114.530 129.755 ;
        RECT 115.810 129.710 116.100 129.755 ;
        RECT 112.140 129.570 116.100 129.710 ;
        RECT 112.140 129.525 112.430 129.570 ;
        RECT 114.240 129.525 114.530 129.570 ;
        RECT 115.810 129.525 116.100 129.570 ;
        RECT 118.555 129.710 118.845 129.755 ;
        RECT 121.390 129.710 121.530 130.590 ;
        RECT 142.000 130.530 142.320 130.590 ;
        RECT 129.595 130.390 129.885 130.435 ;
        RECT 130.040 130.390 130.360 130.450 ;
        RECT 134.180 130.390 134.500 130.450 ;
        RECT 129.595 130.250 134.500 130.390 ;
        RECT 129.595 130.205 129.885 130.250 ;
        RECT 130.040 130.190 130.360 130.250 ;
        RECT 134.180 130.190 134.500 130.250 ;
        RECT 123.155 130.050 123.445 130.095 ;
        RECT 126.360 130.050 126.680 130.110 ;
        RECT 130.500 130.050 130.820 130.110 ;
        RECT 123.155 129.910 130.820 130.050 ;
        RECT 123.155 129.865 123.445 129.910 ;
        RECT 126.360 129.850 126.680 129.910 ;
        RECT 130.500 129.850 130.820 129.910 ;
        RECT 137.875 129.865 138.165 130.095 ;
        RECT 138.320 130.050 138.640 130.110 ;
        RECT 138.795 130.050 139.085 130.095 ;
        RECT 140.620 130.050 140.940 130.110 ;
        RECT 138.320 129.910 140.940 130.050 ;
        RECT 118.555 129.570 121.530 129.710 ;
        RECT 121.775 129.710 122.065 129.755 ;
        RECT 126.820 129.710 127.140 129.770 ;
        RECT 121.775 129.570 127.140 129.710 ;
        RECT 118.555 129.525 118.845 129.570 ;
        RECT 121.775 129.525 122.065 129.570 ;
        RECT 73.000 129.370 73.320 129.430 ;
        RECT 76.235 129.370 76.525 129.415 ;
        RECT 73.000 129.230 76.525 129.370 ;
        RECT 73.000 129.170 73.320 129.230 ;
        RECT 76.235 129.185 76.525 129.230 ;
        RECT 77.140 129.170 77.460 129.430 ;
        RECT 101.075 129.370 101.365 129.415 ;
        RECT 102.440 129.370 102.760 129.430 ;
        RECT 101.075 129.230 102.760 129.370 ;
        RECT 101.075 129.185 101.365 129.230 ;
        RECT 102.440 129.170 102.760 129.230 ;
        RECT 107.960 129.370 108.280 129.430 ;
        RECT 118.630 129.370 118.770 129.525 ;
        RECT 126.820 129.510 127.140 129.570 ;
        RECT 131.435 129.710 131.725 129.755 ;
        RECT 133.720 129.710 134.040 129.770 ;
        RECT 131.435 129.570 134.040 129.710 ;
        RECT 131.435 129.525 131.725 129.570 ;
        RECT 133.720 129.510 134.040 129.570 ;
        RECT 135.100 129.710 135.420 129.770 ;
        RECT 137.950 129.710 138.090 129.865 ;
        RECT 138.320 129.850 138.640 129.910 ;
        RECT 138.795 129.865 139.085 129.910 ;
        RECT 140.620 129.850 140.940 129.910 ;
        RECT 135.100 129.570 138.090 129.710 ;
        RECT 135.100 129.510 135.420 129.570 ;
        RECT 107.960 129.230 118.770 129.370 ;
        RECT 120.855 129.370 121.145 129.415 ;
        RECT 121.300 129.370 121.620 129.430 ;
        RECT 120.855 129.230 121.620 129.370 ;
        RECT 107.960 129.170 108.280 129.230 ;
        RECT 120.855 129.185 121.145 129.230 ;
        RECT 121.300 129.170 121.620 129.230 ;
        RECT 131.880 129.170 132.200 129.430 ;
        RECT 132.340 129.370 132.660 129.430 ;
        RECT 135.575 129.370 135.865 129.415 ;
        RECT 132.340 129.230 135.865 129.370 ;
        RECT 132.340 129.170 132.660 129.230 ;
        RECT 135.575 129.185 135.865 129.230 ;
        RECT 17.270 128.550 146.990 129.030 ;
        RECT 64.720 128.150 65.040 128.410 ;
        RECT 70.700 128.350 71.020 128.410 ;
        RECT 71.635 128.350 71.925 128.395 ;
        RECT 70.700 128.210 71.925 128.350 ;
        RECT 70.700 128.150 71.020 128.210 ;
        RECT 71.635 128.165 71.925 128.210 ;
        RECT 82.215 128.350 82.505 128.395 ;
        RECT 82.660 128.350 82.980 128.410 ;
        RECT 82.215 128.210 82.980 128.350 ;
        RECT 82.215 128.165 82.505 128.210 ;
        RECT 82.660 128.150 82.980 128.210 ;
        RECT 111.195 128.350 111.485 128.395 ;
        RECT 112.100 128.350 112.420 128.410 ;
        RECT 111.195 128.210 112.420 128.350 ;
        RECT 111.195 128.165 111.485 128.210 ;
        RECT 112.100 128.150 112.420 128.210 ;
        RECT 117.620 128.150 117.940 128.410 ;
        RECT 128.660 128.350 128.980 128.410 ;
        RECT 133.735 128.350 134.025 128.395 ;
        RECT 128.660 128.210 134.025 128.350 ;
        RECT 128.660 128.150 128.980 128.210 ;
        RECT 133.735 128.165 134.025 128.210 ;
        RECT 15.960 128.010 16.280 128.070 ;
        RECT 19.195 128.010 19.485 128.055 ;
        RECT 101.520 128.010 101.840 128.070 ;
        RECT 15.400 127.870 19.485 128.010 ;
        RECT 15.960 127.810 16.280 127.870 ;
        RECT 19.195 127.825 19.485 127.870 ;
        RECT 91.030 127.870 101.840 128.010 ;
        RECT 66.100 127.670 66.420 127.730 ;
        RECT 67.495 127.670 67.785 127.715 ;
        RECT 20.190 127.530 25.620 127.670 ;
        RECT 20.190 127.375 20.330 127.530 ;
        RECT 25.480 127.390 25.620 127.530 ;
        RECT 66.100 127.530 67.785 127.670 ;
        RECT 66.100 127.470 66.420 127.530 ;
        RECT 67.495 127.485 67.785 127.530 ;
        RECT 72.540 127.670 72.860 127.730 ;
        RECT 74.395 127.670 74.685 127.715 ;
        RECT 72.540 127.530 74.685 127.670 ;
        RECT 72.540 127.470 72.860 127.530 ;
        RECT 74.395 127.485 74.685 127.530 ;
        RECT 82.200 127.670 82.520 127.730 ;
        RECT 84.975 127.670 85.265 127.715 ;
        RECT 91.030 127.670 91.170 127.870 ;
        RECT 101.520 127.810 101.840 127.870 ;
        RECT 110.735 128.010 111.025 128.055 ;
        RECT 111.655 128.010 111.945 128.055 ;
        RECT 110.735 127.870 111.945 128.010 ;
        RECT 110.735 127.825 111.025 127.870 ;
        RECT 111.655 127.825 111.945 127.870 ;
        RECT 121.340 128.010 121.630 128.055 ;
        RECT 123.440 128.010 123.730 128.055 ;
        RECT 125.010 128.010 125.300 128.055 ;
        RECT 121.340 127.870 125.300 128.010 ;
        RECT 121.340 127.825 121.630 127.870 ;
        RECT 123.440 127.825 123.730 127.870 ;
        RECT 125.010 127.825 125.300 127.870 ;
        RECT 132.340 127.810 132.660 128.070 ;
        RECT 136.020 128.010 136.340 128.070 ;
        RECT 137.900 128.010 138.190 128.055 ;
        RECT 140.000 128.010 140.290 128.055 ;
        RECT 141.570 128.010 141.860 128.055 ;
        RECT 136.020 127.870 137.630 128.010 ;
        RECT 136.020 127.810 136.340 127.870 ;
        RECT 82.200 127.530 85.265 127.670 ;
        RECT 82.200 127.470 82.520 127.530 ;
        RECT 84.975 127.485 85.265 127.530 ;
        RECT 89.190 127.530 91.170 127.670 ;
        RECT 99.695 127.670 99.985 127.715 ;
        RECT 103.360 127.670 103.680 127.730 ;
        RECT 99.695 127.530 103.680 127.670 ;
        RECT 20.115 127.145 20.405 127.375 ;
        RECT 21.940 127.130 22.260 127.390 ;
        RECT 25.480 127.330 25.940 127.390 ;
        RECT 27.015 127.330 27.305 127.375 ;
        RECT 25.480 127.190 27.305 127.330 ;
        RECT 25.620 127.130 25.940 127.190 ;
        RECT 27.015 127.145 27.305 127.190 ;
        RECT 67.035 127.330 67.325 127.375 ;
        RECT 68.860 127.330 69.180 127.390 ;
        RECT 73.935 127.330 74.225 127.375 ;
        RECT 67.035 127.190 74.225 127.330 ;
        RECT 67.035 127.145 67.325 127.190 ;
        RECT 68.860 127.130 69.180 127.190 ;
        RECT 73.935 127.145 74.225 127.190 ;
        RECT 84.055 127.330 84.345 127.375 ;
        RECT 86.340 127.330 86.660 127.390 ;
        RECT 89.190 127.330 89.330 127.530 ;
        RECT 99.695 127.485 99.985 127.530 ;
        RECT 103.360 127.470 103.680 127.530 ;
        RECT 107.960 127.670 108.280 127.730 ;
        RECT 113.955 127.670 114.245 127.715 ;
        RECT 107.960 127.530 114.245 127.670 ;
        RECT 107.960 127.470 108.280 127.530 ;
        RECT 113.955 127.485 114.245 127.530 ;
        RECT 114.860 127.470 115.180 127.730 ;
        RECT 115.320 127.670 115.640 127.730 ;
        RECT 121.735 127.670 122.025 127.715 ;
        RECT 122.925 127.670 123.215 127.715 ;
        RECT 125.445 127.670 125.735 127.715 ;
        RECT 115.320 127.530 118.770 127.670 ;
        RECT 115.320 127.470 115.640 127.530 ;
        RECT 84.055 127.190 86.660 127.330 ;
        RECT 84.055 127.145 84.345 127.190 ;
        RECT 86.340 127.130 86.660 127.190 ;
        RECT 88.270 127.190 89.330 127.330 ;
        RECT 89.560 127.330 89.880 127.390 ;
        RECT 96.015 127.330 96.305 127.375 ;
        RECT 118.080 127.330 118.400 127.390 ;
        RECT 118.630 127.375 118.770 127.530 ;
        RECT 121.735 127.530 125.735 127.670 ;
        RECT 121.735 127.485 122.025 127.530 ;
        RECT 122.925 127.485 123.215 127.530 ;
        RECT 125.445 127.485 125.735 127.530 ;
        RECT 130.500 127.470 130.820 127.730 ;
        RECT 136.940 127.670 137.260 127.730 ;
        RECT 137.490 127.715 137.630 127.870 ;
        RECT 137.900 127.870 141.860 128.010 ;
        RECT 137.900 127.825 138.190 127.870 ;
        RECT 140.000 127.825 140.290 127.870 ;
        RECT 141.570 127.825 141.860 127.870 ;
        RECT 136.110 127.530 137.260 127.670 ;
        RECT 89.560 127.190 118.400 127.330 ;
        RECT 26.095 126.990 26.385 127.035 ;
        RECT 26.540 126.990 26.860 127.050 ;
        RECT 26.095 126.850 26.860 126.990 ;
        RECT 26.095 126.805 26.385 126.850 ;
        RECT 26.540 126.790 26.860 126.850 ;
        RECT 73.000 126.990 73.320 127.050 ;
        RECT 73.475 126.990 73.765 127.035 ;
        RECT 73.000 126.850 73.765 126.990 ;
        RECT 73.000 126.790 73.320 126.850 ;
        RECT 73.475 126.805 73.765 126.850 ;
        RECT 77.140 126.990 77.460 127.050 ;
        RECT 84.515 126.990 84.805 127.035 ;
        RECT 88.270 126.990 88.410 127.190 ;
        RECT 89.560 127.130 89.880 127.190 ;
        RECT 96.015 127.145 96.305 127.190 ;
        RECT 118.080 127.130 118.400 127.190 ;
        RECT 118.555 127.145 118.845 127.375 ;
        RECT 119.015 127.145 119.305 127.375 ;
        RECT 77.140 126.850 88.410 126.990 ;
        RECT 88.640 126.990 88.960 127.050 ;
        RECT 91.875 126.990 92.165 127.035 ;
        RECT 88.640 126.850 92.165 126.990 ;
        RECT 77.140 126.790 77.460 126.850 ;
        RECT 84.515 126.805 84.805 126.850 ;
        RECT 86.430 126.710 86.570 126.850 ;
        RECT 88.640 126.790 88.960 126.850 ;
        RECT 91.875 126.805 92.165 126.850 ;
        RECT 98.300 126.790 98.620 127.050 ;
        RECT 98.775 126.990 99.065 127.035 ;
        RECT 101.980 126.990 102.300 127.050 ;
        RECT 98.775 126.850 102.300 126.990 ;
        RECT 98.775 126.805 99.065 126.850 ;
        RECT 101.980 126.790 102.300 126.850 ;
        RECT 102.440 126.790 102.760 127.050 ;
        RECT 108.880 126.790 109.200 127.050 ;
        RECT 113.480 126.790 113.800 127.050 ;
        RECT 21.020 126.450 21.340 126.710 ;
        RECT 27.935 126.650 28.225 126.695 ;
        RECT 31.600 126.650 31.920 126.710 ;
        RECT 27.935 126.510 31.920 126.650 ;
        RECT 27.935 126.465 28.225 126.510 ;
        RECT 31.600 126.450 31.920 126.510 ;
        RECT 66.575 126.650 66.865 126.695 ;
        RECT 68.400 126.650 68.720 126.710 ;
        RECT 71.620 126.650 71.940 126.710 ;
        RECT 66.575 126.510 71.940 126.650 ;
        RECT 66.575 126.465 66.865 126.510 ;
        RECT 68.400 126.450 68.720 126.510 ;
        RECT 71.620 126.450 71.940 126.510 ;
        RECT 86.340 126.450 86.660 126.710 ;
        RECT 96.460 126.450 96.780 126.710 ;
        RECT 99.220 126.650 99.540 126.710 ;
        RECT 100.615 126.650 100.905 126.695 ;
        RECT 99.220 126.510 100.905 126.650 ;
        RECT 99.220 126.450 99.540 126.510 ;
        RECT 100.615 126.465 100.905 126.510 ;
        RECT 102.915 126.650 103.205 126.695 ;
        RECT 103.820 126.650 104.140 126.710 ;
        RECT 102.915 126.510 104.140 126.650 ;
        RECT 119.090 126.650 119.230 127.145 ;
        RECT 119.920 127.130 120.240 127.390 ;
        RECT 120.395 127.145 120.685 127.375 ;
        RECT 120.840 127.330 121.160 127.390 ;
        RECT 124.980 127.330 125.300 127.390 ;
        RECT 120.840 127.190 125.300 127.330 ;
        RECT 119.460 126.990 119.780 127.050 ;
        RECT 120.470 126.990 120.610 127.145 ;
        RECT 120.840 127.130 121.160 127.190 ;
        RECT 124.980 127.130 125.300 127.190 ;
        RECT 134.640 127.130 134.960 127.390 ;
        RECT 135.100 127.130 135.420 127.390 ;
        RECT 136.110 127.375 136.250 127.530 ;
        RECT 136.940 127.470 137.260 127.530 ;
        RECT 137.415 127.485 137.705 127.715 ;
        RECT 138.295 127.670 138.585 127.715 ;
        RECT 139.485 127.670 139.775 127.715 ;
        RECT 142.005 127.670 142.295 127.715 ;
        RECT 138.295 127.530 142.295 127.670 ;
        RECT 138.295 127.485 138.585 127.530 ;
        RECT 139.485 127.485 139.775 127.530 ;
        RECT 142.005 127.485 142.295 127.530 ;
        RECT 136.035 127.145 136.325 127.375 ;
        RECT 136.495 127.330 136.785 127.375 ;
        RECT 140.620 127.330 140.940 127.390 ;
        RECT 136.495 127.190 140.940 127.330 ;
        RECT 136.495 127.145 136.785 127.190 ;
        RECT 140.620 127.130 140.940 127.190 ;
        RECT 119.460 126.850 120.610 126.990 ;
        RECT 121.300 126.990 121.620 127.050 ;
        RECT 122.080 126.990 122.370 127.035 ;
        RECT 138.640 126.990 138.930 127.035 ;
        RECT 121.300 126.850 122.370 126.990 ;
        RECT 119.460 126.790 119.780 126.850 ;
        RECT 121.300 126.790 121.620 126.850 ;
        RECT 122.080 126.805 122.370 126.850 ;
        RECT 132.890 126.850 138.930 126.990 ;
        RECT 127.755 126.650 128.045 126.695 ;
        RECT 129.120 126.650 129.440 126.710 ;
        RECT 132.890 126.695 133.030 126.850 ;
        RECT 138.640 126.805 138.930 126.850 ;
        RECT 119.090 126.510 129.440 126.650 ;
        RECT 102.915 126.465 103.205 126.510 ;
        RECT 103.820 126.450 104.140 126.510 ;
        RECT 127.755 126.465 128.045 126.510 ;
        RECT 129.120 126.450 129.440 126.510 ;
        RECT 132.815 126.465 133.105 126.695 ;
        RECT 135.100 126.650 135.420 126.710 ;
        RECT 143.840 126.650 144.160 126.710 ;
        RECT 144.315 126.650 144.605 126.695 ;
        RECT 135.100 126.510 144.605 126.650 ;
        RECT 135.100 126.450 135.420 126.510 ;
        RECT 143.840 126.450 144.160 126.510 ;
        RECT 144.315 126.465 144.605 126.510 ;
        RECT 17.270 125.830 146.990 126.310 ;
        RECT 22.875 125.630 23.165 125.675 ;
        RECT 25.620 125.630 25.940 125.690 ;
        RECT 22.875 125.490 25.940 125.630 ;
        RECT 22.875 125.445 23.165 125.490 ;
        RECT 25.620 125.430 25.940 125.490 ;
        RECT 101.980 125.430 102.300 125.690 ;
        RECT 115.780 125.430 116.100 125.690 ;
        RECT 126.820 125.430 127.140 125.690 ;
        RECT 128.200 125.630 128.520 125.690 ;
        RECT 128.675 125.630 128.965 125.675 ;
        RECT 128.200 125.490 128.965 125.630 ;
        RECT 128.200 125.430 128.520 125.490 ;
        RECT 128.675 125.445 128.965 125.490 ;
        RECT 131.880 125.630 132.200 125.690 ;
        RECT 131.880 125.490 133.030 125.630 ;
        RECT 131.880 125.430 132.200 125.490 ;
        RECT 96.460 125.335 96.780 125.350 ;
        RECT 28.550 125.290 28.840 125.335 ;
        RECT 30.235 125.290 30.525 125.335 ;
        RECT 96.430 125.290 96.780 125.335 ;
        RECT 28.550 125.150 30.525 125.290 ;
        RECT 96.265 125.150 96.780 125.290 ;
        RECT 28.550 125.105 28.840 125.150 ;
        RECT 30.235 125.105 30.525 125.150 ;
        RECT 96.430 125.105 96.780 125.150 ;
        RECT 96.460 125.090 96.780 125.105 ;
        RECT 20.100 124.750 20.420 125.010 ;
        RECT 26.080 124.950 26.400 125.010 ;
        RECT 29.775 124.950 30.065 124.995 ;
        RECT 26.080 124.810 30.065 124.950 ;
        RECT 26.080 124.750 26.400 124.810 ;
        RECT 29.775 124.765 30.065 124.810 ;
        RECT 31.600 124.750 31.920 125.010 ;
        RECT 33.915 124.950 34.205 124.995 ;
        RECT 35.280 124.950 35.600 125.010 ;
        RECT 33.915 124.810 35.600 124.950 ;
        RECT 33.915 124.765 34.205 124.810 ;
        RECT 35.280 124.750 35.600 124.810 ;
        RECT 86.800 124.950 87.120 125.010 ;
        RECT 88.640 124.950 88.960 125.010 ;
        RECT 86.800 124.810 88.960 124.950 ;
        RECT 86.800 124.750 87.120 124.810 ;
        RECT 88.640 124.750 88.960 124.810 ;
        RECT 89.560 124.750 89.880 125.010 ;
        RECT 102.070 124.950 102.210 125.430 ;
        RECT 102.455 125.290 102.745 125.335 ;
        RECT 104.280 125.290 104.600 125.350 ;
        RECT 102.455 125.150 104.600 125.290 ;
        RECT 102.455 125.105 102.745 125.150 ;
        RECT 104.280 125.090 104.600 125.150 ;
        RECT 118.080 125.290 118.400 125.350 ;
        RECT 120.380 125.290 120.700 125.350 ;
        RECT 121.775 125.290 122.065 125.335 ;
        RECT 118.080 125.150 122.065 125.290 ;
        RECT 118.080 125.090 118.400 125.150 ;
        RECT 120.380 125.090 120.700 125.150 ;
        RECT 121.775 125.105 122.065 125.150 ;
        RECT 124.980 125.290 125.300 125.350 ;
        RECT 125.455 125.290 125.745 125.335 ;
        RECT 132.890 125.290 133.030 125.490 ;
        RECT 144.760 125.430 145.080 125.690 ;
        RECT 133.580 125.290 133.870 125.335 ;
        RECT 124.980 125.150 132.570 125.290 ;
        RECT 132.890 125.150 133.870 125.290 ;
        RECT 124.980 125.090 125.300 125.150 ;
        RECT 125.455 125.105 125.745 125.150 ;
        RECT 103.375 124.950 103.665 124.995 ;
        RECT 102.070 124.810 103.665 124.950 ;
        RECT 103.375 124.765 103.665 124.810 ;
        RECT 103.820 124.750 104.140 125.010 ;
        RECT 114.860 124.950 115.180 125.010 ;
        RECT 129.120 124.950 129.440 125.010 ;
        RECT 132.430 124.995 132.570 125.150 ;
        RECT 133.580 125.105 133.870 125.150 ;
        RECT 134.270 125.150 144.070 125.290 ;
        RECT 114.860 124.810 117.390 124.950 ;
        RECT 114.860 124.750 115.180 124.810 ;
        RECT 25.185 124.610 25.475 124.655 ;
        RECT 27.705 124.610 27.995 124.655 ;
        RECT 28.895 124.610 29.185 124.655 ;
        RECT 25.185 124.470 29.185 124.610 ;
        RECT 25.185 124.425 25.475 124.470 ;
        RECT 27.705 124.425 27.995 124.470 ;
        RECT 28.895 124.425 29.185 124.470 ;
        RECT 31.140 124.610 31.460 124.670 ;
        RECT 32.075 124.610 32.365 124.655 ;
        RECT 31.140 124.470 32.365 124.610 ;
        RECT 31.140 124.410 31.460 124.470 ;
        RECT 32.075 124.425 32.365 124.470 ;
        RECT 32.535 124.610 32.825 124.655 ;
        RECT 34.820 124.610 35.140 124.670 ;
        RECT 32.535 124.470 35.140 124.610 ;
        RECT 32.535 124.425 32.825 124.470 ;
        RECT 34.820 124.410 35.140 124.470 ;
        RECT 87.720 124.610 88.040 124.670 ;
        RECT 93.240 124.610 93.560 124.670 ;
        RECT 95.095 124.610 95.385 124.655 ;
        RECT 87.720 124.470 95.385 124.610 ;
        RECT 87.720 124.410 88.040 124.470 ;
        RECT 93.240 124.410 93.560 124.470 ;
        RECT 95.095 124.425 95.385 124.470 ;
        RECT 95.975 124.610 96.265 124.655 ;
        RECT 97.165 124.610 97.455 124.655 ;
        RECT 99.685 124.610 99.975 124.655 ;
        RECT 95.975 124.470 99.975 124.610 ;
        RECT 95.975 124.425 96.265 124.470 ;
        RECT 97.165 124.425 97.455 124.470 ;
        RECT 99.685 124.425 99.975 124.470 ;
        RECT 116.240 124.410 116.560 124.670 ;
        RECT 117.250 124.655 117.390 124.810 ;
        RECT 129.120 124.810 130.730 124.950 ;
        RECT 129.120 124.750 129.440 124.810 ;
        RECT 117.175 124.610 117.465 124.655 ;
        RECT 130.055 124.610 130.345 124.655 ;
        RECT 117.175 124.470 130.345 124.610 ;
        RECT 130.590 124.610 130.730 124.810 ;
        RECT 132.355 124.765 132.645 124.995 ;
        RECT 134.270 124.950 134.410 125.150 ;
        RECT 143.930 124.995 144.070 125.150 ;
        RECT 142.015 124.950 142.305 124.995 ;
        RECT 132.890 124.810 134.410 124.950 ;
        RECT 139.330 124.810 142.305 124.950 ;
        RECT 132.890 124.610 133.030 124.810 ;
        RECT 130.590 124.470 133.030 124.610 ;
        RECT 133.235 124.610 133.525 124.655 ;
        RECT 134.425 124.610 134.715 124.655 ;
        RECT 136.945 124.610 137.235 124.655 ;
        RECT 133.235 124.470 137.235 124.610 ;
        RECT 117.175 124.425 117.465 124.470 ;
        RECT 130.055 124.425 130.345 124.470 ;
        RECT 133.235 124.425 133.525 124.470 ;
        RECT 134.425 124.425 134.715 124.470 ;
        RECT 136.945 124.425 137.235 124.470 ;
        RECT 15.880 124.320 16.160 124.350 ;
        RECT 14.970 124.040 16.160 124.320 ;
        RECT 25.620 124.270 25.910 124.315 ;
        RECT 27.190 124.270 27.480 124.315 ;
        RECT 29.290 124.270 29.580 124.315 ;
        RECT 32.995 124.270 33.285 124.315 ;
        RECT 25.620 124.130 29.580 124.270 ;
        RECT 25.620 124.085 25.910 124.130 ;
        RECT 27.190 124.085 27.480 124.130 ;
        RECT 29.290 124.085 29.580 124.130 ;
        RECT 31.690 124.130 33.285 124.270 ;
        RECT 15.480 123.980 16.160 124.040 ;
        RECT 15.480 123.380 16.180 123.980 ;
        RECT 19.180 123.930 19.500 123.990 ;
        RECT 20.575 123.930 20.865 123.975 ;
        RECT 26.080 123.930 26.400 123.990 ;
        RECT 19.180 123.790 26.400 123.930 ;
        RECT 19.180 123.730 19.500 123.790 ;
        RECT 20.575 123.745 20.865 123.790 ;
        RECT 26.080 123.730 26.400 123.790 ;
        RECT 29.760 123.930 30.080 123.990 ;
        RECT 31.690 123.930 31.830 124.130 ;
        RECT 32.995 124.085 33.285 124.130 ;
        RECT 95.580 124.270 95.870 124.315 ;
        RECT 97.680 124.270 97.970 124.315 ;
        RECT 99.250 124.270 99.540 124.315 ;
        RECT 95.580 124.130 99.540 124.270 ;
        RECT 95.580 124.085 95.870 124.130 ;
        RECT 97.680 124.085 97.970 124.130 ;
        RECT 99.250 124.085 99.540 124.130 ;
        RECT 103.835 124.085 104.125 124.315 ;
        RECT 130.130 124.270 130.270 124.425 ;
        RECT 139.330 124.330 139.470 124.810 ;
        RECT 142.015 124.765 142.305 124.810 ;
        RECT 143.855 124.765 144.145 124.995 ;
        RECT 132.840 124.270 133.130 124.315 ;
        RECT 134.940 124.270 135.230 124.315 ;
        RECT 136.510 124.270 136.800 124.315 ;
        RECT 138.320 124.270 138.640 124.330 ;
        RECT 113.570 124.130 114.630 124.270 ;
        RECT 130.130 124.130 132.570 124.270 ;
        RECT 29.760 123.790 31.830 123.930 ;
        RECT 101.520 123.930 101.840 123.990 ;
        RECT 103.910 123.930 104.050 124.085 ;
        RECT 113.570 123.930 113.710 124.130 ;
        RECT 101.520 123.790 113.710 123.930 ;
        RECT 29.760 123.730 30.080 123.790 ;
        RECT 101.520 123.730 101.840 123.790 ;
        RECT 113.940 123.730 114.260 123.990 ;
        RECT 114.490 123.930 114.630 124.130 ;
        RECT 130.960 123.930 131.280 123.990 ;
        RECT 114.490 123.790 131.280 123.930 ;
        RECT 132.430 123.930 132.570 124.130 ;
        RECT 132.840 124.130 136.800 124.270 ;
        RECT 132.840 124.085 133.130 124.130 ;
        RECT 134.940 124.085 135.230 124.130 ;
        RECT 136.510 124.085 136.800 124.130 ;
        RECT 137.030 124.130 138.640 124.270 ;
        RECT 137.030 123.930 137.170 124.130 ;
        RECT 138.320 124.070 138.640 124.130 ;
        RECT 139.240 124.070 139.560 124.330 ;
        RECT 142.920 124.070 143.240 124.330 ;
        RECT 132.430 123.790 137.170 123.930 ;
        RECT 130.960 123.730 131.280 123.790 ;
        RECT 17.270 123.110 146.990 123.590 ;
        RECT 28.840 122.910 29.160 122.970 ;
        RECT 35.280 122.910 35.600 122.970 ;
        RECT 28.470 122.770 35.600 122.910 ;
        RECT 28.470 122.615 28.610 122.770 ;
        RECT 28.840 122.710 29.160 122.770 ;
        RECT 35.280 122.710 35.600 122.770 ;
        RECT 91.860 122.910 92.180 122.970 ;
        RECT 105.660 122.910 105.980 122.970 ;
        RECT 107.975 122.910 108.265 122.955 ;
        RECT 91.860 122.770 105.430 122.910 ;
        RECT 91.860 122.710 92.180 122.770 ;
        RECT 14.650 122.470 15.360 122.610 ;
        RECT 15.220 113.050 15.360 122.470 ;
        RECT 19.680 122.570 19.970 122.615 ;
        RECT 21.780 122.570 22.070 122.615 ;
        RECT 23.350 122.570 23.640 122.615 ;
        RECT 19.680 122.430 23.640 122.570 ;
        RECT 19.680 122.385 19.970 122.430 ;
        RECT 21.780 122.385 22.070 122.430 ;
        RECT 23.350 122.385 23.640 122.430 ;
        RECT 28.395 122.385 28.685 122.615 ;
        RECT 31.180 122.570 31.470 122.615 ;
        RECT 33.280 122.570 33.570 122.615 ;
        RECT 34.850 122.570 35.140 122.615 ;
        RECT 31.180 122.430 35.140 122.570 ;
        RECT 31.180 122.385 31.470 122.430 ;
        RECT 33.280 122.385 33.570 122.430 ;
        RECT 34.850 122.385 35.140 122.430 ;
        RECT 88.640 122.370 88.960 122.630 ;
        RECT 105.290 122.615 105.430 122.770 ;
        RECT 105.660 122.770 108.265 122.910 ;
        RECT 105.660 122.710 105.980 122.770 ;
        RECT 107.975 122.725 108.265 122.770 ;
        RECT 115.320 122.910 115.640 122.970 ;
        RECT 131.420 122.910 131.740 122.970 ;
        RECT 132.815 122.910 133.105 122.955 ;
        RECT 115.320 122.770 120.150 122.910 ;
        RECT 115.320 122.710 115.640 122.770 ;
        RECT 120.010 122.630 120.150 122.770 ;
        RECT 131.420 122.770 133.105 122.910 ;
        RECT 131.420 122.710 131.740 122.770 ;
        RECT 132.815 122.725 133.105 122.770 ;
        RECT 133.720 122.710 134.040 122.970 ;
        RECT 93.740 122.570 94.030 122.615 ;
        RECT 95.840 122.570 96.130 122.615 ;
        RECT 97.410 122.570 97.700 122.615 ;
        RECT 93.740 122.430 97.700 122.570 ;
        RECT 93.740 122.385 94.030 122.430 ;
        RECT 95.840 122.385 96.130 122.430 ;
        RECT 97.410 122.385 97.700 122.430 ;
        RECT 100.155 122.570 100.445 122.615 ;
        RECT 100.155 122.430 103.590 122.570 ;
        RECT 100.155 122.385 100.445 122.430 ;
        RECT 19.180 122.030 19.500 122.290 ;
        RECT 20.075 122.230 20.365 122.275 ;
        RECT 21.265 122.230 21.555 122.275 ;
        RECT 23.785 122.230 24.075 122.275 ;
        RECT 20.075 122.090 24.075 122.230 ;
        RECT 20.075 122.045 20.365 122.090 ;
        RECT 21.265 122.045 21.555 122.090 ;
        RECT 23.785 122.045 24.075 122.090 ;
        RECT 31.575 122.230 31.865 122.275 ;
        RECT 32.765 122.230 33.055 122.275 ;
        RECT 35.285 122.230 35.575 122.275 ;
        RECT 31.575 122.090 35.575 122.230 ;
        RECT 31.575 122.045 31.865 122.090 ;
        RECT 32.765 122.045 33.055 122.090 ;
        RECT 35.285 122.045 35.575 122.090 ;
        RECT 93.240 122.030 93.560 122.290 ;
        RECT 94.135 122.230 94.425 122.275 ;
        RECT 95.325 122.230 95.615 122.275 ;
        RECT 97.845 122.230 98.135 122.275 ;
        RECT 94.135 122.090 98.135 122.230 ;
        RECT 94.135 122.045 94.425 122.090 ;
        RECT 95.325 122.045 95.615 122.090 ;
        RECT 97.845 122.045 98.135 122.090 ;
        RECT 26.080 121.890 26.400 121.950 ;
        RECT 30.695 121.890 30.985 121.935 ;
        RECT 26.080 121.750 30.985 121.890 ;
        RECT 26.080 121.690 26.400 121.750 ;
        RECT 30.695 121.705 30.985 121.750 ;
        RECT 92.335 121.890 92.625 121.935 ;
        RECT 93.330 121.890 93.470 122.030 ;
        RECT 92.335 121.750 93.470 121.890 ;
        RECT 94.590 121.890 94.880 121.935 ;
        RECT 99.220 121.890 99.540 121.950 ;
        RECT 94.590 121.750 99.540 121.890 ;
        RECT 92.335 121.705 92.625 121.750 ;
        RECT 94.590 121.705 94.880 121.750 ;
        RECT 99.220 121.690 99.540 121.750 ;
        RECT 100.615 121.890 100.905 121.935 ;
        RECT 101.980 121.890 102.300 121.950 ;
        RECT 103.450 121.935 103.590 122.430 ;
        RECT 105.215 122.385 105.505 122.615 ;
        RECT 113.980 122.570 114.270 122.615 ;
        RECT 116.080 122.570 116.370 122.615 ;
        RECT 117.650 122.570 117.940 122.615 ;
        RECT 113.980 122.430 117.940 122.570 ;
        RECT 113.980 122.385 114.270 122.430 ;
        RECT 116.080 122.385 116.370 122.430 ;
        RECT 117.650 122.385 117.940 122.430 ;
        RECT 119.920 122.570 120.240 122.630 ;
        RECT 141.540 122.570 141.860 122.630 ;
        RECT 119.920 122.430 141.860 122.570 ;
        RECT 119.920 122.370 120.240 122.430 ;
        RECT 108.420 122.230 108.740 122.290 ;
        RECT 114.375 122.230 114.665 122.275 ;
        RECT 115.565 122.230 115.855 122.275 ;
        RECT 118.085 122.230 118.375 122.275 ;
        RECT 108.420 122.090 110.490 122.230 ;
        RECT 108.420 122.030 108.740 122.090 ;
        RECT 100.615 121.750 102.300 121.890 ;
        RECT 100.615 121.705 100.905 121.750 ;
        RECT 101.980 121.690 102.300 121.750 ;
        RECT 103.375 121.890 103.665 121.935 ;
        RECT 103.820 121.890 104.140 121.950 ;
        RECT 103.375 121.750 104.140 121.890 ;
        RECT 103.375 121.705 103.665 121.750 ;
        RECT 103.820 121.690 104.140 121.750 ;
        RECT 104.280 121.890 104.600 121.950 ;
        RECT 110.350 121.935 110.490 122.090 ;
        RECT 114.375 122.090 118.375 122.230 ;
        RECT 114.375 122.045 114.665 122.090 ;
        RECT 115.565 122.045 115.855 122.090 ;
        RECT 118.085 122.045 118.375 122.090 ;
        RECT 108.895 121.890 109.185 121.935 ;
        RECT 104.280 121.750 109.185 121.890 ;
        RECT 104.280 121.690 104.600 121.750 ;
        RECT 108.895 121.705 109.185 121.750 ;
        RECT 109.355 121.705 109.645 121.935 ;
        RECT 110.275 121.705 110.565 121.935 ;
        RECT 20.530 121.550 20.820 121.595 ;
        RECT 21.480 121.550 21.800 121.610 ;
        RECT 20.530 121.410 21.800 121.550 ;
        RECT 20.530 121.365 20.820 121.410 ;
        RECT 21.480 121.350 21.800 121.410 ;
        RECT 29.760 121.350 30.080 121.610 ;
        RECT 32.060 121.595 32.380 121.610 ;
        RECT 31.920 121.550 32.380 121.595 ;
        RECT 30.310 121.410 32.380 121.550 ;
        RECT 21.940 121.210 22.260 121.270 ;
        RECT 26.095 121.210 26.385 121.255 ;
        RECT 21.940 121.070 26.385 121.210 ;
        RECT 21.940 121.010 22.260 121.070 ;
        RECT 26.095 121.025 26.385 121.070 ;
        RECT 27.460 121.210 27.780 121.270 ;
        RECT 30.310 121.210 30.450 121.410 ;
        RECT 31.920 121.365 32.380 121.410 ;
        RECT 32.060 121.350 32.380 121.365 ;
        RECT 85.880 121.550 86.200 121.610 ;
        RECT 86.815 121.550 87.105 121.595 ;
        RECT 106.135 121.550 106.425 121.595 ;
        RECT 85.880 121.410 87.105 121.550 ;
        RECT 85.880 121.350 86.200 121.410 ;
        RECT 86.815 121.365 87.105 121.410 ;
        RECT 104.370 121.410 106.425 121.550 ;
        RECT 109.430 121.550 109.570 121.705 ;
        RECT 110.720 121.690 111.040 121.950 ;
        RECT 113.480 121.690 113.800 121.950 ;
        RECT 116.240 121.890 116.560 121.950 ;
        RECT 114.490 121.750 116.560 121.890 ;
        RECT 114.490 121.550 114.630 121.750 ;
        RECT 116.240 121.690 116.560 121.750 ;
        RECT 120.380 121.890 120.700 121.950 ;
        RECT 120.855 121.890 121.145 121.935 ;
        RECT 120.380 121.750 121.145 121.890 ;
        RECT 120.380 121.690 120.700 121.750 ;
        RECT 120.855 121.705 121.145 121.750 ;
        RECT 129.120 121.890 129.440 121.950 ;
        RECT 130.500 121.935 130.820 121.950 ;
        RECT 129.595 121.890 129.885 121.935 ;
        RECT 129.120 121.750 129.885 121.890 ;
        RECT 129.120 121.690 129.440 121.750 ;
        RECT 129.595 121.705 129.885 121.750 ;
        RECT 130.335 121.705 130.820 121.935 ;
        RECT 131.920 121.890 132.210 121.935 ;
        RECT 132.430 121.890 132.570 122.430 ;
        RECT 141.540 122.370 141.860 122.430 ;
        RECT 133.260 122.230 133.580 122.290 ;
        RECT 133.260 122.090 135.790 122.230 ;
        RECT 133.260 122.030 133.580 122.090 ;
        RECT 135.650 121.935 135.790 122.090 ;
        RECT 136.020 122.030 136.340 122.290 ;
        RECT 136.955 122.230 137.245 122.275 ;
        RECT 139.700 122.230 140.020 122.290 ;
        RECT 136.955 122.090 140.020 122.230 ;
        RECT 136.955 122.045 137.245 122.090 ;
        RECT 139.700 122.030 140.020 122.090 ;
        RECT 131.920 121.750 132.570 121.890 ;
        RECT 131.920 121.705 132.210 121.750 ;
        RECT 135.575 121.705 135.865 121.935 ;
        RECT 136.110 121.890 136.250 122.030 ;
        RECT 142.015 121.890 142.305 121.935 ;
        RECT 136.110 121.750 142.305 121.890 ;
        RECT 142.015 121.705 142.305 121.750 ;
        RECT 130.500 121.690 130.820 121.705 ;
        RECT 143.840 121.690 144.160 121.950 ;
        RECT 114.860 121.595 115.180 121.610 ;
        RECT 109.430 121.410 114.630 121.550 ;
        RECT 27.460 121.070 30.450 121.210 ;
        RECT 34.820 121.210 35.140 121.270 ;
        RECT 37.595 121.210 37.885 121.255 ;
        RECT 34.820 121.070 37.885 121.210 ;
        RECT 27.460 121.010 27.780 121.070 ;
        RECT 34.820 121.010 35.140 121.070 ;
        RECT 37.595 121.025 37.885 121.070 ;
        RECT 88.180 121.210 88.500 121.270 ;
        RECT 104.370 121.255 104.510 121.410 ;
        RECT 106.135 121.365 106.425 121.410 ;
        RECT 114.830 121.365 115.180 121.595 ;
        RECT 89.115 121.210 89.405 121.255 ;
        RECT 88.180 121.070 89.405 121.210 ;
        RECT 88.180 121.010 88.500 121.070 ;
        RECT 89.115 121.025 89.405 121.070 ;
        RECT 104.295 121.025 104.585 121.255 ;
        RECT 106.210 121.210 106.350 121.365 ;
        RECT 114.860 121.350 115.180 121.365 ;
        RECT 115.320 121.210 115.640 121.270 ;
        RECT 106.210 121.070 115.640 121.210 ;
        RECT 116.330 121.210 116.470 121.690 ;
        RECT 124.520 121.350 124.840 121.610 ;
        RECT 130.960 121.350 131.280 121.610 ;
        RECT 131.435 121.550 131.725 121.595 ;
        RECT 136.035 121.550 136.325 121.595 ;
        RECT 139.240 121.550 139.560 121.610 ;
        RECT 131.435 121.410 139.560 121.550 ;
        RECT 131.435 121.365 131.725 121.410 ;
        RECT 136.035 121.365 136.325 121.410 ;
        RECT 139.240 121.350 139.560 121.410 ;
        RECT 120.395 121.210 120.685 121.255 ;
        RECT 129.580 121.210 129.900 121.270 ;
        RECT 116.330 121.070 129.900 121.210 ;
        RECT 131.050 121.210 131.190 121.350 ;
        RECT 142.460 121.210 142.780 121.270 ;
        RECT 131.050 121.070 142.780 121.210 ;
        RECT 115.320 121.010 115.640 121.070 ;
        RECT 120.395 121.025 120.685 121.070 ;
        RECT 129.580 121.010 129.900 121.070 ;
        RECT 142.460 121.010 142.780 121.070 ;
        RECT 142.920 121.010 143.240 121.270 ;
        RECT 144.760 121.010 145.080 121.270 ;
        RECT 17.270 120.390 146.990 120.870 ;
        RECT 20.100 120.190 20.420 120.250 ;
        RECT 21.035 120.190 21.325 120.235 ;
        RECT 20.100 120.050 21.325 120.190 ;
        RECT 20.100 119.990 20.420 120.050 ;
        RECT 21.035 120.005 21.325 120.050 ;
        RECT 21.480 119.990 21.800 120.250 ;
        RECT 21.940 120.190 22.260 120.250 ;
        RECT 23.335 120.190 23.625 120.235 ;
        RECT 21.940 120.050 23.625 120.190 ;
        RECT 21.940 119.990 22.260 120.050 ;
        RECT 23.335 120.005 23.625 120.050 ;
        RECT 23.795 120.190 24.085 120.235 ;
        RECT 24.240 120.190 24.560 120.250 ;
        RECT 23.795 120.050 24.560 120.190 ;
        RECT 23.795 120.005 24.085 120.050 ;
        RECT 24.240 119.990 24.560 120.050 ;
        RECT 32.995 120.005 33.285 120.235 ;
        RECT 33.070 119.850 33.210 120.005 ;
        RECT 35.740 119.990 36.060 120.250 ;
        RECT 79.915 120.190 80.205 120.235 ;
        RECT 80.360 120.190 80.680 120.250 ;
        RECT 86.340 120.190 86.660 120.250 ;
        RECT 90.020 120.190 90.340 120.250 ;
        RECT 101.520 120.190 101.840 120.250 ;
        RECT 79.915 120.050 90.340 120.190 ;
        RECT 79.915 120.005 80.205 120.050 ;
        RECT 80.360 119.990 80.680 120.050 ;
        RECT 86.340 119.990 86.660 120.050 ;
        RECT 90.020 119.990 90.340 120.050 ;
        RECT 97.470 120.050 101.840 120.190 ;
        RECT 33.455 119.850 33.745 119.895 ;
        RECT 35.280 119.850 35.600 119.910 ;
        RECT 33.070 119.710 35.600 119.850 ;
        RECT 33.455 119.665 33.745 119.710 ;
        RECT 35.280 119.650 35.600 119.710 ;
        RECT 15.960 119.510 16.280 119.570 ;
        RECT 18.735 119.510 19.025 119.555 ;
        RECT 15.960 119.370 19.025 119.510 ;
        RECT 15.960 119.310 16.280 119.370 ;
        RECT 18.735 119.325 19.025 119.370 ;
        RECT 20.100 119.310 20.420 119.570 ;
        RECT 26.540 119.510 26.860 119.570 ;
        RECT 27.430 119.510 27.720 119.555 ;
        RECT 29.300 119.510 29.620 119.570 ;
        RECT 24.790 119.370 29.620 119.510 ;
        RECT 24.790 119.215 24.930 119.370 ;
        RECT 26.540 119.310 26.860 119.370 ;
        RECT 27.430 119.325 27.720 119.370 ;
        RECT 29.300 119.310 29.620 119.370 ;
        RECT 30.220 119.510 30.540 119.570 ;
        RECT 35.830 119.510 35.970 119.990 ;
        RECT 83.580 119.850 83.900 119.910 ;
        RECT 83.580 119.710 92.090 119.850 ;
        RECT 83.580 119.650 83.900 119.710 ;
        RECT 91.950 119.570 92.090 119.710 ;
        RECT 30.220 119.370 35.970 119.510 ;
        RECT 78.980 119.510 79.300 119.570 ;
        RECT 86.815 119.510 87.105 119.555 ;
        RECT 89.100 119.510 89.420 119.570 ;
        RECT 78.980 119.370 81.050 119.510 ;
        RECT 30.220 119.310 30.540 119.370 ;
        RECT 78.980 119.310 79.300 119.370 ;
        RECT 24.715 118.985 25.005 119.215 ;
        RECT 26.080 118.970 26.400 119.230 ;
        RECT 26.975 119.170 27.265 119.215 ;
        RECT 28.165 119.170 28.455 119.215 ;
        RECT 30.685 119.170 30.975 119.215 ;
        RECT 26.975 119.030 30.975 119.170 ;
        RECT 26.975 118.985 27.265 119.030 ;
        RECT 28.165 118.985 28.455 119.030 ;
        RECT 30.685 118.985 30.975 119.030 ;
        RECT 34.360 119.170 34.680 119.230 ;
        RECT 35.280 119.170 35.600 119.230 ;
        RECT 34.360 119.030 35.600 119.170 ;
        RECT 34.360 118.970 34.680 119.030 ;
        RECT 35.280 118.970 35.600 119.030 ;
        RECT 73.920 118.970 74.240 119.230 ;
        RECT 80.910 119.215 81.050 119.370 ;
        RECT 86.815 119.370 89.420 119.510 ;
        RECT 86.815 119.325 87.105 119.370 ;
        RECT 89.100 119.310 89.420 119.370 ;
        RECT 91.860 119.310 92.180 119.570 ;
        RECT 93.700 119.310 94.020 119.570 ;
        RECT 97.470 119.555 97.610 120.050 ;
        RECT 101.520 119.990 101.840 120.050 ;
        RECT 105.200 120.190 105.520 120.250 ;
        RECT 109.355 120.190 109.645 120.235 ;
        RECT 105.200 120.050 114.630 120.190 ;
        RECT 105.200 119.990 105.520 120.050 ;
        RECT 109.355 120.005 109.645 120.050 ;
        RECT 100.615 119.665 100.905 119.895 ;
        RECT 104.280 119.850 104.600 119.910 ;
        RECT 106.135 119.850 106.425 119.895 ;
        RECT 102.070 119.710 104.050 119.850 ;
        RECT 97.395 119.325 97.685 119.555 ;
        RECT 98.315 119.325 98.605 119.555 ;
        RECT 100.155 119.325 100.445 119.555 ;
        RECT 100.690 119.510 100.830 119.665 ;
        RECT 101.520 119.510 101.840 119.570 ;
        RECT 102.070 119.555 102.210 119.710 ;
        RECT 103.910 119.570 104.050 119.710 ;
        RECT 104.280 119.710 106.425 119.850 ;
        RECT 104.280 119.650 104.600 119.710 ;
        RECT 106.135 119.665 106.425 119.710 ;
        RECT 108.880 119.850 109.200 119.910 ;
        RECT 112.575 119.850 112.865 119.895 ;
        RECT 108.880 119.710 112.865 119.850 ;
        RECT 114.490 119.850 114.630 120.050 ;
        RECT 114.860 119.990 115.180 120.250 ;
        RECT 128.215 120.190 128.505 120.235 ;
        RECT 130.500 120.190 130.820 120.250 ;
        RECT 130.975 120.190 131.265 120.235 ;
        RECT 136.020 120.190 136.340 120.250 ;
        RECT 128.215 120.050 136.340 120.190 ;
        RECT 128.215 120.005 128.505 120.050 ;
        RECT 130.500 119.990 130.820 120.050 ;
        RECT 130.975 120.005 131.265 120.050 ;
        RECT 136.020 119.990 136.340 120.050 ;
        RECT 136.955 120.005 137.245 120.235 ;
        RECT 122.650 119.850 122.940 119.895 ;
        RECT 123.600 119.850 123.920 119.910 ;
        RECT 114.490 119.710 122.220 119.850 ;
        RECT 108.880 119.650 109.200 119.710 ;
        RECT 112.575 119.665 112.865 119.710 ;
        RECT 100.690 119.370 101.840 119.510 ;
        RECT 80.375 118.985 80.665 119.215 ;
        RECT 80.835 118.985 81.125 119.215 ;
        RECT 85.420 119.170 85.740 119.230 ;
        RECT 87.275 119.170 87.565 119.215 ;
        RECT 95.080 119.170 95.400 119.230 ;
        RECT 85.420 119.030 95.400 119.170 ;
        RECT 19.655 118.830 19.945 118.875 ;
        RECT 26.580 118.830 26.870 118.875 ;
        RECT 28.680 118.830 28.970 118.875 ;
        RECT 30.250 118.830 30.540 118.875 ;
        RECT 34.820 118.830 35.140 118.890 ;
        RECT 19.655 118.690 25.620 118.830 ;
        RECT 19.655 118.645 19.945 118.690 ;
        RECT 25.480 118.490 25.620 118.690 ;
        RECT 26.580 118.690 30.540 118.830 ;
        RECT 26.580 118.645 26.870 118.690 ;
        RECT 28.680 118.645 28.970 118.690 ;
        RECT 30.250 118.645 30.540 118.690 ;
        RECT 32.610 118.690 35.140 118.830 ;
        RECT 27.920 118.490 28.240 118.550 ;
        RECT 25.480 118.350 28.240 118.490 ;
        RECT 27.920 118.290 28.240 118.350 ;
        RECT 29.760 118.490 30.080 118.550 ;
        RECT 32.610 118.490 32.750 118.690 ;
        RECT 34.820 118.630 35.140 118.690 ;
        RECT 75.775 118.830 76.065 118.875 ;
        RECT 78.075 118.830 78.365 118.875 ;
        RECT 75.775 118.690 78.365 118.830 ;
        RECT 75.775 118.645 76.065 118.690 ;
        RECT 78.075 118.645 78.365 118.690 ;
        RECT 79.900 118.830 80.220 118.890 ;
        RECT 80.450 118.830 80.590 118.985 ;
        RECT 85.420 118.970 85.740 119.030 ;
        RECT 87.275 118.985 87.565 119.030 ;
        RECT 95.080 118.970 95.400 119.030 ;
        RECT 79.900 118.690 80.590 118.830 ;
        RECT 87.720 118.830 88.040 118.890 ;
        RECT 90.955 118.830 91.245 118.875 ;
        RECT 98.390 118.830 98.530 119.325 ;
        RECT 100.230 119.170 100.370 119.325 ;
        RECT 101.520 119.310 101.840 119.370 ;
        RECT 101.995 119.325 102.285 119.555 ;
        RECT 102.440 119.510 102.760 119.570 ;
        RECT 103.375 119.510 103.665 119.555 ;
        RECT 102.440 119.370 103.665 119.510 ;
        RECT 102.440 119.310 102.760 119.370 ;
        RECT 103.375 119.325 103.665 119.370 ;
        RECT 103.820 119.310 104.140 119.570 ;
        RECT 120.840 119.510 121.160 119.570 ;
        RECT 121.315 119.510 121.605 119.555 ;
        RECT 120.840 119.370 121.605 119.510 ;
        RECT 122.080 119.510 122.220 119.710 ;
        RECT 122.650 119.710 123.920 119.850 ;
        RECT 122.650 119.665 122.940 119.710 ;
        RECT 123.600 119.650 123.920 119.710 ;
        RECT 134.180 119.850 134.500 119.910 ;
        RECT 134.655 119.850 134.945 119.895 ;
        RECT 134.180 119.710 134.945 119.850 ;
        RECT 137.030 119.850 137.170 120.005 ;
        RECT 138.640 119.850 138.930 119.895 ;
        RECT 137.030 119.710 138.930 119.850 ;
        RECT 134.180 119.650 134.500 119.710 ;
        RECT 134.655 119.665 134.945 119.710 ;
        RECT 138.640 119.665 138.930 119.710 ;
        RECT 130.515 119.510 130.805 119.555 ;
        RECT 133.260 119.510 133.580 119.570 ;
        RECT 122.080 119.370 133.580 119.510 ;
        RECT 120.840 119.310 121.160 119.370 ;
        RECT 121.315 119.325 121.605 119.370 ;
        RECT 130.515 119.325 130.805 119.370 ;
        RECT 133.260 119.310 133.580 119.370 ;
        RECT 102.530 119.170 102.670 119.310 ;
        RECT 100.230 119.030 102.670 119.170 ;
        RECT 105.200 119.170 105.520 119.230 ;
        RECT 105.675 119.170 105.965 119.215 ;
        RECT 105.200 119.030 105.965 119.170 ;
        RECT 105.200 118.970 105.520 119.030 ;
        RECT 105.675 118.985 105.965 119.030 ;
        RECT 106.120 119.170 106.440 119.230 ;
        RECT 108.435 119.170 108.725 119.215 ;
        RECT 106.120 119.030 108.725 119.170 ;
        RECT 106.120 118.970 106.440 119.030 ;
        RECT 108.435 118.985 108.725 119.030 ;
        RECT 108.880 118.970 109.200 119.230 ;
        RECT 122.195 119.170 122.485 119.215 ;
        RECT 123.385 119.170 123.675 119.215 ;
        RECT 125.905 119.170 126.195 119.215 ;
        RECT 122.195 119.030 126.195 119.170 ;
        RECT 122.195 118.985 122.485 119.030 ;
        RECT 123.385 118.985 123.675 119.030 ;
        RECT 125.905 118.985 126.195 119.030 ;
        RECT 131.895 119.170 132.185 119.215 ;
        RECT 132.800 119.170 133.120 119.230 ;
        RECT 131.895 119.030 133.120 119.170 ;
        RECT 131.895 118.985 132.185 119.030 ;
        RECT 132.800 118.970 133.120 119.030 ;
        RECT 136.020 119.170 136.340 119.230 ;
        RECT 137.415 119.170 137.705 119.215 ;
        RECT 136.020 119.030 137.705 119.170 ;
        RECT 136.020 118.970 136.340 119.030 ;
        RECT 137.415 118.985 137.705 119.030 ;
        RECT 138.295 119.170 138.585 119.215 ;
        RECT 139.485 119.170 139.775 119.215 ;
        RECT 142.005 119.170 142.295 119.215 ;
        RECT 138.295 119.030 142.295 119.170 ;
        RECT 138.295 118.985 138.585 119.030 ;
        RECT 139.485 118.985 139.775 119.030 ;
        RECT 142.005 118.985 142.295 119.030 ;
        RECT 104.280 118.830 104.600 118.890 ;
        RECT 87.720 118.690 97.150 118.830 ;
        RECT 98.390 118.690 104.600 118.830 ;
        RECT 79.900 118.630 80.220 118.690 ;
        RECT 87.720 118.630 88.040 118.690 ;
        RECT 90.955 118.645 91.245 118.690 ;
        RECT 29.760 118.350 32.750 118.490 ;
        RECT 29.760 118.290 30.080 118.350 ;
        RECT 76.220 118.290 76.540 118.550 ;
        RECT 84.040 118.490 84.360 118.550 ;
        RECT 84.515 118.490 84.805 118.535 ;
        RECT 84.040 118.350 84.805 118.490 ;
        RECT 84.040 118.290 84.360 118.350 ;
        RECT 84.515 118.305 84.805 118.350 ;
        RECT 96.460 118.290 96.780 118.550 ;
        RECT 97.010 118.490 97.150 118.690 ;
        RECT 104.280 118.630 104.600 118.690 ;
        RECT 104.830 118.690 111.870 118.830 ;
        RECT 104.830 118.490 104.970 118.690 ;
        RECT 97.010 118.350 104.970 118.490 ;
        RECT 109.800 118.490 110.120 118.550 ;
        RECT 111.195 118.490 111.485 118.535 ;
        RECT 109.800 118.350 111.485 118.490 ;
        RECT 111.730 118.490 111.870 118.690 ;
        RECT 113.940 118.630 114.260 118.890 ;
        RECT 121.800 118.830 122.090 118.875 ;
        RECT 123.900 118.830 124.190 118.875 ;
        RECT 125.470 118.830 125.760 118.875 ;
        RECT 121.800 118.690 125.760 118.830 ;
        RECT 121.800 118.645 122.090 118.690 ;
        RECT 123.900 118.645 124.190 118.690 ;
        RECT 125.470 118.645 125.760 118.690 ;
        RECT 128.290 118.690 129.350 118.830 ;
        RECT 119.000 118.490 119.320 118.550 ;
        RECT 128.290 118.490 128.430 118.690 ;
        RECT 111.730 118.350 128.430 118.490 ;
        RECT 109.800 118.290 110.120 118.350 ;
        RECT 111.195 118.305 111.485 118.350 ;
        RECT 119.000 118.290 119.320 118.350 ;
        RECT 128.660 118.290 128.980 118.550 ;
        RECT 129.210 118.490 129.350 118.690 ;
        RECT 136.480 118.630 136.800 118.890 ;
        RECT 137.900 118.830 138.190 118.875 ;
        RECT 140.000 118.830 140.290 118.875 ;
        RECT 141.570 118.830 141.860 118.875 ;
        RECT 137.900 118.690 141.860 118.830 ;
        RECT 137.900 118.645 138.190 118.690 ;
        RECT 140.000 118.645 140.290 118.690 ;
        RECT 141.570 118.645 141.860 118.690 ;
        RECT 139.240 118.490 139.560 118.550 ;
        RECT 129.210 118.350 139.560 118.490 ;
        RECT 139.240 118.290 139.560 118.350 ;
        RECT 144.300 118.290 144.620 118.550 ;
        RECT 17.270 117.670 146.990 118.150 ;
        RECT 88.640 117.470 88.960 117.530 ;
        RECT 90.495 117.470 90.785 117.515 ;
        RECT 88.640 117.330 90.785 117.470 ;
        RECT 88.640 117.270 88.960 117.330 ;
        RECT 90.495 117.285 90.785 117.330 ;
        RECT 95.080 117.470 95.400 117.530 ;
        RECT 106.120 117.470 106.440 117.530 ;
        RECT 95.080 117.330 106.440 117.470 ;
        RECT 95.080 117.270 95.400 117.330 ;
        RECT 106.120 117.270 106.440 117.330 ;
        RECT 113.480 117.470 113.800 117.530 ;
        RECT 113.480 117.330 115.090 117.470 ;
        RECT 113.480 117.270 113.800 117.330 ;
        RECT 72.555 116.945 72.845 117.175 ;
        RECT 74.420 117.130 74.710 117.175 ;
        RECT 76.520 117.130 76.810 117.175 ;
        RECT 78.090 117.130 78.380 117.175 ;
        RECT 74.420 116.990 78.380 117.130 ;
        RECT 74.420 116.945 74.710 116.990 ;
        RECT 76.520 116.945 76.810 116.990 ;
        RECT 78.090 116.945 78.380 116.990 ;
        RECT 82.700 117.130 82.990 117.175 ;
        RECT 84.800 117.130 85.090 117.175 ;
        RECT 86.370 117.130 86.660 117.175 ;
        RECT 82.700 116.990 86.660 117.130 ;
        RECT 82.700 116.945 82.990 116.990 ;
        RECT 84.800 116.945 85.090 116.990 ;
        RECT 86.370 116.945 86.660 116.990 ;
        RECT 93.700 117.130 94.020 117.190 ;
        RECT 95.540 117.130 95.860 117.190 ;
        RECT 110.720 117.130 111.010 117.175 ;
        RECT 112.290 117.130 112.580 117.175 ;
        RECT 114.390 117.130 114.680 117.175 ;
        RECT 93.700 116.990 97.150 117.130 ;
        RECT 72.630 116.790 72.770 116.945 ;
        RECT 93.700 116.930 94.020 116.990 ;
        RECT 95.540 116.930 95.860 116.990 ;
        RECT 73.000 116.790 73.320 116.850 ;
        RECT 72.630 116.650 73.320 116.790 ;
        RECT 73.000 116.590 73.320 116.650 ;
        RECT 74.815 116.790 75.105 116.835 ;
        RECT 76.005 116.790 76.295 116.835 ;
        RECT 78.525 116.790 78.815 116.835 ;
        RECT 74.815 116.650 78.815 116.790 ;
        RECT 74.815 116.605 75.105 116.650 ;
        RECT 76.005 116.605 76.295 116.650 ;
        RECT 78.525 116.605 78.815 116.650 ;
        RECT 83.095 116.790 83.385 116.835 ;
        RECT 84.285 116.790 84.575 116.835 ;
        RECT 86.805 116.790 87.095 116.835 ;
        RECT 83.095 116.650 87.095 116.790 ;
        RECT 83.095 116.605 83.385 116.650 ;
        RECT 84.285 116.605 84.575 116.650 ;
        RECT 86.805 116.605 87.095 116.650 ;
        RECT 93.255 116.790 93.545 116.835 ;
        RECT 95.080 116.790 95.400 116.850 ;
        RECT 93.255 116.650 95.400 116.790 ;
        RECT 93.255 116.605 93.545 116.650 ;
        RECT 95.080 116.590 95.400 116.650 ;
        RECT 28.840 116.250 29.160 116.510 ;
        RECT 29.760 116.250 30.080 116.510 ;
        RECT 73.935 116.450 74.225 116.495 ;
        RECT 80.820 116.450 81.140 116.510 ;
        RECT 82.215 116.450 82.505 116.495 ;
        RECT 86.340 116.450 86.660 116.510 ;
        RECT 73.935 116.310 86.660 116.450 ;
        RECT 73.935 116.265 74.225 116.310 ;
        RECT 80.820 116.250 81.140 116.310 ;
        RECT 82.215 116.265 82.505 116.310 ;
        RECT 86.340 116.250 86.660 116.310 ;
        RECT 89.560 116.450 89.880 116.510 ;
        RECT 94.635 116.450 94.925 116.495 ;
        RECT 89.560 116.310 94.925 116.450 ;
        RECT 97.010 116.450 97.150 116.990 ;
        RECT 110.720 116.990 114.680 117.130 ;
        RECT 110.720 116.945 111.010 116.990 ;
        RECT 112.290 116.945 112.580 116.990 ;
        RECT 114.390 116.945 114.680 116.990 ;
        RECT 106.135 116.790 106.425 116.835 ;
        RECT 108.420 116.790 108.740 116.850 ;
        RECT 114.950 116.835 115.090 117.330 ;
        RECT 123.600 117.270 123.920 117.530 ;
        RECT 128.660 117.470 128.980 117.530 ;
        RECT 124.150 117.330 128.980 117.470 ;
        RECT 123.155 117.130 123.445 117.175 ;
        RECT 124.150 117.130 124.290 117.330 ;
        RECT 128.660 117.270 128.980 117.330 ;
        RECT 136.480 117.270 136.800 117.530 ;
        RECT 123.155 116.990 124.290 117.130 ;
        RECT 123.155 116.945 123.445 116.990 ;
        RECT 124.980 116.930 125.300 117.190 ;
        RECT 136.020 117.130 136.340 117.190 ;
        RECT 125.530 116.990 136.340 117.130 ;
        RECT 100.690 116.650 108.740 116.790 ;
        RECT 100.690 116.510 100.830 116.650 ;
        RECT 106.135 116.605 106.425 116.650 ;
        RECT 108.420 116.590 108.740 116.650 ;
        RECT 110.285 116.790 110.575 116.835 ;
        RECT 112.805 116.790 113.095 116.835 ;
        RECT 113.995 116.790 114.285 116.835 ;
        RECT 110.285 116.650 114.285 116.790 ;
        RECT 110.285 116.605 110.575 116.650 ;
        RECT 112.805 116.605 113.095 116.650 ;
        RECT 113.995 116.605 114.285 116.650 ;
        RECT 114.875 116.790 115.165 116.835 ;
        RECT 122.220 116.790 122.540 116.850 ;
        RECT 124.520 116.790 124.840 116.850 ;
        RECT 125.530 116.790 125.670 116.990 ;
        RECT 136.020 116.930 136.340 116.990 ;
        RECT 114.875 116.650 125.670 116.790 ;
        RECT 114.875 116.605 115.165 116.650 ;
        RECT 122.220 116.590 122.540 116.650 ;
        RECT 124.520 116.590 124.840 116.650 ;
        RECT 126.360 116.590 126.680 116.850 ;
        RECT 139.700 116.590 140.020 116.850 ;
        RECT 144.300 116.790 144.620 116.850 ;
        RECT 142.090 116.650 144.620 116.790 ;
        RECT 97.395 116.450 97.685 116.495 ;
        RECT 98.775 116.450 99.065 116.495 ;
        RECT 97.010 116.310 99.065 116.450 ;
        RECT 89.560 116.250 89.880 116.310 ;
        RECT 94.635 116.265 94.925 116.310 ;
        RECT 97.395 116.265 97.685 116.310 ;
        RECT 98.775 116.265 99.065 116.310 ;
        RECT 100.600 116.250 100.920 116.510 ;
        RECT 101.060 116.250 101.380 116.510 ;
        RECT 104.740 116.450 105.060 116.510 ;
        RECT 105.215 116.450 105.505 116.495 ;
        RECT 104.740 116.310 105.505 116.450 ;
        RECT 104.740 116.250 105.060 116.310 ;
        RECT 105.215 116.265 105.505 116.310 ;
        RECT 105.675 116.450 105.965 116.495 ;
        RECT 107.960 116.450 108.280 116.510 ;
        RECT 105.675 116.310 108.280 116.450 ;
        RECT 105.675 116.265 105.965 116.310 ;
        RECT 107.960 116.250 108.280 116.310 ;
        RECT 121.315 116.450 121.605 116.495 ;
        RECT 131.420 116.450 131.740 116.510 ;
        RECT 134.180 116.450 134.500 116.510 ;
        RECT 121.315 116.310 134.500 116.450 ;
        RECT 121.315 116.265 121.605 116.310 ;
        RECT 131.420 116.250 131.740 116.310 ;
        RECT 134.180 116.250 134.500 116.310 ;
        RECT 137.400 116.450 137.720 116.510 ;
        RECT 141.540 116.495 141.860 116.510 ;
        RECT 142.090 116.495 142.230 116.650 ;
        RECT 144.300 116.590 144.620 116.650 ;
        RECT 138.335 116.450 138.625 116.495 ;
        RECT 141.530 116.450 141.860 116.495 ;
        RECT 137.400 116.310 138.625 116.450 ;
        RECT 141.345 116.310 141.860 116.450 ;
        RECT 137.400 116.250 137.720 116.310 ;
        RECT 138.335 116.265 138.625 116.310 ;
        RECT 141.530 116.265 141.860 116.310 ;
        RECT 142.015 116.265 142.305 116.495 ;
        RECT 141.540 116.250 141.860 116.265 ;
        RECT 71.175 116.110 71.465 116.155 ;
        RECT 75.270 116.110 75.560 116.155 ;
        RECT 76.220 116.110 76.540 116.170 ;
        RECT 71.175 115.970 74.150 116.110 ;
        RECT 71.175 115.925 71.465 115.970 ;
        RECT 74.010 115.830 74.150 115.970 ;
        RECT 75.270 115.970 76.540 116.110 ;
        RECT 75.270 115.925 75.560 115.970 ;
        RECT 76.220 115.910 76.540 115.970 ;
        RECT 83.550 116.110 83.840 116.155 ;
        RECT 84.500 116.110 84.820 116.170 ;
        RECT 101.150 116.110 101.290 116.250 ;
        RECT 83.550 115.970 84.820 116.110 ;
        RECT 83.550 115.925 83.840 115.970 ;
        RECT 84.500 115.910 84.820 115.970 ;
        RECT 87.350 115.970 101.290 116.110 ;
        RECT 110.260 116.110 110.580 116.170 ;
        RECT 113.540 116.110 113.830 116.155 ;
        RECT 110.260 115.970 113.830 116.110 ;
        RECT 28.840 115.770 29.160 115.830 ;
        RECT 29.315 115.770 29.605 115.815 ;
        RECT 28.840 115.630 29.605 115.770 ;
        RECT 28.840 115.570 29.160 115.630 ;
        RECT 29.315 115.585 29.605 115.630 ;
        RECT 73.460 115.570 73.780 115.830 ;
        RECT 73.920 115.570 74.240 115.830 ;
        RECT 79.900 115.770 80.220 115.830 ;
        RECT 80.835 115.770 81.125 115.815 ;
        RECT 79.900 115.630 81.125 115.770 ;
        RECT 79.900 115.570 80.220 115.630 ;
        RECT 80.835 115.585 81.125 115.630 ;
        RECT 84.960 115.770 85.280 115.830 ;
        RECT 87.350 115.770 87.490 115.970 ;
        RECT 110.260 115.910 110.580 115.970 ;
        RECT 113.540 115.925 113.830 115.970 ;
        RECT 138.795 116.110 139.085 116.155 ;
        RECT 142.090 116.110 142.230 116.265 ;
        RECT 142.460 116.250 142.780 116.510 ;
        RECT 143.380 116.450 143.700 116.510 ;
        RECT 143.185 116.310 143.700 116.450 ;
        RECT 143.380 116.250 143.700 116.310 ;
        RECT 143.855 116.265 144.145 116.495 ;
        RECT 138.795 115.970 142.230 116.110 ;
        RECT 138.795 115.925 139.085 115.970 ;
        RECT 84.960 115.630 87.490 115.770 ;
        RECT 84.960 115.570 85.280 115.630 ;
        RECT 89.100 115.570 89.420 115.830 ;
        RECT 90.020 115.770 90.340 115.830 ;
        RECT 92.335 115.770 92.625 115.815 ;
        RECT 90.020 115.630 92.625 115.770 ;
        RECT 90.020 115.570 90.340 115.630 ;
        RECT 92.335 115.585 92.625 115.630 ;
        RECT 92.795 115.770 93.085 115.815 ;
        RECT 93.700 115.770 94.020 115.830 ;
        RECT 92.795 115.630 94.020 115.770 ;
        RECT 92.795 115.585 93.085 115.630 ;
        RECT 93.700 115.570 94.020 115.630 ;
        RECT 103.360 115.570 103.680 115.830 ;
        RECT 107.975 115.770 108.265 115.815 ;
        RECT 108.880 115.770 109.200 115.830 ;
        RECT 111.180 115.770 111.500 115.830 ;
        RECT 107.975 115.630 111.500 115.770 ;
        RECT 107.975 115.585 108.265 115.630 ;
        RECT 108.880 115.570 109.200 115.630 ;
        RECT 111.180 115.570 111.500 115.630 ;
        RECT 124.060 115.570 124.380 115.830 ;
        RECT 140.620 115.570 140.940 115.830 ;
        RECT 141.080 115.770 141.400 115.830 ;
        RECT 143.930 115.770 144.070 116.265 ;
        RECT 141.080 115.630 144.070 115.770 ;
        RECT 141.080 115.570 141.400 115.630 ;
        RECT 17.270 114.950 146.990 115.430 ;
        RECT 32.060 114.750 32.380 114.810 ;
        RECT 33.915 114.750 34.205 114.795 ;
        RECT 20.190 114.610 34.205 114.750 ;
        RECT 20.190 114.115 20.330 114.610 ;
        RECT 32.060 114.550 32.380 114.610 ;
        RECT 33.915 114.565 34.205 114.610 ;
        RECT 73.000 114.750 73.320 114.810 ;
        RECT 78.535 114.750 78.825 114.795 ;
        RECT 73.000 114.610 78.825 114.750 ;
        RECT 73.000 114.550 73.320 114.610 ;
        RECT 78.535 114.565 78.825 114.610 ;
        RECT 79.900 114.750 80.220 114.810 ;
        RECT 85.895 114.750 86.185 114.795 ;
        RECT 97.380 114.750 97.700 114.810 ;
        RECT 79.900 114.610 84.730 114.750 ;
        RECT 79.900 114.550 80.220 114.610 ;
        RECT 27.460 114.410 27.780 114.470 ;
        RECT 23.410 114.270 27.780 114.410 ;
        RECT 20.115 113.885 20.405 114.115 ;
        RECT 23.410 113.775 23.550 114.270 ;
        RECT 27.460 114.210 27.780 114.270 ;
        RECT 72.510 114.410 72.800 114.455 ;
        RECT 73.460 114.410 73.780 114.470 ;
        RECT 72.510 114.270 73.780 114.410 ;
        RECT 72.510 114.225 72.800 114.270 ;
        RECT 73.460 114.210 73.780 114.270 ;
        RECT 80.360 114.210 80.680 114.470 ;
        RECT 83.580 114.410 83.900 114.470 ;
        RECT 84.590 114.455 84.730 114.610 ;
        RECT 85.895 114.610 97.700 114.750 ;
        RECT 85.895 114.565 86.185 114.610 ;
        RECT 97.380 114.550 97.700 114.610 ;
        RECT 101.060 114.550 101.380 114.810 ;
        RECT 101.520 114.750 101.840 114.810 ;
        RECT 112.575 114.750 112.865 114.795 ;
        RECT 124.980 114.750 125.300 114.810 ;
        RECT 129.595 114.750 129.885 114.795 ;
        RECT 101.520 114.610 110.950 114.750 ;
        RECT 101.520 114.550 101.840 114.610 ;
        RECT 84.055 114.410 84.345 114.455 ;
        RECT 80.910 114.270 83.350 114.410 ;
        RECT 24.240 113.870 24.560 114.130 ;
        RECT 28.350 114.070 28.640 114.115 ;
        RECT 30.680 114.070 31.000 114.130 ;
        RECT 28.350 113.930 31.000 114.070 ;
        RECT 28.350 113.885 28.640 113.930 ;
        RECT 30.680 113.870 31.000 113.930 ;
        RECT 66.560 114.070 66.880 114.130 ;
        RECT 71.175 114.070 71.465 114.115 ;
        RECT 66.560 113.930 71.465 114.070 ;
        RECT 66.560 113.870 66.880 113.930 ;
        RECT 71.175 113.885 71.465 113.930 ;
        RECT 23.335 113.545 23.625 113.775 ;
        RECT 23.780 113.530 24.100 113.790 ;
        RECT 27.000 113.530 27.320 113.790 ;
        RECT 80.910 113.775 81.050 114.270 ;
        RECT 83.210 114.115 83.350 114.270 ;
        RECT 83.580 114.270 84.345 114.410 ;
        RECT 83.580 114.210 83.900 114.270 ;
        RECT 84.055 114.225 84.345 114.270 ;
        RECT 84.515 114.225 84.805 114.455 ;
        RECT 94.620 114.410 94.940 114.470 ;
        RECT 107.960 114.410 108.280 114.470 ;
        RECT 110.810 114.455 110.950 114.610 ;
        RECT 112.575 114.610 124.750 114.750 ;
        RECT 112.575 114.565 112.865 114.610 ;
        RECT 110.735 114.410 111.025 114.455 ;
        RECT 114.860 114.410 115.180 114.470 ;
        RECT 86.890 114.270 102.670 114.410 ;
        RECT 86.890 114.130 87.030 114.270 ;
        RECT 94.620 114.210 94.940 114.270 ;
        RECT 84.960 114.115 85.280 114.130 ;
        RECT 82.675 113.885 82.965 114.115 ;
        RECT 83.140 113.885 83.430 114.115 ;
        RECT 84.960 114.070 85.290 114.115 ;
        RECT 84.960 113.930 85.475 114.070 ;
        RECT 84.960 113.885 85.290 113.930 ;
        RECT 27.895 113.730 28.185 113.775 ;
        RECT 29.085 113.730 29.375 113.775 ;
        RECT 31.605 113.730 31.895 113.775 ;
        RECT 27.895 113.590 31.895 113.730 ;
        RECT 27.895 113.545 28.185 113.590 ;
        RECT 29.085 113.545 29.375 113.590 ;
        RECT 31.605 113.545 31.895 113.590 ;
        RECT 72.055 113.730 72.345 113.775 ;
        RECT 73.245 113.730 73.535 113.775 ;
        RECT 75.765 113.730 76.055 113.775 ;
        RECT 80.835 113.730 81.125 113.775 ;
        RECT 72.055 113.590 76.055 113.730 ;
        RECT 72.055 113.545 72.345 113.590 ;
        RECT 73.245 113.545 73.535 113.590 ;
        RECT 75.765 113.545 76.055 113.590 ;
        RECT 78.150 113.590 81.125 113.730 ;
        RECT 27.500 113.390 27.790 113.435 ;
        RECT 29.600 113.390 29.890 113.435 ;
        RECT 31.170 113.390 31.460 113.435 ;
        RECT 27.500 113.250 31.460 113.390 ;
        RECT 27.500 113.205 27.790 113.250 ;
        RECT 29.600 113.205 29.890 113.250 ;
        RECT 31.170 113.205 31.460 113.250 ;
        RECT 71.660 113.390 71.950 113.435 ;
        RECT 73.760 113.390 74.050 113.435 ;
        RECT 75.330 113.390 75.620 113.435 ;
        RECT 71.660 113.250 75.620 113.390 ;
        RECT 71.660 113.205 71.950 113.250 ;
        RECT 73.760 113.205 74.050 113.250 ;
        RECT 75.330 113.205 75.620 113.250 ;
        RECT 15.960 113.050 16.280 113.110 ;
        RECT 19.195 113.050 19.485 113.095 ;
        RECT 15.220 112.910 19.485 113.050 ;
        RECT 15.960 112.850 16.280 112.910 ;
        RECT 19.195 112.865 19.485 112.910 ;
        RECT 25.620 113.050 25.940 113.110 ;
        RECT 26.095 113.050 26.385 113.095 ;
        RECT 25.620 112.910 26.385 113.050 ;
        RECT 25.620 112.850 25.940 112.910 ;
        RECT 26.095 112.865 26.385 112.910 ;
        RECT 77.600 113.050 77.920 113.110 ;
        RECT 78.150 113.095 78.290 113.590 ;
        RECT 80.835 113.545 81.125 113.590 ;
        RECT 81.755 113.545 82.045 113.775 ;
        RECT 82.750 113.730 82.890 113.885 ;
        RECT 84.960 113.870 85.280 113.885 ;
        RECT 86.800 113.870 87.120 114.130 ;
        RECT 88.180 114.115 88.500 114.130 ;
        RECT 88.150 114.070 88.500 114.115 ;
        RECT 87.985 113.930 88.500 114.070 ;
        RECT 88.150 113.885 88.500 113.930 ;
        RECT 88.180 113.870 88.500 113.885 ;
        RECT 95.540 113.870 95.860 114.130 ;
        RECT 97.380 113.870 97.700 114.130 ;
        RECT 101.520 113.870 101.840 114.130 ;
        RECT 102.530 114.115 102.670 114.270 ;
        RECT 107.960 114.270 110.030 114.410 ;
        RECT 107.960 114.210 108.280 114.270 ;
        RECT 102.455 113.885 102.745 114.115 ;
        RECT 102.900 114.070 103.220 114.130 ;
        RECT 103.735 114.070 104.025 114.115 ;
        RECT 102.900 113.930 104.025 114.070 ;
        RECT 102.900 113.870 103.220 113.930 ;
        RECT 103.735 113.885 104.025 113.930 ;
        RECT 105.200 114.070 105.520 114.130 ;
        RECT 109.890 114.115 110.030 114.270 ;
        RECT 110.735 114.270 115.180 114.410 ;
        RECT 110.735 114.225 111.025 114.270 ;
        RECT 114.860 114.210 115.180 114.270 ;
        RECT 123.570 114.410 123.860 114.455 ;
        RECT 124.060 114.410 124.380 114.470 ;
        RECT 123.570 114.270 124.380 114.410 ;
        RECT 124.610 114.410 124.750 114.610 ;
        RECT 124.980 114.610 129.885 114.750 ;
        RECT 124.980 114.550 125.300 114.610 ;
        RECT 129.595 114.565 129.885 114.610 ;
        RECT 131.435 114.750 131.725 114.795 ;
        RECT 137.400 114.750 137.720 114.810 ;
        RECT 131.435 114.610 137.720 114.750 ;
        RECT 131.435 114.565 131.725 114.610 ;
        RECT 137.400 114.550 137.720 114.610 ;
        RECT 139.700 114.750 140.020 114.810 ;
        RECT 145.220 114.750 145.540 114.810 ;
        RECT 139.700 114.610 145.540 114.750 ;
        RECT 139.700 114.550 140.020 114.610 ;
        RECT 145.220 114.550 145.540 114.610 ;
        RECT 129.120 114.410 129.440 114.470 ;
        RECT 124.610 114.270 129.440 114.410 ;
        RECT 123.570 114.225 123.860 114.270 ;
        RECT 124.060 114.210 124.380 114.270 ;
        RECT 129.120 114.210 129.440 114.270 ;
        RECT 131.895 114.410 132.185 114.455 ;
        RECT 143.380 114.410 143.700 114.470 ;
        RECT 131.895 114.270 143.700 114.410 ;
        RECT 131.895 114.225 132.185 114.270 ;
        RECT 105.200 113.930 109.110 114.070 ;
        RECT 105.200 113.870 105.520 113.930 ;
        RECT 86.340 113.730 86.660 113.790 ;
        RECT 82.750 113.590 86.660 113.730 ;
        RECT 81.830 113.390 81.970 113.545 ;
        RECT 86.340 113.530 86.660 113.590 ;
        RECT 87.695 113.730 87.985 113.775 ;
        RECT 88.885 113.730 89.175 113.775 ;
        RECT 91.405 113.730 91.695 113.775 ;
        RECT 87.695 113.590 91.695 113.730 ;
        RECT 87.695 113.545 87.985 113.590 ;
        RECT 88.885 113.545 89.175 113.590 ;
        RECT 91.405 113.545 91.695 113.590 ;
        RECT 103.335 113.730 103.625 113.775 ;
        RECT 104.525 113.730 104.815 113.775 ;
        RECT 107.045 113.730 107.335 113.775 ;
        RECT 103.335 113.590 107.335 113.730 ;
        RECT 108.970 113.730 109.110 113.930 ;
        RECT 109.815 113.885 110.105 114.115 ;
        RECT 111.180 113.870 111.500 114.130 ;
        RECT 111.655 113.885 111.945 114.115 ;
        RECT 111.730 113.730 111.870 113.885 ;
        RECT 116.700 113.730 117.020 113.790 ;
        RECT 108.970 113.590 117.020 113.730 ;
        RECT 103.335 113.545 103.625 113.590 ;
        RECT 104.525 113.545 104.815 113.590 ;
        RECT 107.045 113.545 107.335 113.590 ;
        RECT 116.700 113.530 117.020 113.590 ;
        RECT 122.220 113.530 122.540 113.790 ;
        RECT 123.115 113.730 123.405 113.775 ;
        RECT 124.305 113.730 124.595 113.775 ;
        RECT 126.825 113.730 127.115 113.775 ;
        RECT 123.115 113.590 127.115 113.730 ;
        RECT 123.115 113.545 123.405 113.590 ;
        RECT 124.305 113.545 124.595 113.590 ;
        RECT 126.825 113.545 127.115 113.590 ;
        RECT 86.800 113.390 87.120 113.450 ;
        RECT 81.830 113.250 87.120 113.390 ;
        RECT 86.800 113.190 87.120 113.250 ;
        RECT 87.300 113.390 87.590 113.435 ;
        RECT 89.400 113.390 89.690 113.435 ;
        RECT 90.970 113.390 91.260 113.435 ;
        RECT 100.600 113.390 100.920 113.450 ;
        RECT 87.300 113.250 91.260 113.390 ;
        RECT 87.300 113.205 87.590 113.250 ;
        RECT 89.400 113.205 89.690 113.250 ;
        RECT 90.970 113.205 91.260 113.250 ;
        RECT 93.330 113.250 100.920 113.390 ;
        RECT 78.075 113.050 78.365 113.095 ;
        RECT 77.600 112.910 78.365 113.050 ;
        RECT 77.600 112.850 77.920 112.910 ;
        RECT 78.075 112.865 78.365 112.910 ;
        RECT 78.980 113.050 79.300 113.110 ;
        RECT 93.330 113.050 93.470 113.250 ;
        RECT 100.600 113.190 100.920 113.250 ;
        RECT 102.940 113.390 103.230 113.435 ;
        RECT 105.040 113.390 105.330 113.435 ;
        RECT 106.610 113.390 106.900 113.435 ;
        RECT 102.940 113.250 106.900 113.390 ;
        RECT 102.940 113.205 103.230 113.250 ;
        RECT 105.040 113.205 105.330 113.250 ;
        RECT 106.610 113.205 106.900 113.250 ;
        RECT 108.420 113.390 108.740 113.450 ;
        RECT 122.720 113.390 123.010 113.435 ;
        RECT 124.820 113.390 125.110 113.435 ;
        RECT 126.390 113.390 126.680 113.435 ;
        RECT 108.420 113.250 122.220 113.390 ;
        RECT 108.420 113.190 108.740 113.250 ;
        RECT 78.980 112.910 93.470 113.050 ;
        RECT 78.980 112.850 79.300 112.910 ;
        RECT 93.700 112.850 94.020 113.110 ;
        RECT 95.080 113.050 95.400 113.110 ;
        RECT 98.300 113.050 98.620 113.110 ;
        RECT 95.080 112.910 98.620 113.050 ;
        RECT 95.080 112.850 95.400 112.910 ;
        RECT 98.300 112.850 98.620 112.910 ;
        RECT 107.960 113.050 108.280 113.110 ;
        RECT 109.355 113.050 109.645 113.095 ;
        RECT 107.960 112.910 109.645 113.050 ;
        RECT 122.080 113.050 122.220 113.250 ;
        RECT 122.720 113.250 126.680 113.390 ;
        RECT 122.720 113.205 123.010 113.250 ;
        RECT 124.820 113.205 125.110 113.250 ;
        RECT 126.390 113.205 126.680 113.250 ;
        RECT 129.135 113.390 129.425 113.435 ;
        RECT 131.970 113.390 132.110 114.225 ;
        RECT 143.380 114.210 143.700 114.270 ;
        RECT 137.400 114.070 137.720 114.130 ;
        RECT 141.555 114.070 141.845 114.115 ;
        RECT 137.400 113.930 141.845 114.070 ;
        RECT 137.400 113.870 137.720 113.930 ;
        RECT 141.555 113.885 141.845 113.930 ;
        RECT 143.855 114.070 144.145 114.115 ;
        RECT 144.300 114.070 144.620 114.130 ;
        RECT 143.855 113.930 144.620 114.070 ;
        RECT 143.855 113.885 144.145 113.930 ;
        RECT 144.300 113.870 144.620 113.930 ;
        RECT 132.800 113.530 133.120 113.790 ;
        RECT 137.860 113.530 138.180 113.790 ;
        RECT 138.795 113.730 139.085 113.775 ;
        RECT 139.700 113.730 140.020 113.790 ;
        RECT 138.795 113.590 140.020 113.730 ;
        RECT 138.795 113.545 139.085 113.590 ;
        RECT 139.700 113.530 140.020 113.590 ;
        RECT 142.000 113.530 142.320 113.790 ;
        RECT 142.475 113.545 142.765 113.775 ;
        RECT 139.240 113.390 139.560 113.450 ;
        RECT 142.550 113.390 142.690 113.545 ;
        RECT 129.135 113.250 132.110 113.390 ;
        RECT 132.430 113.250 142.690 113.390 ;
        RECT 129.135 113.205 129.425 113.250 ;
        RECT 132.430 113.050 132.570 113.250 ;
        RECT 139.240 113.190 139.560 113.250 ;
        RECT 144.760 113.190 145.080 113.450 ;
        RECT 122.080 112.910 132.570 113.050 ;
        RECT 133.260 113.050 133.580 113.110 ;
        RECT 135.575 113.050 135.865 113.095 ;
        RECT 133.260 112.910 135.865 113.050 ;
        RECT 107.960 112.850 108.280 112.910 ;
        RECT 109.355 112.865 109.645 112.910 ;
        RECT 133.260 112.850 133.580 112.910 ;
        RECT 135.575 112.865 135.865 112.910 ;
        RECT 136.480 113.050 136.800 113.110 ;
        RECT 139.715 113.050 140.005 113.095 ;
        RECT 136.480 112.910 140.005 113.050 ;
        RECT 136.480 112.850 136.800 112.910 ;
        RECT 139.715 112.865 140.005 112.910 ;
        RECT 17.270 112.230 146.990 112.710 ;
        RECT 19.195 112.030 19.485 112.075 ;
        RECT 20.100 112.030 20.420 112.090 ;
        RECT 24.240 112.030 24.560 112.090 ;
        RECT 19.195 111.890 24.560 112.030 ;
        RECT 19.195 111.845 19.485 111.890 ;
        RECT 20.100 111.830 20.420 111.890 ;
        RECT 24.240 111.830 24.560 111.890 ;
        RECT 30.680 111.830 31.000 112.090 ;
        RECT 84.500 111.830 84.820 112.090 ;
        RECT 86.340 112.030 86.660 112.090 ;
        RECT 88.655 112.030 88.945 112.075 ;
        RECT 86.340 111.890 88.945 112.030 ;
        RECT 86.340 111.830 86.660 111.890 ;
        RECT 88.655 111.845 88.945 111.890 ;
        RECT 102.900 111.830 103.220 112.090 ;
        RECT 110.260 111.830 110.580 112.090 ;
        RECT 124.520 112.030 124.840 112.090 ;
        RECT 132.800 112.030 133.120 112.090 ;
        RECT 114.490 111.890 133.120 112.030 ;
        RECT 21.940 111.690 22.230 111.735 ;
        RECT 23.510 111.690 23.800 111.735 ;
        RECT 25.610 111.690 25.900 111.735 ;
        RECT 21.940 111.550 25.900 111.690 ;
        RECT 21.940 111.505 22.230 111.550 ;
        RECT 23.510 111.505 23.800 111.550 ;
        RECT 25.610 111.505 25.900 111.550 ;
        RECT 63.840 111.690 64.130 111.735 ;
        RECT 65.940 111.690 66.230 111.735 ;
        RECT 67.510 111.690 67.800 111.735 ;
        RECT 63.840 111.550 67.800 111.690 ;
        RECT 63.840 111.505 64.130 111.550 ;
        RECT 65.940 111.505 66.230 111.550 ;
        RECT 67.510 111.505 67.800 111.550 ;
        RECT 68.400 111.690 68.720 111.750 ;
        RECT 73.920 111.690 74.240 111.750 ;
        RECT 68.400 111.550 82.430 111.690 ;
        RECT 68.400 111.490 68.720 111.550 ;
        RECT 73.920 111.490 74.240 111.550 ;
        RECT 21.505 111.350 21.795 111.395 ;
        RECT 24.025 111.350 24.315 111.395 ;
        RECT 25.215 111.350 25.505 111.395 ;
        RECT 21.505 111.210 25.505 111.350 ;
        RECT 21.505 111.165 21.795 111.210 ;
        RECT 24.025 111.165 24.315 111.210 ;
        RECT 25.215 111.165 25.505 111.210 ;
        RECT 27.460 111.350 27.780 111.410 ;
        RECT 33.455 111.350 33.745 111.395 ;
        RECT 27.460 111.210 33.745 111.350 ;
        RECT 27.460 111.150 27.780 111.210 ;
        RECT 33.455 111.165 33.745 111.210 ;
        RECT 64.235 111.350 64.525 111.395 ;
        RECT 65.425 111.350 65.715 111.395 ;
        RECT 67.945 111.350 68.235 111.395 ;
        RECT 64.235 111.210 68.235 111.350 ;
        RECT 64.235 111.165 64.525 111.210 ;
        RECT 65.425 111.165 65.715 111.210 ;
        RECT 67.945 111.165 68.235 111.210 ;
        RECT 71.160 111.350 71.480 111.410 ;
        RECT 73.475 111.350 73.765 111.395 ;
        RECT 78.980 111.350 79.300 111.410 ;
        RECT 82.290 111.395 82.430 111.550 ;
        RECT 84.040 111.490 84.360 111.750 ;
        RECT 103.360 111.490 103.680 111.750 ;
        RECT 109.800 111.490 110.120 111.750 ;
        RECT 71.160 111.210 79.300 111.350 ;
        RECT 71.160 111.150 71.480 111.210 ;
        RECT 73.475 111.165 73.765 111.210 ;
        RECT 78.980 111.150 79.300 111.210 ;
        RECT 82.215 111.350 82.505 111.395 ;
        RECT 96.460 111.350 96.780 111.410 ;
        RECT 82.215 111.210 96.780 111.350 ;
        RECT 82.215 111.165 82.505 111.210 ;
        RECT 96.460 111.150 96.780 111.210 ;
        RECT 98.300 111.350 98.620 111.410 ;
        RECT 101.060 111.350 101.380 111.410 ;
        RECT 113.955 111.350 114.245 111.395 ;
        RECT 114.490 111.350 114.630 111.890 ;
        RECT 124.520 111.830 124.840 111.890 ;
        RECT 132.800 111.830 133.120 111.890 ;
        RECT 117.660 111.690 117.950 111.735 ;
        RECT 119.760 111.690 120.050 111.735 ;
        RECT 121.330 111.690 121.620 111.735 ;
        RECT 117.660 111.550 121.620 111.690 ;
        RECT 117.660 111.505 117.950 111.550 ;
        RECT 119.760 111.505 120.050 111.550 ;
        RECT 121.330 111.505 121.620 111.550 ;
        RECT 132.355 111.690 132.645 111.735 ;
        RECT 133.260 111.690 133.580 111.750 ;
        RECT 132.355 111.550 133.580 111.690 ;
        RECT 132.355 111.505 132.645 111.550 ;
        RECT 133.260 111.490 133.580 111.550 ;
        RECT 136.520 111.690 136.810 111.735 ;
        RECT 138.620 111.690 138.910 111.735 ;
        RECT 140.190 111.690 140.480 111.735 ;
        RECT 136.520 111.550 140.480 111.690 ;
        RECT 136.520 111.505 136.810 111.550 ;
        RECT 138.620 111.505 138.910 111.550 ;
        RECT 140.190 111.505 140.480 111.550 ;
        RECT 98.300 111.210 114.630 111.350 ;
        RECT 118.055 111.350 118.345 111.395 ;
        RECT 119.245 111.350 119.535 111.395 ;
        RECT 121.765 111.350 122.055 111.395 ;
        RECT 118.055 111.210 122.055 111.350 ;
        RECT 98.300 111.150 98.620 111.210 ;
        RECT 101.060 111.150 101.380 111.210 ;
        RECT 113.955 111.165 114.245 111.210 ;
        RECT 118.055 111.165 118.345 111.210 ;
        RECT 119.245 111.165 119.535 111.210 ;
        RECT 121.765 111.165 122.055 111.210 ;
        RECT 126.360 111.350 126.680 111.410 ;
        RECT 130.515 111.350 130.805 111.395 ;
        RECT 126.360 111.210 130.805 111.350 ;
        RECT 126.360 111.150 126.680 111.210 ;
        RECT 130.515 111.165 130.805 111.210 ;
        RECT 136.020 111.150 136.340 111.410 ;
        RECT 136.915 111.350 137.205 111.395 ;
        RECT 138.105 111.350 138.395 111.395 ;
        RECT 140.625 111.350 140.915 111.395 ;
        RECT 136.915 111.210 140.915 111.350 ;
        RECT 136.915 111.165 137.205 111.210 ;
        RECT 138.105 111.165 138.395 111.210 ;
        RECT 140.625 111.165 140.915 111.210 ;
        RECT 24.815 111.010 25.105 111.055 ;
        RECT 25.620 111.010 25.940 111.070 ;
        RECT 24.815 110.870 25.940 111.010 ;
        RECT 24.815 110.825 25.105 110.870 ;
        RECT 25.620 110.810 25.940 110.870 ;
        RECT 26.095 111.010 26.385 111.055 ;
        RECT 27.000 111.010 27.320 111.070 ;
        RECT 26.095 110.870 27.320 111.010 ;
        RECT 26.095 110.825 26.385 110.870 ;
        RECT 27.000 110.810 27.320 110.870 ;
        RECT 32.060 111.010 32.380 111.070 ;
        RECT 32.535 111.010 32.825 111.055 ;
        RECT 32.060 110.870 32.825 111.010 ;
        RECT 32.060 110.810 32.380 110.870 ;
        RECT 32.535 110.825 32.825 110.870 ;
        RECT 61.500 111.010 61.820 111.070 ;
        RECT 63.355 111.010 63.645 111.055 ;
        RECT 66.560 111.010 66.880 111.070 ;
        RECT 72.540 111.010 72.860 111.070 ;
        RECT 78.060 111.010 78.380 111.070 ;
        RECT 61.500 110.870 66.880 111.010 ;
        RECT 72.345 110.870 78.380 111.010 ;
        RECT 61.500 110.810 61.820 110.870 ;
        RECT 63.355 110.825 63.645 110.870 ;
        RECT 66.560 110.810 66.880 110.870 ;
        RECT 72.540 110.810 72.860 110.870 ;
        RECT 78.060 110.810 78.380 110.870 ;
        RECT 89.560 110.810 89.880 111.070 ;
        RECT 91.415 111.010 91.705 111.055 ;
        RECT 93.700 111.010 94.020 111.070 ;
        RECT 91.415 110.870 94.020 111.010 ;
        RECT 91.415 110.825 91.705 110.870 ;
        RECT 93.700 110.810 94.020 110.870 ;
        RECT 105.215 111.010 105.505 111.055 ;
        RECT 107.975 111.010 108.265 111.055 ;
        RECT 109.340 111.010 109.660 111.070 ;
        RECT 105.215 110.870 109.660 111.010 ;
        RECT 105.215 110.825 105.505 110.870 ;
        RECT 107.975 110.825 108.265 110.870 ;
        RECT 109.340 110.810 109.660 110.870 ;
        RECT 114.400 111.010 114.720 111.070 ;
        RECT 114.875 111.010 115.165 111.055 ;
        RECT 114.400 110.870 115.165 111.010 ;
        RECT 114.400 110.810 114.720 110.870 ;
        RECT 114.875 110.825 115.165 110.870 ;
        RECT 117.175 111.010 117.465 111.055 ;
        RECT 122.220 111.010 122.540 111.070 ;
        RECT 142.460 111.010 142.780 111.070 ;
        RECT 143.855 111.010 144.145 111.055 ;
        RECT 117.175 110.870 122.540 111.010 ;
        RECT 117.175 110.825 117.465 110.870 ;
        RECT 122.220 110.810 122.540 110.870 ;
        RECT 129.670 110.870 142.780 111.010 ;
        RECT 64.720 110.715 65.040 110.730 ;
        RECT 64.690 110.485 65.040 110.715 ;
        RECT 73.015 110.670 73.305 110.715 ;
        RECT 64.720 110.470 65.040 110.485 ;
        RECT 70.330 110.530 73.305 110.670 ;
        RECT 70.330 110.390 70.470 110.530 ;
        RECT 73.015 110.485 73.305 110.530 ;
        RECT 89.100 110.670 89.420 110.730 ;
        RECT 90.035 110.670 90.325 110.715 ;
        RECT 89.100 110.530 90.325 110.670 ;
        RECT 89.100 110.470 89.420 110.530 ;
        RECT 90.035 110.485 90.325 110.530 ;
        RECT 90.480 110.670 90.800 110.730 ;
        RECT 97.380 110.670 97.700 110.730 ;
        RECT 118.540 110.715 118.860 110.730 ;
        RECT 90.480 110.530 97.700 110.670 ;
        RECT 30.680 110.330 31.000 110.390 ;
        RECT 32.995 110.330 33.285 110.375 ;
        RECT 30.680 110.190 33.285 110.330 ;
        RECT 30.680 110.130 31.000 110.190 ;
        RECT 32.995 110.145 33.285 110.190 ;
        RECT 70.240 110.130 70.560 110.390 ;
        RECT 70.700 110.130 71.020 110.390 ;
        RECT 90.110 110.330 90.250 110.485 ;
        RECT 90.480 110.470 90.800 110.530 ;
        RECT 97.380 110.470 97.700 110.530 ;
        RECT 114.490 110.530 118.310 110.670 ;
        RECT 114.490 110.390 114.630 110.530 ;
        RECT 91.860 110.330 92.180 110.390 ;
        RECT 90.110 110.190 92.180 110.330 ;
        RECT 91.860 110.130 92.180 110.190 ;
        RECT 114.400 110.130 114.720 110.390 ;
        RECT 116.715 110.330 117.005 110.375 ;
        RECT 117.620 110.330 117.940 110.390 ;
        RECT 116.715 110.190 117.940 110.330 ;
        RECT 118.170 110.330 118.310 110.530 ;
        RECT 118.510 110.485 118.860 110.715 ;
        RECT 118.540 110.470 118.860 110.485 ;
        RECT 124.075 110.330 124.365 110.375 ;
        RECT 129.670 110.330 129.810 110.870 ;
        RECT 142.460 110.810 142.780 110.870 ;
        RECT 143.010 110.870 144.145 111.010 ;
        RECT 137.260 110.670 137.550 110.715 ;
        RECT 132.890 110.530 137.550 110.670 ;
        RECT 132.890 110.375 133.030 110.530 ;
        RECT 137.260 110.485 137.550 110.530 ;
        RECT 118.170 110.190 129.810 110.330 ;
        RECT 116.715 110.145 117.005 110.190 ;
        RECT 117.620 110.130 117.940 110.190 ;
        RECT 124.075 110.145 124.365 110.190 ;
        RECT 132.815 110.145 133.105 110.375 ;
        RECT 137.860 110.330 138.180 110.390 ;
        RECT 143.010 110.375 143.150 110.870 ;
        RECT 143.855 110.825 144.145 110.870 ;
        RECT 142.935 110.330 143.225 110.375 ;
        RECT 137.860 110.190 143.225 110.330 ;
        RECT 137.860 110.130 138.180 110.190 ;
        RECT 142.935 110.145 143.225 110.190 ;
        RECT 144.760 110.130 145.080 110.390 ;
        RECT 17.270 109.510 146.990 109.990 ;
        RECT 18.260 109.310 18.580 109.370 ;
        RECT 19.195 109.310 19.485 109.355 ;
        RECT 18.260 109.170 19.485 109.310 ;
        RECT 18.260 109.110 18.580 109.170 ;
        RECT 19.195 109.125 19.485 109.170 ;
        RECT 30.680 109.110 31.000 109.370 ;
        RECT 64.275 109.310 64.565 109.355 ;
        RECT 64.720 109.310 65.040 109.370 ;
        RECT 64.275 109.170 65.040 109.310 ;
        RECT 64.275 109.125 64.565 109.170 ;
        RECT 64.720 109.110 65.040 109.170 ;
        RECT 93.700 109.310 94.020 109.370 ;
        RECT 118.080 109.310 118.400 109.370 ;
        RECT 93.700 109.170 118.400 109.310 ;
        RECT 93.700 109.110 94.020 109.170 ;
        RECT 118.080 109.110 118.400 109.170 ;
        RECT 118.540 109.110 118.860 109.370 ;
        RECT 136.035 109.125 136.325 109.355 ;
        RECT 142.000 109.310 142.320 109.370 ;
        RECT 143.395 109.310 143.685 109.355 ;
        RECT 142.000 109.170 143.685 109.310 ;
        RECT 30.235 108.970 30.525 109.015 ;
        RECT 25.480 108.830 30.525 108.970 ;
        RECT 20.100 108.430 20.420 108.690 ;
        RECT 21.940 108.630 22.260 108.690 ;
        RECT 25.480 108.630 25.620 108.830 ;
        RECT 30.235 108.785 30.525 108.830 ;
        RECT 66.575 108.970 66.865 109.015 ;
        RECT 67.020 108.970 67.340 109.030 ;
        RECT 68.400 108.970 68.720 109.030 ;
        RECT 66.575 108.830 68.720 108.970 ;
        RECT 66.575 108.785 66.865 108.830 ;
        RECT 67.020 108.770 67.340 108.830 ;
        RECT 68.400 108.770 68.720 108.830 ;
        RECT 107.055 108.970 107.345 109.015 ;
        RECT 109.340 108.970 109.660 109.030 ;
        RECT 112.560 108.970 112.880 109.030 ;
        RECT 116.255 108.970 116.545 109.015 ;
        RECT 107.055 108.830 116.545 108.970 ;
        RECT 136.110 108.970 136.250 109.125 ;
        RECT 142.000 109.110 142.320 109.170 ;
        RECT 143.395 109.125 143.685 109.170 ;
        RECT 137.720 108.970 138.010 109.015 ;
        RECT 136.110 108.830 138.010 108.970 ;
        RECT 107.055 108.785 107.345 108.830 ;
        RECT 109.340 108.770 109.660 108.830 ;
        RECT 112.560 108.770 112.880 108.830 ;
        RECT 116.255 108.785 116.545 108.830 ;
        RECT 137.720 108.785 138.010 108.830 ;
        RECT 21.110 108.490 25.620 108.630 ;
        RECT 26.655 108.630 26.945 108.675 ;
        RECT 26.655 108.490 28.610 108.630 ;
        RECT 21.110 107.995 21.250 108.490 ;
        RECT 21.940 108.430 22.260 108.490 ;
        RECT 26.655 108.445 26.945 108.490 ;
        RECT 23.345 108.290 23.635 108.335 ;
        RECT 25.865 108.290 26.155 108.335 ;
        RECT 27.055 108.290 27.345 108.335 ;
        RECT 23.345 108.150 27.345 108.290 ;
        RECT 23.345 108.105 23.635 108.150 ;
        RECT 25.865 108.105 26.155 108.150 ;
        RECT 27.055 108.105 27.345 108.150 ;
        RECT 27.935 108.105 28.225 108.335 ;
        RECT 21.035 107.765 21.325 107.995 ;
        RECT 23.780 107.950 24.070 107.995 ;
        RECT 25.350 107.950 25.640 107.995 ;
        RECT 27.450 107.950 27.740 107.995 ;
        RECT 23.780 107.810 27.740 107.950 ;
        RECT 23.780 107.765 24.070 107.810 ;
        RECT 25.350 107.765 25.640 107.810 ;
        RECT 27.450 107.765 27.740 107.810 ;
        RECT 27.000 107.610 27.320 107.670 ;
        RECT 28.010 107.610 28.150 108.105 ;
        RECT 28.470 107.995 28.610 108.490 ;
        RECT 28.840 108.290 29.160 108.350 ;
        RECT 31.155 108.290 31.445 108.335 ;
        RECT 28.840 108.150 31.445 108.290 ;
        RECT 28.840 108.090 29.160 108.150 ;
        RECT 31.155 108.105 31.445 108.150 ;
        RECT 71.620 108.290 71.940 108.350 ;
        RECT 103.820 108.290 104.140 108.350 ;
        RECT 113.940 108.290 114.260 108.350 ;
        RECT 71.620 108.150 104.140 108.290 ;
        RECT 71.620 108.090 71.940 108.150 ;
        RECT 103.820 108.090 104.140 108.150 ;
        RECT 104.370 108.150 114.260 108.290 ;
        RECT 116.330 108.290 116.470 108.785 ;
        RECT 116.700 108.630 117.020 108.690 ;
        RECT 132.340 108.630 132.660 108.690 ;
        RECT 135.560 108.630 135.880 108.690 ;
        RECT 116.700 108.490 135.880 108.630 ;
        RECT 116.700 108.430 117.020 108.490 ;
        RECT 132.340 108.430 132.660 108.490 ;
        RECT 135.560 108.430 135.880 108.490 ;
        RECT 136.020 108.630 136.340 108.690 ;
        RECT 136.495 108.630 136.785 108.675 ;
        RECT 136.020 108.490 136.785 108.630 ;
        RECT 136.020 108.430 136.340 108.490 ;
        RECT 136.495 108.445 136.785 108.490 ;
        RECT 143.380 108.630 143.700 108.690 ;
        RECT 143.855 108.630 144.145 108.675 ;
        RECT 143.380 108.490 144.145 108.630 ;
        RECT 143.380 108.430 143.700 108.490 ;
        RECT 143.855 108.445 144.145 108.490 ;
        RECT 116.330 108.150 118.310 108.290 ;
        RECT 28.395 107.765 28.685 107.995 ;
        RECT 65.195 107.950 65.485 107.995 ;
        RECT 70.700 107.950 71.020 108.010 ;
        RECT 65.195 107.810 71.020 107.950 ;
        RECT 65.195 107.765 65.485 107.810 ;
        RECT 70.700 107.750 71.020 107.810 ;
        RECT 78.060 107.950 78.380 108.010 ;
        RECT 86.340 107.950 86.660 108.010 ;
        RECT 104.370 107.950 104.510 108.150 ;
        RECT 113.940 108.090 114.260 108.150 ;
        RECT 78.060 107.810 104.510 107.950 ;
        RECT 78.060 107.750 78.380 107.810 ;
        RECT 86.340 107.750 86.660 107.810 ;
        RECT 108.880 107.750 109.200 108.010 ;
        RECT 117.620 107.750 117.940 108.010 ;
        RECT 118.170 107.950 118.310 108.150 ;
        RECT 133.720 108.090 134.040 108.350 ;
        RECT 137.375 108.290 137.665 108.335 ;
        RECT 138.565 108.290 138.855 108.335 ;
        RECT 141.085 108.290 141.375 108.335 ;
        RECT 137.375 108.150 141.375 108.290 ;
        RECT 137.375 108.105 137.665 108.150 ;
        RECT 138.565 108.105 138.855 108.150 ;
        RECT 141.085 108.105 141.375 108.150 ;
        RECT 130.960 107.950 131.280 108.010 ;
        RECT 118.170 107.810 131.280 107.950 ;
        RECT 130.960 107.750 131.280 107.810 ;
        RECT 135.575 107.950 135.865 107.995 ;
        RECT 136.480 107.950 136.800 108.010 ;
        RECT 135.575 107.810 136.800 107.950 ;
        RECT 135.575 107.765 135.865 107.810 ;
        RECT 136.480 107.750 136.800 107.810 ;
        RECT 136.980 107.950 137.270 107.995 ;
        RECT 139.080 107.950 139.370 107.995 ;
        RECT 140.650 107.950 140.940 107.995 ;
        RECT 136.980 107.810 140.940 107.950 ;
        RECT 136.980 107.765 137.270 107.810 ;
        RECT 139.080 107.765 139.370 107.810 ;
        RECT 140.650 107.765 140.940 107.810 ;
        RECT 27.000 107.470 28.150 107.610 ;
        RECT 79.440 107.610 79.760 107.670 ;
        RECT 83.120 107.610 83.440 107.670 ;
        RECT 89.560 107.610 89.880 107.670 ;
        RECT 94.620 107.610 94.940 107.670 ;
        RECT 79.440 107.470 94.940 107.610 ;
        RECT 27.000 107.410 27.320 107.470 ;
        RECT 79.440 107.410 79.760 107.470 ;
        RECT 83.120 107.410 83.440 107.470 ;
        RECT 89.560 107.410 89.880 107.470 ;
        RECT 94.620 107.410 94.940 107.470 ;
        RECT 109.340 107.410 109.660 107.670 ;
        RECT 111.640 107.610 111.960 107.670 ;
        RECT 129.580 107.610 129.900 107.670 ;
        RECT 111.640 107.470 129.900 107.610 ;
        RECT 111.640 107.410 111.960 107.470 ;
        RECT 129.580 107.410 129.900 107.470 ;
        RECT 144.760 107.410 145.080 107.670 ;
        RECT 17.270 106.790 146.990 107.270 ;
        RECT 24.700 106.590 25.020 106.650 ;
        RECT 27.935 106.590 28.225 106.635 ;
        RECT 24.700 106.450 28.225 106.590 ;
        RECT 24.700 106.390 25.020 106.450 ;
        RECT 27.935 106.405 28.225 106.450 ;
        RECT 29.775 106.405 30.065 106.635 ;
        RECT 30.695 106.590 30.985 106.635 ;
        RECT 31.140 106.590 31.460 106.650 ;
        RECT 30.695 106.450 31.460 106.590 ;
        RECT 30.695 106.405 30.985 106.450 ;
        RECT 21.940 106.250 22.230 106.295 ;
        RECT 23.510 106.250 23.800 106.295 ;
        RECT 25.610 106.250 25.900 106.295 ;
        RECT 21.940 106.110 25.900 106.250 ;
        RECT 29.850 106.250 29.990 106.405 ;
        RECT 31.140 106.390 31.460 106.450 ;
        RECT 35.755 106.590 36.045 106.635 ;
        RECT 74.395 106.590 74.685 106.635 ;
        RECT 94.160 106.590 94.480 106.650 ;
        RECT 114.400 106.590 114.720 106.650 ;
        RECT 35.755 106.450 36.430 106.590 ;
        RECT 35.755 106.405 36.045 106.450 ;
        RECT 35.280 106.250 35.600 106.310 ;
        RECT 29.850 106.110 35.600 106.250 ;
        RECT 21.940 106.065 22.230 106.110 ;
        RECT 23.510 106.065 23.800 106.110 ;
        RECT 25.610 106.065 25.900 106.110 ;
        RECT 35.280 106.050 35.600 106.110 ;
        RECT 21.505 105.910 21.795 105.955 ;
        RECT 24.025 105.910 24.315 105.955 ;
        RECT 25.215 105.910 25.505 105.955 ;
        RECT 34.835 105.910 35.125 105.955 ;
        RECT 21.505 105.770 25.505 105.910 ;
        RECT 21.505 105.725 21.795 105.770 ;
        RECT 24.025 105.725 24.315 105.770 ;
        RECT 25.215 105.725 25.505 105.770 ;
        RECT 28.930 105.770 35.125 105.910 ;
        RECT 26.095 105.570 26.385 105.615 ;
        RECT 27.000 105.570 27.320 105.630 ;
        RECT 26.095 105.430 27.320 105.570 ;
        RECT 26.095 105.385 26.385 105.430 ;
        RECT 27.000 105.370 27.320 105.430 ;
        RECT 27.920 105.570 28.240 105.630 ;
        RECT 28.930 105.615 29.070 105.770 ;
        RECT 28.855 105.570 29.145 105.615 ;
        RECT 27.920 105.430 29.145 105.570 ;
        RECT 27.920 105.370 28.240 105.430 ;
        RECT 28.855 105.385 29.145 105.430 ;
        RECT 29.760 105.370 30.080 105.630 ;
        RECT 31.690 105.615 31.830 105.770 ;
        RECT 34.835 105.725 35.125 105.770 ;
        RECT 31.615 105.385 31.905 105.615 ;
        RECT 32.520 105.570 32.840 105.630 ;
        RECT 32.995 105.570 33.285 105.615 ;
        RECT 32.520 105.430 33.285 105.570 ;
        RECT 32.520 105.370 32.840 105.430 ;
        RECT 32.995 105.385 33.285 105.430 ;
        RECT 33.915 105.385 34.205 105.615 ;
        RECT 24.870 105.230 25.160 105.275 ;
        RECT 25.620 105.230 25.940 105.290 ;
        RECT 24.870 105.090 25.940 105.230 ;
        RECT 24.870 105.045 25.160 105.090 ;
        RECT 25.620 105.030 25.940 105.090 ;
        RECT 31.140 105.230 31.460 105.290 ;
        RECT 33.990 105.230 34.130 105.385 ;
        RECT 34.360 105.370 34.680 105.630 ;
        RECT 35.280 105.570 35.600 105.630 ;
        RECT 35.755 105.570 36.045 105.615 ;
        RECT 35.280 105.430 36.045 105.570 ;
        RECT 35.280 105.370 35.600 105.430 ;
        RECT 35.755 105.385 36.045 105.430 ;
        RECT 36.290 105.230 36.430 106.450 ;
        RECT 74.395 106.450 94.480 106.590 ;
        RECT 74.395 106.405 74.685 106.450 ;
        RECT 94.160 106.390 94.480 106.450 ;
        RECT 99.770 106.450 114.720 106.590 ;
        RECT 63.815 106.250 64.105 106.295 ;
        RECT 69.320 106.250 69.640 106.310 ;
        RECT 63.815 106.110 69.640 106.250 ;
        RECT 63.815 106.065 64.105 106.110 ;
        RECT 69.320 106.050 69.640 106.110 ;
        RECT 80.835 106.250 81.125 106.295 ;
        RECT 84.055 106.250 84.345 106.295 ;
        RECT 99.770 106.250 99.910 106.450 ;
        RECT 114.400 106.390 114.720 106.450 ;
        RECT 117.635 106.590 117.925 106.635 ;
        RECT 119.460 106.590 119.780 106.650 ;
        RECT 117.635 106.450 119.780 106.590 ;
        RECT 117.635 106.405 117.925 106.450 ;
        RECT 119.460 106.390 119.780 106.450 ;
        RECT 122.080 106.450 144.070 106.590 ;
        RECT 111.640 106.250 111.960 106.310 ;
        RECT 80.835 106.110 84.345 106.250 ;
        RECT 80.835 106.065 81.125 106.110 ;
        RECT 84.055 106.065 84.345 106.110 ;
        RECT 92.410 106.110 99.910 106.250 ;
        RECT 101.610 106.110 111.960 106.250 ;
        RECT 61.040 105.910 61.360 105.970 ;
        RECT 61.975 105.910 62.265 105.955 ;
        RECT 67.020 105.910 67.340 105.970 ;
        RECT 61.040 105.770 67.340 105.910 ;
        RECT 61.040 105.710 61.360 105.770 ;
        RECT 61.975 105.725 62.265 105.770 ;
        RECT 67.020 105.710 67.340 105.770 ;
        RECT 70.715 105.910 71.005 105.955 ;
        RECT 71.160 105.910 71.480 105.970 ;
        RECT 74.380 105.910 74.700 105.970 ;
        RECT 83.580 105.910 83.900 105.970 ;
        RECT 70.715 105.770 71.480 105.910 ;
        RECT 70.715 105.725 71.005 105.770 ;
        RECT 71.160 105.710 71.480 105.770 ;
        RECT 72.630 105.770 83.900 105.910 ;
        RECT 68.400 105.570 68.720 105.630 ;
        RECT 72.630 105.615 72.770 105.770 ;
        RECT 74.380 105.710 74.700 105.770 ;
        RECT 83.580 105.710 83.900 105.770 ;
        RECT 87.275 105.910 87.565 105.955 ;
        RECT 87.720 105.910 88.040 105.970 ;
        RECT 87.275 105.770 88.040 105.910 ;
        RECT 87.275 105.725 87.565 105.770 ;
        RECT 87.720 105.710 88.040 105.770 ;
        RECT 71.635 105.570 71.925 105.615 ;
        RECT 68.400 105.430 71.925 105.570 ;
        RECT 68.400 105.370 68.720 105.430 ;
        RECT 71.635 105.385 71.925 105.430 ;
        RECT 72.555 105.385 72.845 105.615 ;
        RECT 73.475 105.385 73.765 105.615 ;
        RECT 78.995 105.570 79.285 105.615 ;
        RECT 85.880 105.570 86.200 105.630 ;
        RECT 78.995 105.430 86.200 105.570 ;
        RECT 78.995 105.385 79.285 105.430 ;
        RECT 31.140 105.090 36.430 105.230 ;
        RECT 69.335 105.230 69.625 105.275 ;
        RECT 72.080 105.230 72.400 105.290 ;
        RECT 69.335 105.090 72.400 105.230 ;
        RECT 31.140 105.030 31.460 105.090 ;
        RECT 69.335 105.045 69.625 105.090 ;
        RECT 72.080 105.030 72.400 105.090 ;
        RECT 73.000 105.030 73.320 105.290 ;
        RECT 73.550 105.230 73.690 105.385 ;
        RECT 85.880 105.370 86.200 105.430 ;
        RECT 86.340 105.370 86.660 105.630 ;
        RECT 90.480 105.370 90.800 105.630 ;
        RECT 91.235 105.570 91.525 105.615 ;
        RECT 92.410 105.570 92.550 106.110 ;
        RECT 101.610 105.955 101.750 106.110 ;
        RECT 111.640 106.050 111.960 106.110 ;
        RECT 114.860 106.250 115.180 106.310 ;
        RECT 117.160 106.250 117.480 106.310 ;
        RECT 114.860 106.110 117.480 106.250 ;
        RECT 114.860 106.050 115.180 106.110 ;
        RECT 101.535 105.725 101.825 105.955 ;
        RECT 103.360 105.910 103.680 105.970 ;
        RECT 104.755 105.910 105.045 105.955 ;
        RECT 105.660 105.910 105.980 105.970 ;
        RECT 103.360 105.770 105.980 105.910 ;
        RECT 103.360 105.710 103.680 105.770 ;
        RECT 104.755 105.725 105.045 105.770 ;
        RECT 105.660 105.710 105.980 105.770 ;
        RECT 108.420 105.910 108.740 105.970 ;
        RECT 111.195 105.910 111.485 105.955 ;
        RECT 108.420 105.770 111.485 105.910 ;
        RECT 108.420 105.710 108.740 105.770 ;
        RECT 111.195 105.725 111.485 105.770 ;
        RECT 113.570 105.770 115.090 105.910 ;
        RECT 91.235 105.430 92.550 105.570 ;
        RECT 92.780 105.615 93.100 105.630 ;
        RECT 92.780 105.570 93.110 105.615 ;
        RECT 96.000 105.570 96.320 105.630 ;
        RECT 100.155 105.570 100.445 105.615 ;
        RECT 92.780 105.430 93.295 105.570 ;
        RECT 96.000 105.430 100.445 105.570 ;
        RECT 91.235 105.385 91.525 105.430 ;
        RECT 92.780 105.385 93.110 105.430 ;
        RECT 92.780 105.370 93.100 105.385 ;
        RECT 96.000 105.370 96.320 105.430 ;
        RECT 100.155 105.385 100.445 105.430 ;
        RECT 110.735 105.570 111.025 105.615 ;
        RECT 113.570 105.570 113.710 105.770 ;
        RECT 114.950 105.630 115.090 105.770 ;
        RECT 110.735 105.430 113.710 105.570 ;
        RECT 110.735 105.385 111.025 105.430 ;
        RECT 114.415 105.385 114.705 105.615 ;
        RECT 114.860 105.570 115.180 105.630 ;
        RECT 115.870 105.615 116.010 106.110 ;
        RECT 117.160 106.050 117.480 106.110 ;
        RECT 118.080 105.910 118.400 105.970 ;
        RECT 122.080 105.910 122.220 106.450 ;
        RECT 128.215 106.250 128.505 106.295 ;
        RECT 130.500 106.250 130.820 106.310 ;
        RECT 128.215 106.110 130.820 106.250 ;
        RECT 128.215 106.065 128.505 106.110 ;
        RECT 130.500 106.050 130.820 106.110 ;
        RECT 130.960 106.050 131.280 106.310 ;
        RECT 135.575 106.250 135.865 106.295 ;
        RECT 136.480 106.250 136.800 106.310 ;
        RECT 135.575 106.110 136.800 106.250 ;
        RECT 135.575 106.065 135.865 106.110 ;
        RECT 136.480 106.050 136.800 106.110 ;
        RECT 118.080 105.770 122.220 105.910 ;
        RECT 126.360 105.910 126.680 105.970 ;
        RECT 133.720 105.910 134.040 105.970 ;
        RECT 126.360 105.770 134.040 105.910 ;
        RECT 118.080 105.710 118.400 105.770 ;
        RECT 126.360 105.710 126.680 105.770 ;
        RECT 133.720 105.710 134.040 105.770 ;
        RECT 136.035 105.910 136.325 105.955 ;
        RECT 136.940 105.910 137.260 105.970 ;
        RECT 136.035 105.770 137.260 105.910 ;
        RECT 136.035 105.725 136.325 105.770 ;
        RECT 136.940 105.710 137.260 105.770 ;
        RECT 116.700 105.615 117.020 105.630 ;
        RECT 114.860 105.430 115.375 105.570 ;
        RECT 75.300 105.230 75.620 105.290 ;
        RECT 84.960 105.230 85.280 105.290 ;
        RECT 86.430 105.230 86.570 105.370 ;
        RECT 73.550 105.090 85.280 105.230 ;
        RECT 75.300 105.030 75.620 105.090 ;
        RECT 84.960 105.030 85.280 105.090 ;
        RECT 85.970 105.090 86.570 105.230 ;
        RECT 90.020 105.230 90.340 105.290 ;
        RECT 91.875 105.230 92.165 105.275 ;
        RECT 90.020 105.090 92.165 105.230 ;
        RECT 19.180 104.690 19.500 104.950 ;
        RECT 33.900 104.890 34.220 104.950 ;
        RECT 35.740 104.890 36.060 104.950 ;
        RECT 36.675 104.890 36.965 104.935 ;
        RECT 33.900 104.750 36.965 104.890 ;
        RECT 33.900 104.690 34.220 104.750 ;
        RECT 35.740 104.690 36.060 104.750 ;
        RECT 36.675 104.705 36.965 104.750 ;
        RECT 64.260 104.690 64.580 104.950 ;
        RECT 67.020 104.890 67.340 104.950 ;
        RECT 67.495 104.890 67.785 104.935 ;
        RECT 67.020 104.750 67.785 104.890 ;
        RECT 67.020 104.690 67.340 104.750 ;
        RECT 67.495 104.705 67.785 104.750 ;
        RECT 68.860 104.890 69.180 104.950 ;
        RECT 69.795 104.890 70.085 104.935 ;
        RECT 68.860 104.750 70.085 104.890 ;
        RECT 68.860 104.690 69.180 104.750 ;
        RECT 69.795 104.705 70.085 104.750 ;
        RECT 81.295 104.890 81.585 104.935 ;
        RECT 81.740 104.890 82.060 104.950 ;
        RECT 85.970 104.935 86.110 105.090 ;
        RECT 90.020 105.030 90.340 105.090 ;
        RECT 91.875 105.045 92.165 105.090 ;
        RECT 92.335 105.045 92.625 105.275 ;
        RECT 99.680 105.230 100.000 105.290 ;
        RECT 93.790 105.090 100.000 105.230 ;
        RECT 81.295 104.750 82.060 104.890 ;
        RECT 81.295 104.705 81.585 104.750 ;
        RECT 81.740 104.690 82.060 104.750 ;
        RECT 85.895 104.705 86.185 104.935 ;
        RECT 86.355 104.890 86.645 104.935 ;
        RECT 87.260 104.890 87.580 104.950 ;
        RECT 92.410 104.890 92.550 105.045 ;
        RECT 93.790 104.935 93.930 105.090 ;
        RECT 99.680 105.030 100.000 105.090 ;
        RECT 103.820 105.230 104.140 105.290 ;
        RECT 113.020 105.230 113.340 105.290 ;
        RECT 103.820 105.090 113.340 105.230 ;
        RECT 103.820 105.030 104.140 105.090 ;
        RECT 113.020 105.030 113.340 105.090 ;
        RECT 86.355 104.750 92.550 104.890 ;
        RECT 86.355 104.705 86.645 104.750 ;
        RECT 87.260 104.690 87.580 104.750 ;
        RECT 93.715 104.705 94.005 104.935 ;
        RECT 96.460 104.890 96.780 104.950 ;
        RECT 99.220 104.890 99.540 104.950 ;
        RECT 96.460 104.750 99.540 104.890 ;
        RECT 96.460 104.690 96.780 104.750 ;
        RECT 99.220 104.690 99.540 104.750 ;
        RECT 101.980 104.690 102.300 104.950 ;
        RECT 104.280 104.690 104.600 104.950 ;
        RECT 108.420 104.690 108.740 104.950 ;
        RECT 110.260 104.690 110.580 104.950 ;
        RECT 114.490 104.890 114.630 105.385 ;
        RECT 114.860 105.370 115.180 105.430 ;
        RECT 115.795 105.385 116.085 105.615 ;
        RECT 116.700 105.570 117.030 105.615 ;
        RECT 130.515 105.570 130.805 105.615 ;
        RECT 131.420 105.570 131.740 105.630 ;
        RECT 131.895 105.570 132.185 105.615 ;
        RECT 116.700 105.430 117.215 105.570 ;
        RECT 130.515 105.430 132.185 105.570 ;
        RECT 116.700 105.385 117.030 105.430 ;
        RECT 130.515 105.385 130.805 105.430 ;
        RECT 116.700 105.370 117.020 105.385 ;
        RECT 131.420 105.370 131.740 105.430 ;
        RECT 131.895 105.385 132.185 105.430 ;
        RECT 135.560 105.570 135.880 105.630 ;
        RECT 137.415 105.570 137.705 105.615 ;
        RECT 135.560 105.430 137.705 105.570 ;
        RECT 135.560 105.370 135.880 105.430 ;
        RECT 137.415 105.385 137.705 105.430 ;
        RECT 137.860 105.370 138.180 105.630 ;
        RECT 139.255 105.570 139.545 105.615 ;
        RECT 142.000 105.570 142.320 105.630 ;
        RECT 143.930 105.615 144.070 106.450 ;
        RECT 139.255 105.430 142.320 105.570 ;
        RECT 139.255 105.385 139.545 105.430 ;
        RECT 142.000 105.370 142.320 105.430 ;
        RECT 143.855 105.385 144.145 105.615 ;
        RECT 116.255 105.045 116.545 105.275 ;
        RECT 115.320 104.890 115.640 104.950 ;
        RECT 114.490 104.750 115.640 104.890 ;
        RECT 116.330 104.890 116.470 105.045 ;
        RECT 129.580 105.030 129.900 105.290 ;
        RECT 138.320 105.030 138.640 105.290 ;
        RECT 147.060 105.230 147.380 105.290 ;
        RECT 143.010 105.090 147.380 105.230 ;
        RECT 116.700 104.890 117.020 104.950 ;
        RECT 116.330 104.750 117.020 104.890 ;
        RECT 115.320 104.690 115.640 104.750 ;
        RECT 116.700 104.690 117.020 104.750 ;
        RECT 128.660 104.690 128.980 104.950 ;
        RECT 136.495 104.890 136.785 104.935 ;
        RECT 141.080 104.890 141.400 104.950 ;
        RECT 143.010 104.935 143.150 105.090 ;
        RECT 147.060 105.030 147.380 105.090 ;
        RECT 136.495 104.750 141.400 104.890 ;
        RECT 136.495 104.705 136.785 104.750 ;
        RECT 141.080 104.690 141.400 104.750 ;
        RECT 142.935 104.705 143.225 104.935 ;
        RECT 144.775 104.890 145.065 104.935 ;
        RECT 150.280 104.890 150.600 104.950 ;
        RECT 144.775 104.750 150.600 104.890 ;
        RECT 144.775 104.705 145.065 104.750 ;
        RECT 150.280 104.690 150.600 104.750 ;
        RECT 17.270 104.070 146.990 104.550 ;
        RECT 147.590 104.220 147.910 104.280 ;
        RECT 147.310 104.080 147.910 104.220 ;
        RECT 25.620 103.870 25.940 103.930 ;
        RECT 26.095 103.870 26.385 103.915 ;
        RECT 25.620 103.730 26.385 103.870 ;
        RECT 25.620 103.670 25.940 103.730 ;
        RECT 26.095 103.685 26.385 103.730 ;
        RECT 68.415 103.685 68.705 103.915 ;
        RECT 24.255 103.530 24.545 103.575 ;
        RECT 20.190 103.390 24.545 103.530 ;
        RECT 19.180 103.190 19.500 103.250 ;
        RECT 20.190 103.235 20.330 103.390 ;
        RECT 24.255 103.345 24.545 103.390 ;
        RECT 28.840 103.330 29.160 103.590 ;
        RECT 35.280 103.530 35.600 103.590 ;
        RECT 33.070 103.390 35.600 103.530 ;
        RECT 20.115 103.190 20.405 103.235 ;
        RECT 19.180 103.050 20.405 103.190 ;
        RECT 19.180 102.990 19.500 103.050 ;
        RECT 20.115 103.005 20.405 103.050 ;
        RECT 21.940 102.990 22.260 103.250 ;
        RECT 23.780 102.990 24.100 103.250 ;
        RECT 25.620 103.190 25.940 103.250 ;
        RECT 28.395 103.190 28.685 103.235 ;
        RECT 25.620 103.050 28.685 103.190 ;
        RECT 28.930 103.190 29.070 103.330 ;
        RECT 31.140 103.190 31.460 103.250 ;
        RECT 28.930 103.050 31.460 103.190 ;
        RECT 25.620 102.990 25.940 103.050 ;
        RECT 28.395 103.005 28.685 103.050 ;
        RECT 31.140 102.990 31.460 103.050 ;
        RECT 32.060 103.190 32.380 103.250 ;
        RECT 33.070 103.190 33.210 103.390 ;
        RECT 35.280 103.330 35.600 103.390 ;
        RECT 35.755 103.530 36.045 103.575 ;
        RECT 36.660 103.530 36.980 103.590 ;
        RECT 61.040 103.530 61.360 103.590 ;
        RECT 62.850 103.530 63.140 103.575 ;
        RECT 64.260 103.530 64.580 103.590 ;
        RECT 35.755 103.390 41.950 103.530 ;
        RECT 35.755 103.345 36.045 103.390 ;
        RECT 36.660 103.330 36.980 103.390 ;
        RECT 32.060 103.050 33.210 103.190 ;
        RECT 32.060 102.990 32.380 103.050 ;
        RECT 33.440 102.990 33.760 103.250 ;
        RECT 37.595 103.190 37.885 103.235 ;
        RECT 38.500 103.190 38.820 103.250 ;
        RECT 37.595 103.050 38.820 103.190 ;
        RECT 37.595 103.005 37.885 103.050 ;
        RECT 38.500 102.990 38.820 103.050 ;
        RECT 38.975 103.190 39.265 103.235 ;
        RECT 39.510 103.190 39.650 103.390 ;
        RECT 41.810 103.250 41.950 103.390 ;
        RECT 61.040 103.390 62.650 103.530 ;
        RECT 61.040 103.330 61.360 103.390 ;
        RECT 38.975 103.050 39.650 103.190 ;
        RECT 39.880 103.190 40.200 103.250 ;
        RECT 40.355 103.190 40.645 103.235 ;
        RECT 39.880 103.050 40.645 103.190 ;
        RECT 38.975 103.005 39.265 103.050 ;
        RECT 39.880 102.990 40.200 103.050 ;
        RECT 40.355 103.005 40.645 103.050 ;
        RECT 41.260 102.990 41.580 103.250 ;
        RECT 41.720 102.990 42.040 103.250 ;
        RECT 61.500 102.990 61.820 103.250 ;
        RECT 62.510 103.190 62.650 103.390 ;
        RECT 62.850 103.390 64.580 103.530 ;
        RECT 68.490 103.530 68.630 103.685 ;
        RECT 69.320 103.670 69.640 103.930 ;
        RECT 70.700 103.870 71.020 103.930 ;
        RECT 71.175 103.870 71.465 103.915 ;
        RECT 70.700 103.730 71.465 103.870 ;
        RECT 70.700 103.670 71.020 103.730 ;
        RECT 71.175 103.685 71.465 103.730 ;
        RECT 71.635 103.870 71.925 103.915 ;
        RECT 73.000 103.870 73.320 103.930 ;
        RECT 71.635 103.730 73.320 103.870 ;
        RECT 71.635 103.685 71.925 103.730 ;
        RECT 71.710 103.530 71.850 103.685 ;
        RECT 73.000 103.670 73.320 103.730 ;
        RECT 73.920 103.870 74.240 103.930 ;
        RECT 87.720 103.870 88.040 103.930 ;
        RECT 73.920 103.730 88.040 103.870 ;
        RECT 73.920 103.670 74.240 103.730 ;
        RECT 87.720 103.670 88.040 103.730 ;
        RECT 89.560 103.670 89.880 103.930 ;
        RECT 90.020 103.670 90.340 103.930 ;
        RECT 92.780 103.870 93.100 103.930 ;
        RECT 103.360 103.870 103.680 103.930 ;
        RECT 92.780 103.730 103.680 103.870 ;
        RECT 92.780 103.670 93.100 103.730 ;
        RECT 103.360 103.670 103.680 103.730 ;
        RECT 103.820 103.870 104.140 103.930 ;
        RECT 104.295 103.870 104.585 103.915 ;
        RECT 103.820 103.730 104.585 103.870 ;
        RECT 103.820 103.670 104.140 103.730 ;
        RECT 104.295 103.685 104.585 103.730 ;
        RECT 108.880 103.870 109.200 103.930 ;
        RECT 114.415 103.870 114.705 103.915 ;
        RECT 117.620 103.870 117.940 103.930 ;
        RECT 122.695 103.870 122.985 103.915 ;
        RECT 126.820 103.870 127.140 103.930 ;
        RECT 136.035 103.870 136.325 103.915 ;
        RECT 136.480 103.870 136.800 103.930 ;
        RECT 108.880 103.730 114.705 103.870 ;
        RECT 108.880 103.670 109.200 103.730 ;
        RECT 114.415 103.685 114.705 103.730 ;
        RECT 116.330 103.730 127.140 103.870 ;
        RECT 68.490 103.390 71.850 103.530 ;
        RECT 72.080 103.530 72.400 103.590 ;
        RECT 79.440 103.530 79.760 103.590 ;
        RECT 72.080 103.390 79.760 103.530 ;
        RECT 62.850 103.345 63.140 103.390 ;
        RECT 64.260 103.330 64.580 103.390 ;
        RECT 72.080 103.330 72.400 103.390 ;
        RECT 79.440 103.330 79.760 103.390 ;
        RECT 85.880 103.530 86.200 103.590 ;
        RECT 108.390 103.530 108.680 103.575 ;
        RECT 109.340 103.530 109.660 103.590 ;
        RECT 85.880 103.390 91.170 103.530 ;
        RECT 85.880 103.330 86.200 103.390 ;
        RECT 64.720 103.190 65.040 103.250 ;
        RECT 62.510 103.050 65.040 103.190 ;
        RECT 64.720 102.990 65.040 103.050 ;
        RECT 73.460 102.990 73.780 103.250 ;
        RECT 78.060 102.990 78.380 103.250 ;
        RECT 80.375 103.190 80.665 103.235 ;
        RECT 80.820 103.190 81.140 103.250 ;
        RECT 81.740 103.235 82.060 103.250 ;
        RECT 81.710 103.190 82.060 103.235 ;
        RECT 80.375 103.050 81.140 103.190 ;
        RECT 81.545 103.050 82.060 103.190 ;
        RECT 91.030 103.190 91.170 103.390 ;
        RECT 103.910 103.390 104.970 103.530 ;
        RECT 91.875 103.190 92.165 103.235 ;
        RECT 93.700 103.190 94.020 103.250 ;
        RECT 96.375 103.190 96.665 103.235 ;
        RECT 91.030 103.050 94.020 103.190 ;
        RECT 80.375 103.005 80.665 103.050 ;
        RECT 80.820 102.990 81.140 103.050 ;
        RECT 81.710 103.005 82.060 103.050 ;
        RECT 91.875 103.005 92.165 103.050 ;
        RECT 81.740 102.990 82.060 103.005 ;
        RECT 93.700 102.990 94.020 103.050 ;
        RECT 94.250 103.050 96.665 103.190 ;
        RECT 23.335 102.665 23.625 102.895 ;
        RECT 23.870 102.850 24.010 102.990 ;
        RECT 28.855 102.850 29.145 102.895 ;
        RECT 23.870 102.710 29.145 102.850 ;
        RECT 28.855 102.665 29.145 102.710 ;
        RECT 16.880 102.510 17.200 102.570 ;
        RECT 21.035 102.510 21.325 102.555 ;
        RECT 16.880 102.370 21.325 102.510 ;
        RECT 23.410 102.510 23.550 102.665 ;
        RECT 28.380 102.510 28.700 102.570 ;
        RECT 23.410 102.370 28.700 102.510 ;
        RECT 28.930 102.510 29.070 102.665 ;
        RECT 29.300 102.650 29.620 102.910 ;
        RECT 31.615 102.850 31.905 102.895 ;
        RECT 34.375 102.850 34.665 102.895 ;
        RECT 35.280 102.850 35.600 102.910 ;
        RECT 31.615 102.710 34.130 102.850 ;
        RECT 31.615 102.665 31.905 102.710 ;
        RECT 32.535 102.510 32.825 102.555 ;
        RECT 28.930 102.370 32.825 102.510 ;
        RECT 33.990 102.510 34.130 102.710 ;
        RECT 34.375 102.710 35.600 102.850 ;
        RECT 34.375 102.665 34.665 102.710 ;
        RECT 35.280 102.650 35.600 102.710 ;
        RECT 38.055 102.850 38.345 102.895 ;
        RECT 40.800 102.850 41.120 102.910 ;
        RECT 38.055 102.710 41.120 102.850 ;
        RECT 38.055 102.665 38.345 102.710 ;
        RECT 40.800 102.650 41.120 102.710 ;
        RECT 62.395 102.850 62.685 102.895 ;
        RECT 63.585 102.850 63.875 102.895 ;
        RECT 66.105 102.850 66.395 102.895 ;
        RECT 62.395 102.710 66.395 102.850 ;
        RECT 62.395 102.665 62.685 102.710 ;
        RECT 63.585 102.665 63.875 102.710 ;
        RECT 66.105 102.665 66.395 102.710 ;
        RECT 71.620 102.850 71.940 102.910 ;
        RECT 72.095 102.850 72.385 102.895 ;
        RECT 71.620 102.710 72.385 102.850 ;
        RECT 71.620 102.650 71.940 102.710 ;
        RECT 72.095 102.665 72.385 102.710 ;
        RECT 78.535 102.665 78.825 102.895 ;
        RECT 79.455 102.665 79.745 102.895 ;
        RECT 81.255 102.850 81.545 102.895 ;
        RECT 82.445 102.850 82.735 102.895 ;
        RECT 84.965 102.850 85.255 102.895 ;
        RECT 90.495 102.850 90.785 102.895 ;
        RECT 92.780 102.850 93.100 102.910 ;
        RECT 94.250 102.895 94.390 103.050 ;
        RECT 96.375 103.005 96.665 103.050 ;
        RECT 101.060 103.190 101.380 103.250 ;
        RECT 103.910 103.190 104.050 103.390 ;
        RECT 101.060 103.050 104.050 103.190 ;
        RECT 104.830 103.190 104.970 103.390 ;
        RECT 108.390 103.390 109.660 103.530 ;
        RECT 108.390 103.345 108.680 103.390 ;
        RECT 109.340 103.330 109.660 103.390 ;
        RECT 110.260 103.530 110.580 103.590 ;
        RECT 116.330 103.575 116.470 103.730 ;
        RECT 117.620 103.670 117.940 103.730 ;
        RECT 122.695 103.685 122.985 103.730 ;
        RECT 126.820 103.670 127.140 103.730 ;
        RECT 127.370 103.730 135.790 103.870 ;
        RECT 116.255 103.530 116.545 103.575 ;
        RECT 110.260 103.390 116.545 103.530 ;
        RECT 110.260 103.330 110.580 103.390 ;
        RECT 116.255 103.345 116.545 103.390 ;
        RECT 117.160 103.530 117.480 103.590 ;
        RECT 127.370 103.530 127.510 103.730 ;
        RECT 117.160 103.390 127.510 103.530 ;
        RECT 127.710 103.530 128.000 103.575 ;
        RECT 128.660 103.530 128.980 103.590 ;
        RECT 127.710 103.390 128.980 103.530 ;
        RECT 117.160 103.330 117.480 103.390 ;
        RECT 127.710 103.345 128.000 103.390 ;
        RECT 128.660 103.330 128.980 103.390 ;
        RECT 130.960 103.530 131.280 103.590 ;
        RECT 134.195 103.530 134.485 103.575 ;
        RECT 130.960 103.390 134.485 103.530 ;
        RECT 135.650 103.530 135.790 103.730 ;
        RECT 136.035 103.730 136.800 103.870 ;
        RECT 136.035 103.685 136.325 103.730 ;
        RECT 136.480 103.670 136.800 103.730 ;
        RECT 137.400 103.870 137.720 103.930 ;
        RECT 137.875 103.870 138.165 103.915 ;
        RECT 137.400 103.730 138.165 103.870 ;
        RECT 137.400 103.670 137.720 103.730 ;
        RECT 137.875 103.685 138.165 103.730 ;
        RECT 138.320 103.670 138.640 103.930 ;
        RECT 138.410 103.530 138.550 103.670 ;
        RECT 135.650 103.390 141.310 103.530 ;
        RECT 130.960 103.330 131.280 103.390 ;
        RECT 134.195 103.345 134.485 103.390 ;
        RECT 105.660 103.190 105.980 103.250 ;
        RECT 116.700 103.190 117.020 103.250 ;
        RECT 120.840 103.190 121.160 103.250 ;
        RECT 141.170 103.235 141.310 103.390 ;
        RECT 138.335 103.190 138.625 103.235 ;
        RECT 104.830 103.050 105.430 103.190 ;
        RECT 101.060 102.990 101.380 103.050 ;
        RECT 81.255 102.710 85.255 102.850 ;
        RECT 81.255 102.665 81.545 102.710 ;
        RECT 82.445 102.665 82.735 102.710 ;
        RECT 84.965 102.665 85.255 102.710 ;
        RECT 86.890 102.710 93.100 102.850 ;
        RECT 38.515 102.510 38.805 102.555 ;
        RECT 43.560 102.510 43.880 102.570 ;
        RECT 33.990 102.370 38.270 102.510 ;
        RECT 16.880 102.310 17.200 102.370 ;
        RECT 21.035 102.325 21.325 102.370 ;
        RECT 28.380 102.310 28.700 102.370 ;
        RECT 32.535 102.325 32.825 102.370 ;
        RECT 38.130 102.230 38.270 102.370 ;
        RECT 38.515 102.370 43.880 102.510 ;
        RECT 38.515 102.325 38.805 102.370 ;
        RECT 43.560 102.310 43.880 102.370 ;
        RECT 59.675 102.325 59.965 102.555 ;
        RECT 62.000 102.510 62.290 102.555 ;
        RECT 64.100 102.510 64.390 102.555 ;
        RECT 65.670 102.510 65.960 102.555 ;
        RECT 62.000 102.370 65.960 102.510 ;
        RECT 62.000 102.325 62.290 102.370 ;
        RECT 64.100 102.325 64.390 102.370 ;
        RECT 65.670 102.325 65.960 102.370 ;
        RECT 75.315 102.510 75.605 102.555 ;
        RECT 76.235 102.510 76.525 102.555 ;
        RECT 75.315 102.370 76.525 102.510 ;
        RECT 75.315 102.325 75.605 102.370 ;
        RECT 76.235 102.325 76.525 102.370 ;
        RECT 78.060 102.510 78.380 102.570 ;
        RECT 78.610 102.510 78.750 102.665 ;
        RECT 78.060 102.370 78.750 102.510 ;
        RECT 18.260 102.170 18.580 102.230 ;
        RECT 19.195 102.170 19.485 102.215 ;
        RECT 18.260 102.030 19.485 102.170 ;
        RECT 18.260 101.970 18.580 102.030 ;
        RECT 19.195 101.985 19.485 102.030 ;
        RECT 26.080 102.170 26.400 102.230 ;
        RECT 26.555 102.170 26.845 102.215 ;
        RECT 26.080 102.030 26.845 102.170 ;
        RECT 26.080 101.970 26.400 102.030 ;
        RECT 26.555 101.985 26.845 102.030 ;
        RECT 27.460 102.170 27.780 102.230 ;
        RECT 33.440 102.170 33.760 102.230 ;
        RECT 27.460 102.030 33.760 102.170 ;
        RECT 27.460 101.970 27.780 102.030 ;
        RECT 33.440 101.970 33.760 102.030 ;
        RECT 33.900 101.970 34.220 102.230 ;
        RECT 34.820 102.170 35.140 102.230 ;
        RECT 36.675 102.170 36.965 102.215 ;
        RECT 34.820 102.030 36.965 102.170 ;
        RECT 34.820 101.970 35.140 102.030 ;
        RECT 36.675 101.985 36.965 102.030 ;
        RECT 38.040 101.970 38.360 102.230 ;
        RECT 41.275 102.170 41.565 102.215 ;
        RECT 44.480 102.170 44.800 102.230 ;
        RECT 41.275 102.030 44.800 102.170 ;
        RECT 41.275 101.985 41.565 102.030 ;
        RECT 44.480 101.970 44.800 102.030 ;
        RECT 58.740 101.970 59.060 102.230 ;
        RECT 59.750 102.170 59.890 102.325 ;
        RECT 78.060 102.310 78.380 102.370 ;
        RECT 66.100 102.170 66.420 102.230 ;
        RECT 59.750 102.030 66.420 102.170 ;
        RECT 66.100 101.970 66.420 102.030 ;
        RECT 75.760 101.970 76.080 102.230 ;
        RECT 79.530 102.170 79.670 102.665 ;
        RECT 80.860 102.510 81.150 102.555 ;
        RECT 82.960 102.510 83.250 102.555 ;
        RECT 84.530 102.510 84.820 102.555 ;
        RECT 80.860 102.370 84.820 102.510 ;
        RECT 80.860 102.325 81.150 102.370 ;
        RECT 82.960 102.325 83.250 102.370 ;
        RECT 84.530 102.325 84.820 102.370 ;
        RECT 85.420 102.170 85.740 102.230 ;
        RECT 86.890 102.170 87.030 102.710 ;
        RECT 90.495 102.665 90.785 102.710 ;
        RECT 92.780 102.650 93.100 102.710 ;
        RECT 94.175 102.665 94.465 102.895 ;
        RECT 95.080 102.650 95.400 102.910 ;
        RECT 105.290 102.895 105.430 103.050 ;
        RECT 105.660 103.050 112.330 103.190 ;
        RECT 105.660 102.990 105.980 103.050 ;
        RECT 95.975 102.850 96.265 102.895 ;
        RECT 97.165 102.850 97.455 102.895 ;
        RECT 99.685 102.850 99.975 102.895 ;
        RECT 95.975 102.710 99.975 102.850 ;
        RECT 95.975 102.665 96.265 102.710 ;
        RECT 97.165 102.665 97.455 102.710 ;
        RECT 99.685 102.665 99.975 102.710 ;
        RECT 104.755 102.665 105.045 102.895 ;
        RECT 105.215 102.665 105.505 102.895 ;
        RECT 93.255 102.325 93.545 102.555 ;
        RECT 95.580 102.510 95.870 102.555 ;
        RECT 97.680 102.510 97.970 102.555 ;
        RECT 99.250 102.510 99.540 102.555 ;
        RECT 102.455 102.510 102.745 102.555 ;
        RECT 95.580 102.370 99.540 102.510 ;
        RECT 95.580 102.325 95.870 102.370 ;
        RECT 97.680 102.325 97.970 102.370 ;
        RECT 99.250 102.325 99.540 102.370 ;
        RECT 99.770 102.370 102.745 102.510 ;
        RECT 79.530 102.030 87.030 102.170 ;
        RECT 85.420 101.970 85.740 102.030 ;
        RECT 87.260 101.970 87.580 102.230 ;
        RECT 87.720 101.970 88.040 102.230 ;
        RECT 93.330 102.170 93.470 102.325 ;
        RECT 99.770 102.170 99.910 102.370 ;
        RECT 102.455 102.325 102.745 102.370 ;
        RECT 93.330 102.030 99.910 102.170 ;
        RECT 101.995 102.170 102.285 102.215 ;
        RECT 102.900 102.170 103.220 102.230 ;
        RECT 104.830 102.170 104.970 102.665 ;
        RECT 107.040 102.650 107.360 102.910 ;
        RECT 107.935 102.850 108.225 102.895 ;
        RECT 109.125 102.850 109.415 102.895 ;
        RECT 111.645 102.850 111.935 102.895 ;
        RECT 107.935 102.710 111.935 102.850 ;
        RECT 112.190 102.850 112.330 103.050 ;
        RECT 116.700 103.050 121.160 103.190 ;
        RECT 116.700 102.990 117.020 103.050 ;
        RECT 120.840 102.990 121.160 103.050 ;
        RECT 125.990 103.050 136.705 103.190 ;
        RECT 117.635 102.850 117.925 102.895 ;
        RECT 112.190 102.710 117.925 102.850 ;
        RECT 107.935 102.665 108.225 102.710 ;
        RECT 109.125 102.665 109.415 102.710 ;
        RECT 111.645 102.665 111.935 102.710 ;
        RECT 117.635 102.665 117.925 102.710 ;
        RECT 123.155 102.850 123.445 102.895 ;
        RECT 123.600 102.850 123.920 102.910 ;
        RECT 123.155 102.710 123.920 102.850 ;
        RECT 123.155 102.665 123.445 102.710 ;
        RECT 107.540 102.510 107.830 102.555 ;
        RECT 109.640 102.510 109.930 102.555 ;
        RECT 111.210 102.510 111.500 102.555 ;
        RECT 107.540 102.370 111.500 102.510 ;
        RECT 107.540 102.325 107.830 102.370 ;
        RECT 109.640 102.325 109.930 102.370 ;
        RECT 111.210 102.325 111.500 102.370 ;
        RECT 113.955 102.510 114.245 102.555 ;
        RECT 116.700 102.510 117.020 102.570 ;
        RECT 113.955 102.370 117.020 102.510 ;
        RECT 117.710 102.510 117.850 102.665 ;
        RECT 123.600 102.650 123.920 102.710 ;
        RECT 124.075 102.850 124.365 102.895 ;
        RECT 124.520 102.850 124.840 102.910 ;
        RECT 124.075 102.710 124.840 102.850 ;
        RECT 124.075 102.665 124.365 102.710 ;
        RECT 124.520 102.650 124.840 102.710 ;
        RECT 125.990 102.510 126.130 103.050 ;
        RECT 126.375 102.665 126.665 102.895 ;
        RECT 127.255 102.850 127.545 102.895 ;
        RECT 128.445 102.850 128.735 102.895 ;
        RECT 130.965 102.850 131.255 102.895 ;
        RECT 127.255 102.710 131.255 102.850 ;
        RECT 127.255 102.665 127.545 102.710 ;
        RECT 128.445 102.665 128.735 102.710 ;
        RECT 130.965 102.665 131.255 102.710 ;
        RECT 133.720 102.850 134.040 102.910 ;
        RECT 135.115 102.850 135.405 102.895 ;
        RECT 133.720 102.710 135.405 102.850 ;
        RECT 117.710 102.370 126.130 102.510 ;
        RECT 113.955 102.325 114.245 102.370 ;
        RECT 116.700 102.310 117.020 102.370 ;
        RECT 101.995 102.030 104.970 102.170 ;
        RECT 116.240 102.170 116.560 102.230 ;
        RECT 120.855 102.170 121.145 102.215 ;
        RECT 116.240 102.030 121.145 102.170 ;
        RECT 126.450 102.170 126.590 102.665 ;
        RECT 133.720 102.650 134.040 102.710 ;
        RECT 135.115 102.665 135.405 102.710 ;
        RECT 126.860 102.510 127.150 102.555 ;
        RECT 128.960 102.510 129.250 102.555 ;
        RECT 130.530 102.510 130.820 102.555 ;
        RECT 136.020 102.510 136.340 102.570 ;
        RECT 126.860 102.370 130.820 102.510 ;
        RECT 126.860 102.325 127.150 102.370 ;
        RECT 128.960 102.325 129.250 102.370 ;
        RECT 130.530 102.325 130.820 102.370 ;
        RECT 131.050 102.370 136.340 102.510 ;
        RECT 136.565 102.510 136.705 103.050 ;
        RECT 138.335 103.050 140.850 103.190 ;
        RECT 138.335 103.005 138.625 103.050 ;
        RECT 139.240 102.650 139.560 102.910 ;
        RECT 140.710 102.850 140.850 103.050 ;
        RECT 141.095 103.005 141.385 103.235 ;
        RECT 141.555 103.005 141.845 103.235 ;
        RECT 141.630 102.850 141.770 103.005 ;
        RECT 142.000 102.990 142.320 103.250 ;
        RECT 142.935 103.190 143.225 103.235 ;
        RECT 143.840 103.190 144.160 103.250 ;
        RECT 142.935 103.050 144.160 103.190 ;
        RECT 142.935 103.005 143.225 103.050 ;
        RECT 143.840 102.990 144.160 103.050 ;
        RECT 140.710 102.710 141.770 102.850 ;
        RECT 141.170 102.570 141.310 102.710 ;
        RECT 139.700 102.510 140.020 102.570 ;
        RECT 136.565 102.370 140.020 102.510 ;
        RECT 131.050 102.170 131.190 102.370 ;
        RECT 136.020 102.310 136.340 102.370 ;
        RECT 139.700 102.310 140.020 102.370 ;
        RECT 141.080 102.310 141.400 102.570 ;
        RECT 126.450 102.030 131.190 102.170 ;
        RECT 101.995 101.985 102.285 102.030 ;
        RECT 102.900 101.970 103.220 102.030 ;
        RECT 116.240 101.970 116.560 102.030 ;
        RECT 120.855 101.985 121.145 102.030 ;
        RECT 133.260 101.970 133.580 102.230 ;
        RECT 137.400 102.170 137.720 102.230 ;
        RECT 140.175 102.170 140.465 102.215 ;
        RECT 137.400 102.030 140.465 102.170 ;
        RECT 137.400 101.970 137.720 102.030 ;
        RECT 140.175 101.985 140.465 102.030 ;
        RECT 144.300 102.170 144.620 102.230 ;
        RECT 144.775 102.170 145.065 102.215 ;
        RECT 144.300 102.030 145.065 102.170 ;
        RECT 144.300 101.970 144.620 102.030 ;
        RECT 144.775 101.985 145.065 102.030 ;
        RECT 17.270 101.350 146.990 101.830 ;
        RECT 31.615 101.150 31.905 101.195 ;
        RECT 32.060 101.150 32.380 101.210 ;
        RECT 42.180 101.150 42.500 101.210 ;
        RECT 61.500 101.150 61.820 101.210 ;
        RECT 31.615 101.010 32.380 101.150 ;
        RECT 31.615 100.965 31.905 101.010 ;
        RECT 32.060 100.950 32.380 101.010 ;
        RECT 36.290 101.010 42.500 101.150 ;
        RECT 21.980 100.810 22.270 100.855 ;
        RECT 24.080 100.810 24.370 100.855 ;
        RECT 25.650 100.810 25.940 100.855 ;
        RECT 21.980 100.670 25.940 100.810 ;
        RECT 21.980 100.625 22.270 100.670 ;
        RECT 24.080 100.625 24.370 100.670 ;
        RECT 25.650 100.625 25.940 100.670 ;
        RECT 22.375 100.470 22.665 100.515 ;
        RECT 23.565 100.470 23.855 100.515 ;
        RECT 26.085 100.470 26.375 100.515 ;
        RECT 35.280 100.470 35.600 100.530 ;
        RECT 22.375 100.330 26.375 100.470 ;
        RECT 22.375 100.285 22.665 100.330 ;
        RECT 23.565 100.285 23.855 100.330 ;
        RECT 26.085 100.285 26.375 100.330 ;
        RECT 32.150 100.330 35.600 100.470 ;
        RECT 32.150 100.190 32.290 100.330 ;
        RECT 21.495 100.130 21.785 100.175 ;
        RECT 27.000 100.130 27.320 100.190 ;
        RECT 21.495 99.990 27.320 100.130 ;
        RECT 21.495 99.945 21.785 99.990 ;
        RECT 27.000 99.930 27.320 99.990 ;
        RECT 27.460 100.130 27.780 100.190 ;
        RECT 28.855 100.130 29.145 100.175 ;
        RECT 27.460 99.990 29.145 100.130 ;
        RECT 27.460 99.930 27.780 99.990 ;
        RECT 28.855 99.945 29.145 99.990 ;
        RECT 29.775 100.130 30.065 100.175 ;
        RECT 32.060 100.130 32.380 100.190 ;
        RECT 29.775 99.990 32.380 100.130 ;
        RECT 29.775 99.945 30.065 99.990 ;
        RECT 32.060 99.930 32.380 99.990 ;
        RECT 32.520 99.930 32.840 100.190 ;
        RECT 33.900 99.930 34.220 100.190 ;
        RECT 34.910 100.175 35.050 100.330 ;
        RECT 35.280 100.270 35.600 100.330 ;
        RECT 36.290 100.175 36.430 101.010 ;
        RECT 42.180 100.950 42.500 101.010 ;
        RECT 57.910 101.010 61.820 101.150 ;
        RECT 41.260 100.610 41.580 100.870 ;
        RECT 48.160 100.610 48.480 100.870 ;
        RECT 38.975 100.470 39.265 100.515 ;
        RECT 37.670 100.330 39.265 100.470 ;
        RECT 37.670 100.175 37.810 100.330 ;
        RECT 38.975 100.285 39.265 100.330 ;
        RECT 39.420 100.470 39.740 100.530 ;
        RECT 41.350 100.470 41.490 100.610 ;
        RECT 57.910 100.515 58.050 101.010 ;
        RECT 61.500 100.950 61.820 101.010 ;
        RECT 64.735 101.150 65.025 101.195 ;
        RECT 68.400 101.150 68.720 101.210 ;
        RECT 71.160 101.150 71.480 101.210 ;
        RECT 84.975 101.150 85.265 101.195 ;
        RECT 90.480 101.150 90.800 101.210 ;
        RECT 64.735 101.010 71.480 101.150 ;
        RECT 64.735 100.965 65.025 101.010 ;
        RECT 68.400 100.950 68.720 101.010 ;
        RECT 71.160 100.950 71.480 101.010 ;
        RECT 71.710 101.010 82.430 101.150 ;
        RECT 58.320 100.810 58.610 100.855 ;
        RECT 60.420 100.810 60.710 100.855 ;
        RECT 61.990 100.810 62.280 100.855 ;
        RECT 58.320 100.670 62.280 100.810 ;
        RECT 58.320 100.625 58.610 100.670 ;
        RECT 60.420 100.625 60.710 100.670 ;
        RECT 61.990 100.625 62.280 100.670 ;
        RECT 65.680 100.810 65.970 100.855 ;
        RECT 67.780 100.810 68.070 100.855 ;
        RECT 69.350 100.810 69.640 100.855 ;
        RECT 65.680 100.670 69.640 100.810 ;
        RECT 65.680 100.625 65.970 100.670 ;
        RECT 67.780 100.625 68.070 100.670 ;
        RECT 69.350 100.625 69.640 100.670 ;
        RECT 48.635 100.470 48.925 100.515 ;
        RECT 39.420 100.330 42.410 100.470 ;
        RECT 39.420 100.270 39.740 100.330 ;
        RECT 34.835 99.945 35.125 100.175 ;
        RECT 36.215 99.945 36.505 100.175 ;
        RECT 37.595 99.945 37.885 100.175 ;
        RECT 38.515 99.945 38.805 100.175 ;
        RECT 39.895 100.130 40.185 100.175 ;
        RECT 40.340 100.130 40.660 100.190 ;
        RECT 42.270 100.175 42.410 100.330 ;
        RECT 45.030 100.330 48.925 100.470 ;
        RECT 45.030 100.175 45.170 100.330 ;
        RECT 48.635 100.285 48.925 100.330 ;
        RECT 57.835 100.285 58.125 100.515 ;
        RECT 58.715 100.470 59.005 100.515 ;
        RECT 59.905 100.470 60.195 100.515 ;
        RECT 62.425 100.470 62.715 100.515 ;
        RECT 58.715 100.330 62.715 100.470 ;
        RECT 58.715 100.285 59.005 100.330 ;
        RECT 59.905 100.285 60.195 100.330 ;
        RECT 62.425 100.285 62.715 100.330 ;
        RECT 66.075 100.470 66.365 100.515 ;
        RECT 67.265 100.470 67.555 100.515 ;
        RECT 69.785 100.470 70.075 100.515 ;
        RECT 66.075 100.330 70.075 100.470 ;
        RECT 66.075 100.285 66.365 100.330 ;
        RECT 67.265 100.285 67.555 100.330 ;
        RECT 69.785 100.285 70.075 100.330 ;
        RECT 39.895 99.990 40.660 100.130 ;
        RECT 39.895 99.945 40.185 99.990 ;
        RECT 22.830 99.790 23.120 99.835 ;
        RECT 26.540 99.790 26.860 99.850 ;
        RECT 22.830 99.650 26.860 99.790 ;
        RECT 22.830 99.605 23.120 99.650 ;
        RECT 26.540 99.590 26.860 99.650 ;
        RECT 33.440 99.790 33.760 99.850 ;
        RECT 36.660 99.790 36.980 99.850 ;
        RECT 33.440 99.650 36.980 99.790 ;
        RECT 38.590 99.790 38.730 99.945 ;
        RECT 40.340 99.930 40.660 99.990 ;
        RECT 41.275 99.945 41.565 100.175 ;
        RECT 42.195 99.945 42.485 100.175 ;
        RECT 43.575 99.945 43.865 100.175 ;
        RECT 44.955 99.945 45.245 100.175 ;
        RECT 45.875 100.130 46.165 100.175 ;
        RECT 46.780 100.130 47.100 100.190 ;
        RECT 45.875 99.990 47.100 100.130 ;
        RECT 45.875 99.945 46.165 99.990 ;
        RECT 40.800 99.790 41.120 99.850 ;
        RECT 38.590 99.650 41.120 99.790 ;
        RECT 41.350 99.790 41.490 99.945 ;
        RECT 42.655 99.790 42.945 99.835 ;
        RECT 41.350 99.650 42.945 99.790 ;
        RECT 33.440 99.590 33.760 99.650 ;
        RECT 36.660 99.590 36.980 99.650 ;
        RECT 40.800 99.590 41.120 99.650 ;
        RECT 42.655 99.605 42.945 99.650 ;
        RECT 28.380 99.250 28.700 99.510 ;
        RECT 29.315 99.450 29.605 99.495 ;
        RECT 31.140 99.450 31.460 99.510 ;
        RECT 29.315 99.310 31.460 99.450 ;
        RECT 29.315 99.265 29.605 99.310 ;
        RECT 31.140 99.250 31.460 99.310 ;
        RECT 35.280 99.250 35.600 99.510 ;
        RECT 39.880 99.450 40.200 99.510 ;
        RECT 43.650 99.450 43.790 99.945 ;
        RECT 46.780 99.930 47.100 99.990 ;
        RECT 59.170 99.945 59.460 100.175 ;
        RECT 61.500 100.130 61.820 100.190 ;
        RECT 65.195 100.130 65.485 100.175 ;
        RECT 61.500 99.990 65.485 100.130 ;
        RECT 46.335 99.605 46.625 99.835 ;
        RECT 58.740 99.790 59.060 99.850 ;
        RECT 59.290 99.790 59.430 99.945 ;
        RECT 61.500 99.930 61.820 99.990 ;
        RECT 65.195 99.945 65.485 99.990 ;
        RECT 68.400 100.130 68.720 100.190 ;
        RECT 70.240 100.130 70.560 100.190 ;
        RECT 71.710 100.130 71.850 101.010 ;
        RECT 74.880 100.810 75.170 100.855 ;
        RECT 76.980 100.810 77.270 100.855 ;
        RECT 78.550 100.810 78.840 100.855 ;
        RECT 74.880 100.670 78.840 100.810 ;
        RECT 74.880 100.625 75.170 100.670 ;
        RECT 76.980 100.625 77.270 100.670 ;
        RECT 78.550 100.625 78.840 100.670 ;
        RECT 75.275 100.470 75.565 100.515 ;
        RECT 76.465 100.470 76.755 100.515 ;
        RECT 78.985 100.470 79.275 100.515 ;
        RECT 75.275 100.330 79.275 100.470 ;
        RECT 75.275 100.285 75.565 100.330 ;
        RECT 76.465 100.285 76.755 100.330 ;
        RECT 78.985 100.285 79.275 100.330 ;
        RECT 68.400 99.990 71.850 100.130 ;
        RECT 72.555 100.130 72.845 100.175 ;
        RECT 73.000 100.130 73.320 100.190 ;
        RECT 72.555 99.990 73.320 100.130 ;
        RECT 68.400 99.930 68.720 99.990 ;
        RECT 70.240 99.930 70.560 99.990 ;
        RECT 72.555 99.945 72.845 99.990 ;
        RECT 73.000 99.930 73.320 99.990 ;
        RECT 74.395 100.130 74.685 100.175 ;
        RECT 80.820 100.130 81.140 100.190 ;
        RECT 82.290 100.175 82.430 101.010 ;
        RECT 84.975 101.010 90.800 101.150 ;
        RECT 84.975 100.965 85.265 101.010 ;
        RECT 90.480 100.950 90.800 101.010 ;
        RECT 92.320 101.150 92.640 101.210 ;
        RECT 94.175 101.150 94.465 101.195 ;
        RECT 92.320 101.010 94.465 101.150 ;
        RECT 92.320 100.950 92.640 101.010 ;
        RECT 94.175 100.965 94.465 101.010 ;
        RECT 102.915 101.150 103.205 101.195 ;
        RECT 104.280 101.150 104.600 101.210 ;
        RECT 102.915 101.010 104.600 101.150 ;
        RECT 102.915 100.965 103.205 101.010 ;
        RECT 104.280 100.950 104.600 101.010 ;
        RECT 106.580 100.950 106.900 101.210 ;
        RECT 123.600 101.150 123.920 101.210 ;
        RECT 125.900 101.150 126.220 101.210 ;
        RECT 129.595 101.150 129.885 101.195 ;
        RECT 136.020 101.150 136.340 101.210 ;
        RECT 123.600 101.010 129.885 101.150 ;
        RECT 123.600 100.950 123.920 101.010 ;
        RECT 125.900 100.950 126.220 101.010 ;
        RECT 129.595 100.965 129.885 101.010 ;
        RECT 134.270 101.010 136.340 101.150 ;
        RECT 87.760 100.810 88.050 100.855 ;
        RECT 89.860 100.810 90.150 100.855 ;
        RECT 91.430 100.810 91.720 100.855 ;
        RECT 82.795 100.670 87.490 100.810 ;
        RECT 74.395 99.990 81.140 100.130 ;
        RECT 74.395 99.945 74.685 99.990 ;
        RECT 80.820 99.930 81.140 99.990 ;
        RECT 82.215 99.945 82.505 100.175 ;
        RECT 58.740 99.650 59.430 99.790 ;
        RECT 66.530 99.790 66.820 99.835 ;
        RECT 67.940 99.790 68.260 99.850 ;
        RECT 66.530 99.650 68.260 99.790 ;
        RECT 39.880 99.310 43.790 99.450 ;
        RECT 45.860 99.450 46.180 99.510 ;
        RECT 46.410 99.450 46.550 99.605 ;
        RECT 58.740 99.590 59.060 99.650 ;
        RECT 66.530 99.605 66.820 99.650 ;
        RECT 67.940 99.590 68.260 99.650 ;
        RECT 69.780 99.790 70.100 99.850 ;
        RECT 75.760 99.835 76.080 99.850 ;
        RECT 75.730 99.790 76.080 99.835 ;
        RECT 69.780 99.650 73.690 99.790 ;
        RECT 75.565 99.650 76.080 99.790 ;
        RECT 80.910 99.790 81.050 99.930 ;
        RECT 82.795 99.850 82.935 100.670 ;
        RECT 84.960 100.470 85.280 100.530 ;
        RECT 87.350 100.515 87.490 100.670 ;
        RECT 87.760 100.670 91.720 100.810 ;
        RECT 87.760 100.625 88.050 100.670 ;
        RECT 89.860 100.625 90.150 100.670 ;
        RECT 91.430 100.625 91.720 100.670 ;
        RECT 93.700 100.810 94.020 100.870 ;
        RECT 94.635 100.810 94.925 100.855 ;
        RECT 93.700 100.670 94.925 100.810 ;
        RECT 93.700 100.610 94.020 100.670 ;
        RECT 94.635 100.625 94.925 100.670 ;
        RECT 96.500 100.810 96.790 100.855 ;
        RECT 98.600 100.810 98.890 100.855 ;
        RECT 100.170 100.810 100.460 100.855 ;
        RECT 105.200 100.810 105.520 100.870 ;
        RECT 108.460 100.810 108.750 100.855 ;
        RECT 110.560 100.810 110.850 100.855 ;
        RECT 112.130 100.810 112.420 100.855 ;
        RECT 96.500 100.670 100.460 100.810 ;
        RECT 96.500 100.625 96.790 100.670 ;
        RECT 98.600 100.625 98.890 100.670 ;
        RECT 100.170 100.625 100.460 100.670 ;
        RECT 102.530 100.670 105.890 100.810 ;
        RECT 83.210 100.330 85.280 100.470 ;
        RECT 83.210 100.175 83.350 100.330 ;
        RECT 84.960 100.270 85.280 100.330 ;
        RECT 87.275 100.285 87.565 100.515 ;
        RECT 88.155 100.470 88.445 100.515 ;
        RECT 89.345 100.470 89.635 100.515 ;
        RECT 91.865 100.470 92.155 100.515 ;
        RECT 88.155 100.330 92.155 100.470 ;
        RECT 88.155 100.285 88.445 100.330 ;
        RECT 89.345 100.285 89.635 100.330 ;
        RECT 91.865 100.285 92.155 100.330 ;
        RECT 95.080 100.470 95.400 100.530 ;
        RECT 96.015 100.470 96.305 100.515 ;
        RECT 95.080 100.330 96.305 100.470 ;
        RECT 95.080 100.270 95.400 100.330 ;
        RECT 96.015 100.285 96.305 100.330 ;
        RECT 96.895 100.470 97.185 100.515 ;
        RECT 98.085 100.470 98.375 100.515 ;
        RECT 100.605 100.470 100.895 100.515 ;
        RECT 96.895 100.330 100.895 100.470 ;
        RECT 96.895 100.285 97.185 100.330 ;
        RECT 98.085 100.285 98.375 100.330 ;
        RECT 100.605 100.285 100.895 100.330 ;
        RECT 83.135 99.945 83.425 100.175 ;
        RECT 84.055 99.945 84.345 100.175 ;
        RECT 82.660 99.790 82.980 99.850 ;
        RECT 80.910 99.650 82.980 99.790 ;
        RECT 69.780 99.590 70.100 99.650 ;
        RECT 45.860 99.310 46.550 99.450 ;
        RECT 39.880 99.250 40.200 99.310 ;
        RECT 45.860 99.250 46.180 99.310 ;
        RECT 72.080 99.250 72.400 99.510 ;
        RECT 73.550 99.495 73.690 99.650 ;
        RECT 75.730 99.605 76.080 99.650 ;
        RECT 75.760 99.590 76.080 99.605 ;
        RECT 82.660 99.590 82.980 99.650 ;
        RECT 83.595 99.605 83.885 99.835 ;
        RECT 73.475 99.265 73.765 99.495 ;
        RECT 78.060 99.450 78.380 99.510 ;
        RECT 81.295 99.450 81.585 99.495 ;
        RECT 83.670 99.450 83.810 99.605 ;
        RECT 78.060 99.310 83.810 99.450 ;
        RECT 84.130 99.450 84.270 99.945 ;
        RECT 95.540 99.930 95.860 100.190 ;
        RECT 102.530 100.130 102.670 100.670 ;
        RECT 105.200 100.610 105.520 100.670 ;
        RECT 102.900 100.470 103.220 100.530 ;
        RECT 102.900 100.330 104.050 100.470 ;
        RECT 102.900 100.270 103.220 100.330 ;
        RECT 103.910 100.175 104.050 100.330 ;
        RECT 103.375 100.130 103.665 100.175 ;
        RECT 97.010 99.990 102.670 100.130 ;
        RECT 102.990 99.990 103.665 100.130 ;
        RECT 88.610 99.790 88.900 99.835 ;
        RECT 89.560 99.790 89.880 99.850 ;
        RECT 93.240 99.790 93.560 99.850 ;
        RECT 97.010 99.790 97.150 99.990 ;
        RECT 88.610 99.650 89.880 99.790 ;
        RECT 88.610 99.605 88.900 99.650 ;
        RECT 89.560 99.590 89.880 99.650 ;
        RECT 90.570 99.650 97.150 99.790 ;
        RECT 97.350 99.790 97.640 99.835 ;
        RECT 101.520 99.790 101.840 99.850 ;
        RECT 97.350 99.650 101.840 99.790 ;
        RECT 89.100 99.450 89.420 99.510 ;
        RECT 90.570 99.450 90.710 99.650 ;
        RECT 93.240 99.590 93.560 99.650 ;
        RECT 97.350 99.605 97.640 99.650 ;
        RECT 101.520 99.590 101.840 99.650 ;
        RECT 84.130 99.310 90.710 99.450 ;
        RECT 94.160 99.450 94.480 99.510 ;
        RECT 102.990 99.450 103.130 99.990 ;
        RECT 103.375 99.945 103.665 99.990 ;
        RECT 103.840 99.945 104.130 100.175 ;
        RECT 104.280 100.130 104.600 100.190 ;
        RECT 105.750 100.175 105.890 100.670 ;
        RECT 108.460 100.670 112.420 100.810 ;
        RECT 108.460 100.625 108.750 100.670 ;
        RECT 110.560 100.625 110.850 100.670 ;
        RECT 112.130 100.625 112.420 100.670 ;
        RECT 115.820 100.810 116.110 100.855 ;
        RECT 117.920 100.810 118.210 100.855 ;
        RECT 119.490 100.810 119.780 100.855 ;
        RECT 115.820 100.670 119.780 100.810 ;
        RECT 115.820 100.625 116.110 100.670 ;
        RECT 117.920 100.625 118.210 100.670 ;
        RECT 119.490 100.625 119.780 100.670 ;
        RECT 123.180 100.810 123.470 100.855 ;
        RECT 125.280 100.810 125.570 100.855 ;
        RECT 126.850 100.810 127.140 100.855 ;
        RECT 123.180 100.670 127.140 100.810 ;
        RECT 123.180 100.625 123.470 100.670 ;
        RECT 125.280 100.625 125.570 100.670 ;
        RECT 126.850 100.625 127.140 100.670 ;
        RECT 130.960 100.610 131.280 100.870 ;
        RECT 108.855 100.470 109.145 100.515 ;
        RECT 110.045 100.470 110.335 100.515 ;
        RECT 112.565 100.470 112.855 100.515 ;
        RECT 108.855 100.330 112.855 100.470 ;
        RECT 108.855 100.285 109.145 100.330 ;
        RECT 110.045 100.285 110.335 100.330 ;
        RECT 112.565 100.285 112.855 100.330 ;
        RECT 116.215 100.470 116.505 100.515 ;
        RECT 117.405 100.470 117.695 100.515 ;
        RECT 119.925 100.470 120.215 100.515 ;
        RECT 116.215 100.330 120.215 100.470 ;
        RECT 116.215 100.285 116.505 100.330 ;
        RECT 117.405 100.285 117.695 100.330 ;
        RECT 119.925 100.285 120.215 100.330 ;
        RECT 123.575 100.470 123.865 100.515 ;
        RECT 124.765 100.470 125.055 100.515 ;
        RECT 127.285 100.470 127.575 100.515 ;
        RECT 123.575 100.330 127.575 100.470 ;
        RECT 123.575 100.285 123.865 100.330 ;
        RECT 124.765 100.285 125.055 100.330 ;
        RECT 127.285 100.285 127.575 100.330 ;
        RECT 132.355 100.470 132.645 100.515 ;
        RECT 133.720 100.470 134.040 100.530 ;
        RECT 134.270 100.515 134.410 101.010 ;
        RECT 136.020 100.950 136.340 101.010 ;
        RECT 141.080 100.950 141.400 101.210 ;
        RECT 134.680 100.810 134.970 100.855 ;
        RECT 136.780 100.810 137.070 100.855 ;
        RECT 138.350 100.810 138.640 100.855 ;
        RECT 134.680 100.670 138.640 100.810 ;
        RECT 134.680 100.625 134.970 100.670 ;
        RECT 136.780 100.625 137.070 100.670 ;
        RECT 138.350 100.625 138.640 100.670 ;
        RECT 132.355 100.330 134.040 100.470 ;
        RECT 132.355 100.285 132.645 100.330 ;
        RECT 133.720 100.270 134.040 100.330 ;
        RECT 134.195 100.285 134.485 100.515 ;
        RECT 135.075 100.470 135.365 100.515 ;
        RECT 136.265 100.470 136.555 100.515 ;
        RECT 138.785 100.470 139.075 100.515 ;
        RECT 135.075 100.330 139.075 100.470 ;
        RECT 135.075 100.285 135.365 100.330 ;
        RECT 136.265 100.285 136.555 100.330 ;
        RECT 138.785 100.285 139.075 100.330 ;
        RECT 144.775 100.470 145.065 100.515 ;
        RECT 145.220 100.470 145.540 100.530 ;
        RECT 144.775 100.330 145.540 100.470 ;
        RECT 144.775 100.285 145.065 100.330 ;
        RECT 145.220 100.270 145.540 100.330 ;
        RECT 105.215 100.130 105.505 100.175 ;
        RECT 104.280 99.990 105.505 100.130 ;
        RECT 104.280 99.930 104.600 99.990 ;
        RECT 105.215 99.945 105.505 99.990 ;
        RECT 105.700 99.945 105.990 100.175 ;
        RECT 107.040 100.130 107.360 100.190 ;
        RECT 107.975 100.130 108.265 100.175 ;
        RECT 115.335 100.130 115.625 100.175 ;
        RECT 122.680 100.130 123.000 100.190 ;
        RECT 107.040 99.990 123.000 100.130 ;
        RECT 107.040 99.930 107.360 99.990 ;
        RECT 107.975 99.945 108.265 99.990 ;
        RECT 115.335 99.945 115.625 99.990 ;
        RECT 122.680 99.930 123.000 99.990 ;
        RECT 135.530 100.130 135.820 100.175 ;
        RECT 136.940 100.130 137.260 100.190 ;
        RECT 135.530 99.990 137.260 100.130 ;
        RECT 135.530 99.945 135.820 99.990 ;
        RECT 136.940 99.930 137.260 99.990 ;
        RECT 104.740 99.590 105.060 99.850 ;
        RECT 107.500 99.790 107.820 99.850 ;
        RECT 109.200 99.790 109.490 99.835 ;
        RECT 107.500 99.650 109.490 99.790 ;
        RECT 107.500 99.590 107.820 99.650 ;
        RECT 109.200 99.605 109.490 99.650 ;
        RECT 115.780 99.790 116.100 99.850 ;
        RECT 124.060 99.835 124.380 99.850 ;
        RECT 116.560 99.790 116.850 99.835 ;
        RECT 115.780 99.650 116.850 99.790 ;
        RECT 115.780 99.590 116.100 99.650 ;
        RECT 116.560 99.605 116.850 99.650 ;
        RECT 124.030 99.605 124.380 99.835 ;
        RECT 143.395 99.790 143.685 99.835 ;
        RECT 124.060 99.590 124.380 99.605 ;
        RECT 137.950 99.650 143.685 99.790 ;
        RECT 137.950 99.510 138.090 99.650 ;
        RECT 143.395 99.605 143.685 99.650 ;
        RECT 94.160 99.310 103.130 99.450 ;
        RECT 113.020 99.450 113.340 99.510 ;
        RECT 114.860 99.450 115.180 99.510 ;
        RECT 113.020 99.310 115.180 99.450 ;
        RECT 78.060 99.250 78.380 99.310 ;
        RECT 81.295 99.265 81.585 99.310 ;
        RECT 89.100 99.250 89.420 99.310 ;
        RECT 94.160 99.250 94.480 99.310 ;
        RECT 113.020 99.250 113.340 99.310 ;
        RECT 114.860 99.250 115.180 99.310 ;
        RECT 118.080 99.450 118.400 99.510 ;
        RECT 122.235 99.450 122.525 99.495 ;
        RECT 118.080 99.310 122.525 99.450 ;
        RECT 118.080 99.250 118.400 99.310 ;
        RECT 122.235 99.265 122.525 99.310 ;
        RECT 130.040 99.250 130.360 99.510 ;
        RECT 132.800 99.450 133.120 99.510 ;
        RECT 137.860 99.450 138.180 99.510 ;
        RECT 132.800 99.310 138.180 99.450 ;
        RECT 132.800 99.250 133.120 99.310 ;
        RECT 137.860 99.250 138.180 99.310 ;
        RECT 141.540 99.250 141.860 99.510 ;
        RECT 143.840 99.250 144.160 99.510 ;
        RECT 17.270 98.630 146.990 99.110 ;
        RECT 19.195 98.430 19.485 98.475 ;
        RECT 25.620 98.430 25.940 98.490 ;
        RECT 19.195 98.290 25.940 98.430 ;
        RECT 19.195 98.245 19.485 98.290 ;
        RECT 25.620 98.230 25.940 98.290 ;
        RECT 26.540 98.230 26.860 98.490 ;
        RECT 28.380 98.230 28.700 98.490 ;
        RECT 28.855 98.430 29.145 98.475 ;
        RECT 30.680 98.430 31.000 98.490 ;
        RECT 31.615 98.430 31.905 98.475 ;
        RECT 28.855 98.290 31.905 98.430 ;
        RECT 28.855 98.245 29.145 98.290 ;
        RECT 30.680 98.230 31.000 98.290 ;
        RECT 31.615 98.245 31.905 98.290 ;
        RECT 33.900 98.430 34.220 98.490 ;
        RECT 33.900 98.290 34.590 98.430 ;
        RECT 33.900 98.230 34.220 98.290 ;
        RECT 24.870 98.090 25.160 98.135 ;
        RECT 26.080 98.090 26.400 98.150 ;
        RECT 24.870 97.950 26.400 98.090 ;
        RECT 24.870 97.905 25.160 97.950 ;
        RECT 26.080 97.890 26.400 97.950 ;
        RECT 27.460 98.090 27.780 98.150 ;
        RECT 34.450 98.090 34.590 98.290 ;
        RECT 41.720 98.230 42.040 98.490 ;
        RECT 43.560 98.230 43.880 98.490 ;
        RECT 48.160 98.430 48.480 98.490 ;
        RECT 57.375 98.430 57.665 98.475 ;
        RECT 48.160 98.290 57.665 98.430 ;
        RECT 48.160 98.230 48.480 98.290 ;
        RECT 57.375 98.245 57.665 98.290 ;
        RECT 67.480 98.430 67.800 98.490 ;
        RECT 68.860 98.430 69.180 98.490 ;
        RECT 67.480 98.290 69.180 98.430 ;
        RECT 67.480 98.230 67.800 98.290 ;
        RECT 68.860 98.230 69.180 98.290 ;
        RECT 71.635 98.430 71.925 98.475 ;
        RECT 72.080 98.430 72.400 98.490 ;
        RECT 71.635 98.290 72.400 98.430 ;
        RECT 71.635 98.245 71.925 98.290 ;
        RECT 72.080 98.230 72.400 98.290 ;
        RECT 76.235 98.430 76.525 98.475 ;
        RECT 91.400 98.430 91.720 98.490 ;
        RECT 94.175 98.430 94.465 98.475 ;
        RECT 76.235 98.290 91.170 98.430 ;
        RECT 76.235 98.245 76.525 98.290 ;
        RECT 34.835 98.090 35.125 98.135 ;
        RECT 27.460 97.950 34.130 98.090 ;
        RECT 34.450 97.950 35.125 98.090 ;
        RECT 27.460 97.890 27.780 97.950 ;
        RECT 31.140 97.750 31.460 97.810 ;
        RECT 32.995 97.750 33.285 97.795 ;
        RECT 31.140 97.610 33.285 97.750 ;
        RECT 31.140 97.550 31.460 97.610 ;
        RECT 32.995 97.565 33.285 97.610 ;
        RECT 33.440 97.550 33.760 97.810 ;
        RECT 33.990 97.770 34.130 97.950 ;
        RECT 34.835 97.905 35.125 97.950 ;
        RECT 35.280 98.090 35.600 98.150 ;
        RECT 61.500 98.090 61.820 98.150 ;
        RECT 35.280 97.950 37.350 98.090 ;
        RECT 35.280 97.890 35.600 97.950 ;
        RECT 37.210 97.795 37.350 97.950 ;
        RECT 38.130 97.950 41.490 98.090 ;
        RECT 33.990 97.700 34.590 97.770 ;
        RECT 35.755 97.750 36.045 97.795 ;
        RECT 34.910 97.700 36.045 97.750 ;
        RECT 33.990 97.630 36.045 97.700 ;
        RECT 34.450 97.610 36.045 97.630 ;
        RECT 34.450 97.560 35.050 97.610 ;
        RECT 35.755 97.565 36.045 97.610 ;
        RECT 37.135 97.565 37.425 97.795 ;
        RECT 37.580 97.750 37.900 97.810 ;
        RECT 38.130 97.795 38.270 97.950 ;
        RECT 38.055 97.750 38.345 97.795 ;
        RECT 37.580 97.610 38.345 97.750 ;
        RECT 37.580 97.550 37.900 97.610 ;
        RECT 38.055 97.565 38.345 97.610 ;
        RECT 38.500 97.550 38.820 97.810 ;
        RECT 39.420 97.550 39.740 97.810 ;
        RECT 40.800 97.550 41.120 97.810 ;
        RECT 41.350 97.795 41.490 97.950 ;
        RECT 60.670 97.950 61.820 98.090 ;
        RECT 41.275 97.565 41.565 97.795 ;
        RECT 42.180 97.550 42.500 97.810 ;
        RECT 44.480 97.550 44.800 97.810 ;
        RECT 45.860 97.550 46.180 97.810 ;
        RECT 56.900 97.750 57.220 97.810 ;
        RECT 60.670 97.795 60.810 97.950 ;
        RECT 61.500 97.890 61.820 97.950 ;
        RECT 61.960 97.795 62.280 97.810 ;
        RECT 58.295 97.750 58.585 97.795 ;
        RECT 56.900 97.610 58.585 97.750 ;
        RECT 56.900 97.550 57.220 97.610 ;
        RECT 58.295 97.565 58.585 97.610 ;
        RECT 60.595 97.565 60.885 97.795 ;
        RECT 61.930 97.565 62.280 97.795 ;
        RECT 71.175 97.750 71.465 97.795 ;
        RECT 71.620 97.750 71.940 97.810 ;
        RECT 71.175 97.610 71.940 97.750 ;
        RECT 72.170 97.750 72.310 98.230 ;
        RECT 74.380 97.890 74.700 98.150 ;
        RECT 84.930 98.090 85.220 98.135 ;
        RECT 85.880 98.090 86.200 98.150 ;
        RECT 84.930 97.950 86.200 98.090 ;
        RECT 84.930 97.905 85.220 97.950 ;
        RECT 85.880 97.890 86.200 97.950 ;
        RECT 73.460 97.750 73.780 97.810 ;
        RECT 72.170 97.610 73.780 97.750 ;
        RECT 71.175 97.565 71.465 97.610 ;
        RECT 61.960 97.550 62.280 97.565 ;
        RECT 71.620 97.550 71.940 97.610 ;
        RECT 73.460 97.550 73.780 97.610 ;
        RECT 74.855 97.565 75.145 97.795 ;
        RECT 21.505 97.410 21.795 97.455 ;
        RECT 24.025 97.410 24.315 97.455 ;
        RECT 25.215 97.410 25.505 97.455 ;
        RECT 21.505 97.270 25.505 97.410 ;
        RECT 21.505 97.225 21.795 97.270 ;
        RECT 24.025 97.225 24.315 97.270 ;
        RECT 25.215 97.225 25.505 97.270 ;
        RECT 26.095 97.410 26.385 97.455 ;
        RECT 27.000 97.410 27.320 97.470 ;
        RECT 26.095 97.270 27.320 97.410 ;
        RECT 26.095 97.225 26.385 97.270 ;
        RECT 27.000 97.210 27.320 97.270 ;
        RECT 29.300 97.210 29.620 97.470 ;
        RECT 32.535 97.225 32.825 97.455 ;
        RECT 33.915 97.410 34.205 97.455 ;
        RECT 35.280 97.410 35.600 97.470 ;
        RECT 33.915 97.270 35.600 97.410 ;
        RECT 33.915 97.225 34.205 97.270 ;
        RECT 21.940 97.070 22.230 97.115 ;
        RECT 23.510 97.070 23.800 97.115 ;
        RECT 25.610 97.070 25.900 97.115 ;
        RECT 21.940 96.930 25.900 97.070 ;
        RECT 32.610 97.070 32.750 97.225 ;
        RECT 35.280 97.210 35.600 97.270 ;
        RECT 36.200 97.410 36.520 97.470 ;
        RECT 38.590 97.410 38.730 97.550 ;
        RECT 39.895 97.410 40.185 97.455 ;
        RECT 40.340 97.410 40.660 97.470 ;
        RECT 36.200 97.270 40.660 97.410 ;
        RECT 36.200 97.210 36.520 97.270 ;
        RECT 39.895 97.225 40.185 97.270 ;
        RECT 40.340 97.210 40.660 97.270 ;
        RECT 61.475 97.410 61.765 97.455 ;
        RECT 62.665 97.410 62.955 97.455 ;
        RECT 65.185 97.410 65.475 97.455 ;
        RECT 72.540 97.410 72.860 97.470 ;
        RECT 73.920 97.410 74.240 97.470 ;
        RECT 61.475 97.270 65.475 97.410 ;
        RECT 72.345 97.270 74.240 97.410 ;
        RECT 61.475 97.225 61.765 97.270 ;
        RECT 62.665 97.225 62.955 97.270 ;
        RECT 65.185 97.225 65.475 97.270 ;
        RECT 72.540 97.210 72.860 97.270 ;
        RECT 73.920 97.210 74.240 97.270 ;
        RECT 38.515 97.070 38.805 97.115 ;
        RECT 32.610 96.930 38.805 97.070 ;
        RECT 21.940 96.885 22.230 96.930 ;
        RECT 23.510 96.885 23.800 96.930 ;
        RECT 25.610 96.885 25.900 96.930 ;
        RECT 38.515 96.885 38.805 96.930 ;
        RECT 61.080 97.070 61.370 97.115 ;
        RECT 63.180 97.070 63.470 97.115 ;
        RECT 64.750 97.070 65.040 97.115 ;
        RECT 61.080 96.930 65.040 97.070 ;
        RECT 61.080 96.885 61.370 96.930 ;
        RECT 63.180 96.885 63.470 96.930 ;
        RECT 64.750 96.885 65.040 96.930 ;
        RECT 68.860 97.070 69.180 97.130 ;
        RECT 74.930 97.070 75.070 97.565 ;
        RECT 75.300 97.550 75.620 97.810 ;
        RECT 82.660 97.750 82.980 97.810 ;
        RECT 91.030 97.795 91.170 98.290 ;
        RECT 91.400 98.290 92.550 98.430 ;
        RECT 91.400 98.230 91.720 98.290 ;
        RECT 92.410 98.135 92.550 98.290 ;
        RECT 94.175 98.290 101.290 98.430 ;
        RECT 94.175 98.245 94.465 98.290 ;
        RECT 92.335 98.090 92.625 98.135 ;
        RECT 101.150 98.090 101.290 98.290 ;
        RECT 101.520 98.230 101.840 98.490 ;
        RECT 107.055 98.430 107.345 98.475 ;
        RECT 107.500 98.430 107.820 98.490 ;
        RECT 107.055 98.290 107.820 98.430 ;
        RECT 107.055 98.245 107.345 98.290 ;
        RECT 107.500 98.230 107.820 98.290 ;
        RECT 114.875 98.430 115.165 98.475 ;
        RECT 115.780 98.430 116.100 98.490 ;
        RECT 114.875 98.290 116.100 98.430 ;
        RECT 114.875 98.245 115.165 98.290 ;
        RECT 115.780 98.230 116.100 98.290 ;
        RECT 117.620 98.230 117.940 98.490 ;
        RECT 118.080 98.230 118.400 98.490 ;
        RECT 130.500 98.430 130.820 98.490 ;
        RECT 130.975 98.430 131.265 98.475 ;
        RECT 130.500 98.290 131.265 98.430 ;
        RECT 130.500 98.230 130.820 98.290 ;
        RECT 130.975 98.245 131.265 98.290 ;
        RECT 132.800 98.230 133.120 98.490 ;
        RECT 133.260 98.430 133.580 98.490 ;
        RECT 135.100 98.430 135.420 98.490 ;
        RECT 139.700 98.430 140.020 98.490 ;
        RECT 133.260 98.290 135.420 98.430 ;
        RECT 133.260 98.230 133.580 98.290 ;
        RECT 135.100 98.230 135.420 98.290 ;
        RECT 137.030 98.290 140.020 98.430 ;
        RECT 110.720 98.090 111.040 98.150 ;
        RECT 92.335 97.950 98.070 98.090 ;
        RECT 101.150 97.950 111.040 98.090 ;
        RECT 92.335 97.905 92.625 97.950 ;
        RECT 83.595 97.750 83.885 97.795 ;
        RECT 82.660 97.610 83.885 97.750 ;
        RECT 82.660 97.550 82.980 97.610 ;
        RECT 83.595 97.565 83.885 97.610 ;
        RECT 90.955 97.565 91.245 97.795 ;
        RECT 91.695 97.750 91.985 97.795 ;
        RECT 91.695 97.610 92.550 97.750 ;
        RECT 91.695 97.565 91.985 97.610 ;
        RECT 92.410 97.470 92.550 97.610 ;
        RECT 92.780 97.550 93.100 97.810 ;
        RECT 93.240 97.795 93.560 97.810 ;
        RECT 93.240 97.750 93.570 97.795 ;
        RECT 94.620 97.750 94.940 97.810 ;
        RECT 96.935 97.750 97.225 97.795 ;
        RECT 93.240 97.610 93.755 97.750 ;
        RECT 94.620 97.610 97.225 97.750 ;
        RECT 93.240 97.565 93.570 97.610 ;
        RECT 93.240 97.550 93.560 97.565 ;
        RECT 94.620 97.550 94.940 97.610 ;
        RECT 96.935 97.565 97.225 97.610 ;
        RECT 84.475 97.410 84.765 97.455 ;
        RECT 85.665 97.410 85.955 97.455 ;
        RECT 88.185 97.410 88.475 97.455 ;
        RECT 84.475 97.270 88.475 97.410 ;
        RECT 84.475 97.225 84.765 97.270 ;
        RECT 85.665 97.225 85.955 97.270 ;
        RECT 88.185 97.225 88.475 97.270 ;
        RECT 92.320 97.210 92.640 97.470 ;
        RECT 93.700 97.410 94.020 97.470 ;
        RECT 97.380 97.410 97.700 97.470 ;
        RECT 93.700 97.270 97.700 97.410 ;
        RECT 93.700 97.210 94.020 97.270 ;
        RECT 97.380 97.210 97.700 97.270 ;
        RECT 68.860 96.930 75.070 97.070 ;
        RECT 84.080 97.070 84.370 97.115 ;
        RECT 86.180 97.070 86.470 97.115 ;
        RECT 87.750 97.070 88.040 97.115 ;
        RECT 84.080 96.930 88.040 97.070 ;
        RECT 68.860 96.870 69.180 96.930 ;
        RECT 84.080 96.885 84.370 96.930 ;
        RECT 86.180 96.885 86.470 96.930 ;
        RECT 87.750 96.885 88.040 96.930 ;
        RECT 90.020 97.070 90.340 97.130 ;
        RECT 90.495 97.070 90.785 97.115 ;
        RECT 90.020 96.930 90.785 97.070 ;
        RECT 90.020 96.870 90.340 96.930 ;
        RECT 90.495 96.885 90.785 96.930 ;
        RECT 32.520 96.730 32.840 96.790 ;
        RECT 36.660 96.730 36.980 96.790 ;
        RECT 32.520 96.590 36.980 96.730 ;
        RECT 32.520 96.530 32.840 96.590 ;
        RECT 36.660 96.530 36.980 96.590 ;
        RECT 38.960 96.730 39.280 96.790 ;
        RECT 39.435 96.730 39.725 96.775 ;
        RECT 38.960 96.590 39.725 96.730 ;
        RECT 38.960 96.530 39.280 96.590 ;
        RECT 39.435 96.545 39.725 96.590 ;
        RECT 45.415 96.730 45.705 96.775 ;
        RECT 46.780 96.730 47.100 96.790 ;
        RECT 48.620 96.730 48.940 96.790 ;
        RECT 45.415 96.590 48.940 96.730 ;
        RECT 45.415 96.545 45.705 96.590 ;
        RECT 46.780 96.530 47.100 96.590 ;
        RECT 48.620 96.530 48.940 96.590 ;
        RECT 69.320 96.530 69.640 96.790 ;
        RECT 95.080 96.530 95.400 96.790 ;
        RECT 97.930 96.730 98.070 97.950 ;
        RECT 110.720 97.890 111.040 97.950 ;
        RECT 112.560 97.890 112.880 98.150 ;
        RECT 122.680 98.090 123.000 98.150 ;
        RECT 122.680 97.950 136.710 98.090 ;
        RECT 122.680 97.890 123.000 97.950 ;
        RECT 99.220 97.550 99.540 97.810 ;
        RECT 98.315 97.410 98.605 97.455 ;
        RECT 100.600 97.410 100.920 97.470 ;
        RECT 98.315 97.270 100.920 97.410 ;
        RECT 98.315 97.225 98.605 97.270 ;
        RECT 100.600 97.210 100.920 97.270 ;
        RECT 104.755 97.410 105.045 97.455 ;
        RECT 112.650 97.410 112.790 97.890 ;
        RECT 123.690 97.795 123.830 97.950 ;
        RECT 136.570 97.810 136.710 97.950 ;
        RECT 123.615 97.565 123.905 97.795 ;
        RECT 124.950 97.750 125.240 97.795 ;
        RECT 130.040 97.750 130.360 97.810 ;
        RECT 124.950 97.610 130.360 97.750 ;
        RECT 124.950 97.565 125.240 97.610 ;
        RECT 130.040 97.550 130.360 97.610 ;
        RECT 136.020 97.550 136.340 97.810 ;
        RECT 136.480 97.550 136.800 97.810 ;
        RECT 113.480 97.410 113.800 97.470 ;
        RECT 104.755 97.270 113.800 97.410 ;
        RECT 104.755 97.225 105.045 97.270 ;
        RECT 113.480 97.210 113.800 97.270 ;
        RECT 119.000 97.210 119.320 97.470 ;
        RECT 124.495 97.410 124.785 97.455 ;
        RECT 125.685 97.410 125.975 97.455 ;
        RECT 128.205 97.410 128.495 97.455 ;
        RECT 124.495 97.270 128.495 97.410 ;
        RECT 124.495 97.225 124.785 97.270 ;
        RECT 125.685 97.225 125.975 97.270 ;
        RECT 128.205 97.225 128.495 97.270 ;
        RECT 134.195 97.410 134.485 97.455 ;
        RECT 137.030 97.410 137.170 98.290 ;
        RECT 139.700 98.230 140.020 98.290 ;
        RECT 143.395 98.430 143.685 98.475 ;
        RECT 143.840 98.430 144.160 98.490 ;
        RECT 143.395 98.290 144.160 98.430 ;
        RECT 143.395 98.245 143.685 98.290 ;
        RECT 143.840 98.230 144.160 98.290 ;
        RECT 141.080 98.090 141.400 98.150 ;
        RECT 141.080 97.950 144.070 98.090 ;
        RECT 141.080 97.890 141.400 97.950 ;
        RECT 137.830 97.750 138.120 97.795 ;
        RECT 139.700 97.750 140.020 97.810 ;
        RECT 143.930 97.795 144.070 97.950 ;
        RECT 137.830 97.610 140.020 97.750 ;
        RECT 137.830 97.565 138.120 97.610 ;
        RECT 139.700 97.550 140.020 97.610 ;
        RECT 143.855 97.565 144.145 97.795 ;
        RECT 134.195 97.270 137.170 97.410 ;
        RECT 137.375 97.410 137.665 97.455 ;
        RECT 138.565 97.410 138.855 97.455 ;
        RECT 141.085 97.410 141.375 97.455 ;
        RECT 137.375 97.270 141.375 97.410 ;
        RECT 134.195 97.225 134.485 97.270 ;
        RECT 137.375 97.225 137.665 97.270 ;
        RECT 138.565 97.225 138.855 97.270 ;
        RECT 141.085 97.225 141.375 97.270 ;
        RECT 101.075 97.070 101.365 97.115 ;
        RECT 101.980 97.070 102.300 97.130 ;
        RECT 101.075 96.930 102.300 97.070 ;
        RECT 101.075 96.885 101.365 96.930 ;
        RECT 101.980 96.870 102.300 96.930 ;
        RECT 106.595 97.070 106.885 97.115 ;
        RECT 108.420 97.070 108.740 97.130 ;
        RECT 106.595 96.930 108.740 97.070 ;
        RECT 106.595 96.885 106.885 96.930 ;
        RECT 108.420 96.870 108.740 96.930 ;
        RECT 114.415 97.070 114.705 97.115 ;
        RECT 115.795 97.070 116.085 97.115 ;
        RECT 114.415 96.930 116.085 97.070 ;
        RECT 114.415 96.885 114.705 96.930 ;
        RECT 115.795 96.885 116.085 96.930 ;
        RECT 124.100 97.070 124.390 97.115 ;
        RECT 126.200 97.070 126.490 97.115 ;
        RECT 127.770 97.070 128.060 97.115 ;
        RECT 124.100 96.930 128.060 97.070 ;
        RECT 124.100 96.885 124.390 96.930 ;
        RECT 126.200 96.885 126.490 96.930 ;
        RECT 127.770 96.885 128.060 96.930 ;
        RECT 129.120 97.070 129.440 97.130 ;
        RECT 130.040 97.070 130.360 97.130 ;
        RECT 129.120 96.930 130.360 97.070 ;
        RECT 129.120 96.870 129.440 96.930 ;
        RECT 130.040 96.870 130.360 96.930 ;
        RECT 130.515 97.070 130.805 97.115 ;
        RECT 131.420 97.070 131.740 97.130 ;
        RECT 130.515 96.930 131.740 97.070 ;
        RECT 130.515 96.885 130.805 96.930 ;
        RECT 131.420 96.870 131.740 96.930 ;
        RECT 133.720 97.070 134.040 97.130 ;
        RECT 136.480 97.070 136.800 97.130 ;
        RECT 133.720 96.930 136.800 97.070 ;
        RECT 133.720 96.870 134.040 96.930 ;
        RECT 136.480 96.870 136.800 96.930 ;
        RECT 136.980 97.070 137.270 97.115 ;
        RECT 139.080 97.070 139.370 97.115 ;
        RECT 140.650 97.070 140.940 97.115 ;
        RECT 136.980 96.930 140.940 97.070 ;
        RECT 136.980 96.885 137.270 96.930 ;
        RECT 139.080 96.885 139.370 96.930 ;
        RECT 140.650 96.885 140.940 96.930 ;
        RECT 104.740 96.730 105.060 96.790 ;
        RECT 97.930 96.590 105.060 96.730 ;
        RECT 104.740 96.530 105.060 96.590 ;
        RECT 129.580 96.730 129.900 96.790 ;
        RECT 135.115 96.730 135.405 96.775 ;
        RECT 129.580 96.590 135.405 96.730 ;
        RECT 129.580 96.530 129.900 96.590 ;
        RECT 135.115 96.545 135.405 96.590 ;
        RECT 144.760 96.530 145.080 96.790 ;
        RECT 17.270 95.910 146.990 96.390 ;
        RECT 26.095 95.710 26.385 95.755 ;
        RECT 28.840 95.710 29.160 95.770 ;
        RECT 26.095 95.570 29.160 95.710 ;
        RECT 26.095 95.525 26.385 95.570 ;
        RECT 28.840 95.510 29.160 95.570 ;
        RECT 29.760 95.710 30.080 95.770 ;
        RECT 32.075 95.710 32.365 95.755 ;
        RECT 29.760 95.570 32.365 95.710 ;
        RECT 29.760 95.510 30.080 95.570 ;
        RECT 32.075 95.525 32.365 95.570 ;
        RECT 33.530 95.570 35.970 95.710 ;
        RECT 21.035 95.370 21.325 95.415 ;
        RECT 24.715 95.370 25.005 95.415 ;
        RECT 33.530 95.370 33.670 95.570 ;
        RECT 21.035 95.230 24.470 95.370 ;
        RECT 21.035 95.185 21.325 95.230 ;
        RECT 15.040 95.030 15.360 95.090 ;
        RECT 24.330 95.030 24.470 95.230 ;
        RECT 24.715 95.230 33.670 95.370 ;
        RECT 33.915 95.370 34.205 95.415 ;
        RECT 34.820 95.370 35.140 95.430 ;
        RECT 33.915 95.230 35.140 95.370 ;
        RECT 35.830 95.370 35.970 95.570 ;
        RECT 36.200 95.510 36.520 95.770 ;
        RECT 36.660 95.710 36.980 95.770 ;
        RECT 38.975 95.710 39.265 95.755 ;
        RECT 39.420 95.710 39.740 95.770 ;
        RECT 36.660 95.570 38.730 95.710 ;
        RECT 36.660 95.510 36.980 95.570 ;
        RECT 37.580 95.370 37.900 95.430 ;
        RECT 35.830 95.230 37.900 95.370 ;
        RECT 24.715 95.185 25.005 95.230 ;
        RECT 33.915 95.185 34.205 95.230 ;
        RECT 34.820 95.170 35.140 95.230 ;
        RECT 37.580 95.170 37.900 95.230 ;
        RECT 38.040 95.170 38.360 95.430 ;
        RECT 38.590 95.370 38.730 95.570 ;
        RECT 38.975 95.570 39.740 95.710 ;
        RECT 38.975 95.525 39.265 95.570 ;
        RECT 39.420 95.510 39.740 95.570 ;
        RECT 40.800 95.710 41.120 95.770 ;
        RECT 41.275 95.710 41.565 95.755 ;
        RECT 44.495 95.710 44.785 95.755 ;
        RECT 40.800 95.570 41.565 95.710 ;
        RECT 40.800 95.510 41.120 95.570 ;
        RECT 41.275 95.525 41.565 95.570 ;
        RECT 41.810 95.570 44.785 95.710 ;
        RECT 41.810 95.370 41.950 95.570 ;
        RECT 44.495 95.525 44.785 95.570 ;
        RECT 48.620 95.710 48.940 95.770 ;
        RECT 54.155 95.710 54.445 95.755 ;
        RECT 48.620 95.570 54.445 95.710 ;
        RECT 48.620 95.510 48.940 95.570 ;
        RECT 54.155 95.525 54.445 95.570 ;
        RECT 61.960 95.510 62.280 95.770 ;
        RECT 67.940 95.510 68.260 95.770 ;
        RECT 85.880 95.510 86.200 95.770 ;
        RECT 89.560 95.510 89.880 95.770 ;
        RECT 115.320 95.710 115.640 95.770 ;
        RECT 117.175 95.710 117.465 95.755 ;
        RECT 115.320 95.570 117.465 95.710 ;
        RECT 115.320 95.510 115.640 95.570 ;
        RECT 117.175 95.525 117.465 95.570 ;
        RECT 119.920 95.710 120.240 95.770 ;
        RECT 125.900 95.710 126.220 95.770 ;
        RECT 119.920 95.570 126.220 95.710 ;
        RECT 119.920 95.510 120.240 95.570 ;
        RECT 125.900 95.510 126.220 95.570 ;
        RECT 130.055 95.710 130.345 95.755 ;
        RECT 130.960 95.710 131.280 95.770 ;
        RECT 130.055 95.570 131.280 95.710 ;
        RECT 130.055 95.525 130.345 95.570 ;
        RECT 130.960 95.510 131.280 95.570 ;
        RECT 133.735 95.710 134.025 95.755 ;
        RECT 138.780 95.710 139.100 95.770 ;
        RECT 133.735 95.570 139.100 95.710 ;
        RECT 133.735 95.525 134.025 95.570 ;
        RECT 138.780 95.510 139.100 95.570 ;
        RECT 139.700 95.510 140.020 95.770 ;
        RECT 38.590 95.230 41.950 95.370 ;
        RECT 42.180 95.370 42.500 95.430 ;
        RECT 50.935 95.370 51.225 95.415 ;
        RECT 42.180 95.230 51.225 95.370 ;
        RECT 42.180 95.170 42.500 95.230 ;
        RECT 50.935 95.185 51.225 95.230 ;
        RECT 56.915 95.370 57.205 95.415 ;
        RECT 60.120 95.370 60.440 95.430 ;
        RECT 56.915 95.230 60.440 95.370 ;
        RECT 56.915 95.185 57.205 95.230 ;
        RECT 60.120 95.170 60.440 95.230 ;
        RECT 62.895 95.370 63.185 95.415 ;
        RECT 67.020 95.370 67.340 95.430 ;
        RECT 62.895 95.230 67.340 95.370 ;
        RECT 62.895 95.185 63.185 95.230 ;
        RECT 67.020 95.170 67.340 95.230 ;
        RECT 67.495 95.370 67.785 95.415 ;
        RECT 69.320 95.370 69.640 95.430 ;
        RECT 67.495 95.230 69.640 95.370 ;
        RECT 67.495 95.185 67.785 95.230 ;
        RECT 69.320 95.170 69.640 95.230 ;
        RECT 85.435 95.370 85.725 95.415 ;
        RECT 87.720 95.370 88.040 95.430 ;
        RECT 85.435 95.230 88.040 95.370 ;
        RECT 85.435 95.185 85.725 95.230 ;
        RECT 87.720 95.170 88.040 95.230 ;
        RECT 89.115 95.370 89.405 95.415 ;
        RECT 95.080 95.370 95.400 95.430 ;
        RECT 89.115 95.230 95.400 95.370 ;
        RECT 89.115 95.185 89.405 95.230 ;
        RECT 95.080 95.170 95.400 95.230 ;
        RECT 95.540 95.370 95.860 95.430 ;
        RECT 97.855 95.370 98.145 95.415 ;
        RECT 95.540 95.230 98.145 95.370 ;
        RECT 95.540 95.170 95.860 95.230 ;
        RECT 97.855 95.185 98.145 95.230 ;
        RECT 113.480 95.370 113.800 95.430 ;
        RECT 115.795 95.370 116.085 95.415 ;
        RECT 116.240 95.370 116.560 95.430 ;
        RECT 113.480 95.230 114.170 95.370 ;
        RECT 113.480 95.170 113.800 95.230 ;
        RECT 38.130 95.030 38.270 95.170 ;
        RECT 71.620 95.030 71.940 95.090 ;
        RECT 15.040 94.890 24.010 95.030 ;
        RECT 24.330 94.890 34.130 95.030 ;
        RECT 15.040 94.830 15.360 94.890 ;
        RECT 18.260 94.690 18.580 94.750 ;
        RECT 23.870 94.735 24.010 94.890 ;
        RECT 18.735 94.690 19.025 94.735 ;
        RECT 18.260 94.550 19.025 94.690 ;
        RECT 18.260 94.490 18.580 94.550 ;
        RECT 18.735 94.505 19.025 94.550 ;
        RECT 20.115 94.505 20.405 94.735 ;
        RECT 23.335 94.505 23.625 94.735 ;
        RECT 23.795 94.505 24.085 94.735 ;
        RECT 24.700 94.690 25.020 94.750 ;
        RECT 25.175 94.690 25.465 94.735 ;
        RECT 24.700 94.550 25.465 94.690 ;
        RECT 11.820 94.350 12.140 94.410 ;
        RECT 20.190 94.350 20.330 94.505 ;
        RECT 23.410 94.350 23.550 94.505 ;
        RECT 24.700 94.490 25.020 94.550 ;
        RECT 25.175 94.505 25.465 94.550 ;
        RECT 28.380 94.490 28.700 94.750 ;
        RECT 30.695 94.690 30.985 94.735 ;
        RECT 31.140 94.690 31.460 94.750 ;
        RECT 30.695 94.550 31.460 94.690 ;
        RECT 30.695 94.505 30.985 94.550 ;
        RECT 31.140 94.490 31.460 94.550 ;
        RECT 32.995 94.505 33.285 94.735 ;
        RECT 25.620 94.350 25.940 94.410 ;
        RECT 11.820 94.210 20.330 94.350 ;
        RECT 21.110 94.210 23.090 94.350 ;
        RECT 23.410 94.210 25.940 94.350 ;
        RECT 11.820 94.150 12.140 94.210 ;
        RECT 19.655 94.010 19.945 94.055 ;
        RECT 21.110 94.010 21.250 94.210 ;
        RECT 19.655 93.870 21.250 94.010 ;
        RECT 21.480 94.010 21.800 94.070 ;
        RECT 22.415 94.010 22.705 94.055 ;
        RECT 21.480 93.870 22.705 94.010 ;
        RECT 22.950 94.010 23.090 94.210 ;
        RECT 25.620 94.150 25.940 94.210 ;
        RECT 27.460 94.350 27.780 94.410 ;
        RECT 33.070 94.350 33.210 94.505 ;
        RECT 33.440 94.490 33.760 94.750 ;
        RECT 27.460 94.210 33.210 94.350 ;
        RECT 33.990 94.350 34.130 94.890 ;
        RECT 34.450 94.890 38.270 95.030 ;
        RECT 59.750 94.890 71.940 95.030 ;
        RECT 34.450 94.735 34.590 94.890 ;
        RECT 34.375 94.505 34.665 94.735 ;
        RECT 34.820 94.690 35.140 94.750 ;
        RECT 35.295 94.690 35.585 94.735 ;
        RECT 34.820 94.550 35.585 94.690 ;
        RECT 34.820 94.490 35.140 94.550 ;
        RECT 35.295 94.505 35.585 94.550 ;
        RECT 38.040 94.490 38.360 94.750 ;
        RECT 40.800 94.690 41.120 94.750 ;
        RECT 42.195 94.690 42.485 94.735 ;
        RECT 40.800 94.550 42.485 94.690 ;
        RECT 40.800 94.490 41.120 94.550 ;
        RECT 42.195 94.505 42.485 94.550 ;
        RECT 44.020 94.690 44.340 94.750 ;
        RECT 45.415 94.690 45.705 94.735 ;
        RECT 44.020 94.550 45.705 94.690 ;
        RECT 44.020 94.490 44.340 94.550 ;
        RECT 45.415 94.505 45.705 94.550 ;
        RECT 47.240 94.690 47.560 94.750 ;
        RECT 48.635 94.690 48.925 94.735 ;
        RECT 47.240 94.550 48.925 94.690 ;
        RECT 47.240 94.490 47.560 94.550 ;
        RECT 48.635 94.505 48.925 94.550 ;
        RECT 50.460 94.690 50.780 94.750 ;
        RECT 51.855 94.690 52.145 94.735 ;
        RECT 50.460 94.550 52.145 94.690 ;
        RECT 50.460 94.490 50.780 94.550 ;
        RECT 51.855 94.505 52.145 94.550 ;
        RECT 53.680 94.690 54.000 94.750 ;
        RECT 55.075 94.690 55.365 94.735 ;
        RECT 53.680 94.550 55.365 94.690 ;
        RECT 53.680 94.490 54.000 94.550 ;
        RECT 55.075 94.505 55.365 94.550 ;
        RECT 57.820 94.490 58.140 94.750 ;
        RECT 59.750 94.735 59.890 94.890 ;
        RECT 71.620 94.830 71.940 94.890 ;
        RECT 72.540 94.830 72.860 95.090 ;
        RECT 83.595 95.030 83.885 95.075 ;
        RECT 86.800 95.030 87.120 95.090 ;
        RECT 83.595 94.890 87.120 95.030 ;
        RECT 83.595 94.845 83.885 94.890 ;
        RECT 86.800 94.830 87.120 94.890 ;
        RECT 87.260 95.030 87.580 95.090 ;
        RECT 114.030 95.075 114.170 95.230 ;
        RECT 115.795 95.230 116.560 95.370 ;
        RECT 115.795 95.185 116.085 95.230 ;
        RECT 116.240 95.170 116.560 95.230 ;
        RECT 118.080 95.370 118.400 95.430 ;
        RECT 123.615 95.370 123.905 95.415 ;
        RECT 118.080 95.230 123.905 95.370 ;
        RECT 118.080 95.170 118.400 95.230 ;
        RECT 123.615 95.185 123.905 95.230 ;
        RECT 124.980 95.370 125.300 95.430 ;
        RECT 131.435 95.370 131.725 95.415 ;
        RECT 137.400 95.370 137.720 95.430 ;
        RECT 124.980 95.230 131.725 95.370 ;
        RECT 124.980 95.170 125.300 95.230 ;
        RECT 131.435 95.185 131.725 95.230 ;
        RECT 137.085 95.230 137.720 95.370 ;
        RECT 87.260 94.890 91.630 95.030 ;
        RECT 87.260 94.830 87.580 94.890 ;
        RECT 59.675 94.505 59.965 94.735 ;
        RECT 61.515 94.690 61.805 94.735 ;
        RECT 67.480 94.690 67.800 94.750 ;
        RECT 61.515 94.550 67.800 94.690 ;
        RECT 61.515 94.505 61.805 94.550 ;
        RECT 67.480 94.490 67.800 94.550 ;
        RECT 71.160 94.490 71.480 94.750 ;
        RECT 73.460 94.490 73.780 94.750 ;
        RECT 77.600 94.490 77.920 94.750 ;
        RECT 78.060 94.490 78.380 94.750 ;
        RECT 79.900 94.490 80.220 94.750 ;
        RECT 45.860 94.350 46.180 94.410 ;
        RECT 63.340 94.350 63.660 94.410 ;
        RECT 33.990 94.210 46.180 94.350 ;
        RECT 27.460 94.150 27.780 94.210 ;
        RECT 45.860 94.150 46.180 94.210 ;
        RECT 58.830 94.210 63.660 94.350 ;
        RECT 27.550 94.010 27.690 94.150 ;
        RECT 22.950 93.870 27.690 94.010 ;
        RECT 27.920 94.010 28.240 94.070 ;
        RECT 29.315 94.010 29.605 94.055 ;
        RECT 27.920 93.870 29.605 94.010 ;
        RECT 19.655 93.825 19.945 93.870 ;
        RECT 21.480 93.810 21.800 93.870 ;
        RECT 22.415 93.825 22.705 93.870 ;
        RECT 27.920 93.810 28.240 93.870 ;
        RECT 29.315 93.825 29.605 93.870 ;
        RECT 31.615 94.010 31.905 94.055 ;
        RECT 38.960 94.010 39.280 94.070 ;
        RECT 31.615 93.870 39.280 94.010 ;
        RECT 31.615 93.825 31.905 93.870 ;
        RECT 38.960 93.810 39.280 93.870 ;
        RECT 47.700 93.810 48.020 94.070 ;
        RECT 58.830 94.055 58.970 94.210 ;
        RECT 63.340 94.150 63.660 94.210 ;
        RECT 64.275 94.350 64.565 94.395 ;
        RECT 64.720 94.350 65.040 94.410 ;
        RECT 65.655 94.350 65.945 94.395 ;
        RECT 64.275 94.210 65.945 94.350 ;
        RECT 64.275 94.165 64.565 94.210 ;
        RECT 64.720 94.150 65.040 94.210 ;
        RECT 65.655 94.165 65.945 94.210 ;
        RECT 66.100 94.350 66.420 94.410 ;
        RECT 86.890 94.350 87.030 94.830 ;
        RECT 91.490 94.735 91.630 94.890 ;
        RECT 113.955 94.845 114.245 95.075 ;
        RECT 118.540 95.030 118.860 95.090 ;
        RECT 124.520 95.030 124.840 95.090 ;
        RECT 126.835 95.030 127.125 95.075 ;
        RECT 118.540 94.890 122.220 95.030 ;
        RECT 118.540 94.830 118.860 94.890 ;
        RECT 91.415 94.505 91.705 94.735 ;
        RECT 91.860 94.490 92.180 94.750 ;
        RECT 94.160 94.690 94.480 94.750 ;
        RECT 95.095 94.690 95.385 94.735 ;
        RECT 94.160 94.550 95.385 94.690 ;
        RECT 94.160 94.490 94.480 94.550 ;
        RECT 95.095 94.505 95.385 94.550 ;
        RECT 96.935 94.690 97.225 94.735 ;
        RECT 97.380 94.690 97.700 94.750 ;
        RECT 96.935 94.550 97.700 94.690 ;
        RECT 96.935 94.505 97.225 94.550 ;
        RECT 97.380 94.490 97.700 94.550 ;
        RECT 100.615 94.690 100.905 94.735 ;
        RECT 102.900 94.690 103.220 94.750 ;
        RECT 100.615 94.550 103.220 94.690 ;
        RECT 100.615 94.505 100.905 94.550 ;
        RECT 102.900 94.490 103.220 94.550 ;
        RECT 103.835 94.690 104.125 94.735 ;
        RECT 104.280 94.690 104.600 94.750 ;
        RECT 103.835 94.550 104.600 94.690 ;
        RECT 103.835 94.505 104.125 94.550 ;
        RECT 104.280 94.490 104.600 94.550 ;
        RECT 107.055 94.690 107.345 94.735 ;
        RECT 107.960 94.690 108.280 94.750 ;
        RECT 107.055 94.550 108.280 94.690 ;
        RECT 107.055 94.505 107.345 94.550 ;
        RECT 107.960 94.490 108.280 94.550 ;
        RECT 110.275 94.690 110.565 94.735 ;
        RECT 111.180 94.690 111.500 94.750 ;
        RECT 110.275 94.550 111.500 94.690 ;
        RECT 110.275 94.505 110.565 94.550 ;
        RECT 111.180 94.490 111.500 94.550 ;
        RECT 113.020 94.690 113.340 94.750 ;
        RECT 113.495 94.690 113.785 94.735 ;
        RECT 113.020 94.550 113.785 94.690 ;
        RECT 113.020 94.490 113.340 94.550 ;
        RECT 113.495 94.505 113.785 94.550 ;
        RECT 118.095 94.690 118.385 94.735 ;
        RECT 119.460 94.690 119.780 94.750 ;
        RECT 118.095 94.550 119.780 94.690 ;
        RECT 118.095 94.505 118.385 94.550 ;
        RECT 119.460 94.490 119.780 94.550 ;
        RECT 119.920 94.490 120.240 94.750 ;
        RECT 120.840 94.490 121.160 94.750 ;
        RECT 122.080 94.690 122.220 94.890 ;
        RECT 124.520 94.890 127.125 95.030 ;
        RECT 124.520 94.830 124.840 94.890 ;
        RECT 126.835 94.845 127.125 94.890 ;
        RECT 127.755 95.030 128.045 95.075 ;
        RECT 130.960 95.030 131.280 95.090 ;
        RECT 127.755 94.890 131.280 95.030 ;
        RECT 127.755 94.845 128.045 94.890 ;
        RECT 130.960 94.830 131.280 94.890 ;
        RECT 122.695 94.690 122.985 94.735 ;
        RECT 122.080 94.550 122.985 94.690 ;
        RECT 122.695 94.505 122.985 94.550 ;
        RECT 125.900 94.490 126.220 94.750 ;
        RECT 130.500 94.490 130.820 94.750 ;
        RECT 132.340 94.690 132.660 94.750 ;
        RECT 134.425 94.690 134.715 94.735 ;
        RECT 132.340 94.550 134.715 94.690 ;
        RECT 132.340 94.490 132.660 94.550 ;
        RECT 134.425 94.505 134.715 94.550 ;
        RECT 135.100 94.490 135.420 94.750 ;
        RECT 135.560 94.490 135.880 94.750 ;
        RECT 136.480 94.690 136.800 94.750 ;
        RECT 137.085 94.735 137.225 95.230 ;
        RECT 137.400 95.170 137.720 95.230 ;
        RECT 139.255 95.370 139.545 95.415 ;
        RECT 141.540 95.370 141.860 95.430 ;
        RECT 139.255 95.230 141.860 95.370 ;
        RECT 139.255 95.185 139.545 95.230 ;
        RECT 141.540 95.170 141.860 95.230 ;
        RECT 144.775 95.185 145.065 95.415 ;
        RECT 138.320 95.030 138.640 95.090 ;
        RECT 144.850 95.030 144.990 95.185 ;
        RECT 138.320 94.890 144.990 95.030 ;
        RECT 138.320 94.830 138.640 94.890 ;
        RECT 136.285 94.550 136.800 94.690 ;
        RECT 136.480 94.490 136.800 94.550 ;
        RECT 136.955 94.505 137.245 94.735 ;
        RECT 137.400 94.490 137.720 94.750 ;
        RECT 140.160 94.490 140.480 94.750 ;
        RECT 142.000 94.490 142.320 94.750 ;
        RECT 142.920 94.690 143.240 94.750 ;
        RECT 143.855 94.690 144.145 94.735 ;
        RECT 142.920 94.550 144.145 94.690 ;
        RECT 142.920 94.490 143.240 94.550 ;
        RECT 143.855 94.505 144.145 94.550 ;
        RECT 87.275 94.350 87.565 94.395 ;
        RECT 66.100 94.210 69.550 94.350 ;
        RECT 86.890 94.210 87.565 94.350 ;
        RECT 66.100 94.150 66.420 94.210 ;
        RECT 58.755 93.825 59.045 94.055 ;
        RECT 60.595 94.010 60.885 94.055 ;
        RECT 66.560 94.010 66.880 94.070 ;
        RECT 69.410 94.055 69.550 94.210 ;
        RECT 87.275 94.165 87.565 94.210 ;
        RECT 89.100 94.350 89.420 94.410 ;
        RECT 92.320 94.350 92.640 94.410 ;
        RECT 114.860 94.350 115.180 94.410 ;
        RECT 89.100 94.210 91.170 94.350 ;
        RECT 89.100 94.150 89.420 94.210 ;
        RECT 60.595 93.870 66.880 94.010 ;
        RECT 60.595 93.825 60.885 93.870 ;
        RECT 66.560 93.810 66.880 93.870 ;
        RECT 69.335 93.825 69.625 94.055 ;
        RECT 73.000 94.010 73.320 94.070 ;
        RECT 74.395 94.010 74.685 94.055 ;
        RECT 73.000 93.870 74.685 94.010 ;
        RECT 73.000 93.810 73.320 93.870 ;
        RECT 74.395 93.825 74.685 93.870 ;
        RECT 76.220 94.010 76.540 94.070 ;
        RECT 76.695 94.010 76.985 94.055 ;
        RECT 76.220 93.870 76.985 94.010 ;
        RECT 76.220 93.810 76.540 93.870 ;
        RECT 76.695 93.825 76.985 93.870 ;
        RECT 78.995 94.010 79.285 94.055 ;
        RECT 79.440 94.010 79.760 94.070 ;
        RECT 78.995 93.870 79.760 94.010 ;
        RECT 78.995 93.825 79.285 93.870 ;
        RECT 79.440 93.810 79.760 93.870 ;
        RECT 80.835 94.010 81.125 94.055 ;
        RECT 82.660 94.010 82.980 94.070 ;
        RECT 80.835 93.870 82.980 94.010 ;
        RECT 80.835 93.825 81.125 93.870 ;
        RECT 82.660 93.810 82.980 93.870 ;
        RECT 85.880 94.010 86.200 94.070 ;
        RECT 90.495 94.010 90.785 94.055 ;
        RECT 85.880 93.870 90.785 94.010 ;
        RECT 91.030 94.010 91.170 94.210 ;
        RECT 92.320 94.210 94.620 94.350 ;
        RECT 92.320 94.150 92.640 94.210 ;
        RECT 92.795 94.010 93.085 94.055 ;
        RECT 91.030 93.870 93.085 94.010 ;
        RECT 94.480 94.010 94.620 94.210 ;
        RECT 114.860 94.210 117.850 94.350 ;
        RECT 114.860 94.150 115.180 94.210 ;
        RECT 96.015 94.010 96.305 94.055 ;
        RECT 94.480 93.870 96.305 94.010 ;
        RECT 85.880 93.810 86.200 93.870 ;
        RECT 90.495 93.825 90.785 93.870 ;
        RECT 92.795 93.825 93.085 93.870 ;
        RECT 96.015 93.825 96.305 93.870 ;
        RECT 98.760 94.010 99.080 94.070 ;
        RECT 99.695 94.010 99.985 94.055 ;
        RECT 98.760 93.870 99.985 94.010 ;
        RECT 98.760 93.810 99.080 93.870 ;
        RECT 99.695 93.825 99.985 93.870 ;
        RECT 101.980 94.010 102.300 94.070 ;
        RECT 102.915 94.010 103.205 94.055 ;
        RECT 101.980 93.870 103.205 94.010 ;
        RECT 101.980 93.810 102.300 93.870 ;
        RECT 102.915 93.825 103.205 93.870 ;
        RECT 105.200 94.010 105.520 94.070 ;
        RECT 106.135 94.010 106.425 94.055 ;
        RECT 105.200 93.870 106.425 94.010 ;
        RECT 105.200 93.810 105.520 93.870 ;
        RECT 106.135 93.825 106.425 93.870 ;
        RECT 108.420 94.010 108.740 94.070 ;
        RECT 109.355 94.010 109.645 94.055 ;
        RECT 108.420 93.870 109.645 94.010 ;
        RECT 108.420 93.810 108.740 93.870 ;
        RECT 109.355 93.825 109.645 93.870 ;
        RECT 111.640 94.010 111.960 94.070 ;
        RECT 112.575 94.010 112.865 94.055 ;
        RECT 111.640 93.870 112.865 94.010 ;
        RECT 111.640 93.810 111.960 93.870 ;
        RECT 112.575 93.825 112.865 93.870 ;
        RECT 116.240 93.810 116.560 94.070 ;
        RECT 117.710 94.010 117.850 94.210 ;
        RECT 118.540 94.150 118.860 94.410 ;
        RECT 119.000 94.150 119.320 94.410 ;
        RECT 121.300 94.350 121.620 94.410 ;
        RECT 130.960 94.350 131.280 94.410 ;
        RECT 121.300 94.210 125.210 94.350 ;
        RECT 121.300 94.150 121.620 94.210 ;
        RECT 125.070 94.055 125.210 94.210 ;
        RECT 130.960 94.210 134.410 94.350 ;
        RECT 130.960 94.150 131.280 94.210 ;
        RECT 121.775 94.010 122.065 94.055 ;
        RECT 117.710 93.870 122.065 94.010 ;
        RECT 121.775 93.825 122.065 93.870 ;
        RECT 124.995 93.825 125.285 94.055 ;
        RECT 128.215 94.010 128.505 94.055 ;
        RECT 132.800 94.010 133.120 94.070 ;
        RECT 128.215 93.870 133.120 94.010 ;
        RECT 134.270 94.010 134.410 94.210 ;
        RECT 141.095 94.010 141.385 94.055 ;
        RECT 134.270 93.870 141.385 94.010 ;
        RECT 128.215 93.825 128.505 93.870 ;
        RECT 132.800 93.810 133.120 93.870 ;
        RECT 141.095 93.825 141.385 93.870 ;
        RECT 142.920 93.810 143.240 94.070 ;
        RECT 17.270 93.190 146.990 93.670 ;
        RECT 33.440 92.990 33.760 93.050 ;
        RECT 47.700 92.990 48.020 93.050 ;
        RECT 13.660 92.890 13.980 92.950 ;
        RECT 27.950 92.890 28.210 92.980 ;
        RECT 13.660 92.750 28.210 92.890 ;
        RECT 33.440 92.850 48.020 92.990 ;
        RECT 33.440 92.790 33.760 92.850 ;
        RECT 47.700 92.790 48.020 92.850 ;
        RECT 57.820 92.990 58.140 93.050 ;
        RECT 68.860 92.990 69.180 93.050 ;
        RECT 57.820 92.850 69.180 92.990 ;
        RECT 57.820 92.790 58.140 92.850 ;
        RECT 68.860 92.790 69.180 92.850 ;
        RECT 116.240 92.990 116.560 93.050 ;
        RECT 124.060 92.990 124.380 93.050 ;
        RECT 116.240 92.850 124.380 92.990 ;
        RECT 116.240 92.790 116.560 92.850 ;
        RECT 124.060 92.790 124.380 92.850 ;
        RECT 13.660 92.690 13.980 92.750 ;
        RECT 27.950 92.660 28.210 92.750 ;
        RECT 104.740 92.650 105.060 92.710 ;
        RECT 119.000 92.650 119.320 92.710 ;
        RECT 135.560 92.650 135.880 92.710 ;
        RECT 104.740 92.510 135.880 92.650 ;
        RECT 104.740 92.450 105.060 92.510 ;
        RECT 119.000 92.450 119.320 92.510 ;
        RECT 135.560 92.450 135.880 92.510 ;
        RECT 12.910 92.250 13.330 92.390 ;
        RECT 21.470 92.250 21.810 92.350 ;
        RECT 12.910 92.110 21.810 92.250 ;
        RECT 12.910 91.970 13.330 92.110 ;
        RECT 21.470 92.020 21.810 92.110 ;
        RECT 147.310 89.460 147.450 104.080 ;
        RECT 147.590 104.020 147.910 104.080 ;
        RECT 136.120 89.320 147.450 89.460 ;
        RECT 136.120 89.310 136.440 89.320 ;
        RECT 127.740 89.250 128.060 89.310 ;
        RECT 136.020 89.250 136.440 89.310 ;
        RECT 127.740 89.190 136.440 89.250 ;
        RECT 127.740 89.110 136.340 89.190 ;
        RECT 127.740 89.050 128.060 89.110 ;
        RECT 136.020 89.050 136.340 89.110 ;
        RECT 140.620 88.910 140.940 88.970 ;
        RECT 144.760 88.910 145.080 88.970 ;
        RECT 140.620 88.770 145.080 88.910 ;
        RECT 140.620 88.710 140.940 88.770 ;
        RECT 144.760 88.710 145.080 88.770 ;
        RECT 134.180 88.230 134.500 88.290 ;
        RECT 142.920 88.230 143.240 88.290 ;
        RECT 134.180 88.090 143.240 88.230 ;
        RECT 134.180 88.030 134.500 88.090 ;
        RECT 142.920 88.030 143.240 88.090 ;
        RECT 147.540 85.605 147.860 85.660 ;
        RECT 147.445 85.400 147.860 85.605 ;
        RECT 56.880 83.580 57.250 83.660 ;
        RECT 53.165 83.365 57.250 83.580 ;
        RECT 37.570 82.630 37.910 82.910 ;
        RECT 37.600 81.080 37.880 82.630 ;
        RECT 53.165 77.640 53.380 83.365 ;
        RECT 56.880 83.290 57.250 83.365 ;
        RECT 53.700 80.740 53.980 82.960 ;
        RECT 53.035 77.425 53.380 77.640 ;
        RECT 53.035 28.890 53.250 77.425 ;
        RECT 53.735 76.915 53.945 80.740 ;
        RECT 147.445 77.640 147.595 85.400 ;
        RECT 147.965 85.025 148.225 85.095 ;
        RECT 147.855 84.775 148.225 85.025 ;
        RECT 147.855 79.425 148.030 84.775 ;
        RECT 148.480 84.395 148.800 84.420 ;
        RECT 148.325 84.160 148.800 84.395 ;
        RECT 148.325 80.020 148.535 84.160 ;
        RECT 148.820 80.510 149.080 83.720 ;
        RECT 149.440 82.670 149.700 82.990 ;
        RECT 149.470 81.060 149.670 82.670 ;
        RECT 149.440 80.740 149.700 81.060 ;
        RECT 148.790 80.250 149.110 80.510 ;
        RECT 148.300 79.700 148.560 80.020 ;
        RECT 147.815 79.105 148.075 79.425 ;
        RECT 151.810 78.185 152.045 174.575 ;
        RECT 152.430 142.270 152.750 142.530 ;
        RECT 152.475 78.860 152.705 142.270 ;
        RECT 152.460 78.540 152.720 78.860 ;
        RECT 151.800 77.865 152.060 78.185 ;
        RECT 147.390 77.320 147.650 77.640 ;
        RECT 53.625 76.705 53.945 76.915 ;
        RECT 53.625 29.275 53.835 76.705 ;
        RECT 73.730 76.490 75.490 76.500 ;
        RECT 73.730 76.470 90.620 76.490 ;
        RECT 102.030 76.470 105.400 76.480 ;
        RECT 68.260 76.415 68.580 76.470 ;
        RECT 54.055 76.265 68.580 76.415 ;
        RECT 54.055 29.655 54.205 76.265 ;
        RECT 68.260 76.210 68.580 76.265 ;
        RECT 73.730 76.420 117.930 76.470 ;
        RECT 120.090 76.460 132.940 76.470 ;
        RECT 135.080 76.460 147.930 76.470 ;
        RECT 120.090 76.420 147.930 76.460 ;
        RECT 73.730 76.340 147.930 76.420 ;
        RECT 73.730 76.040 147.960 76.340 ;
        RECT 54.680 76.020 147.960 76.040 ;
        RECT 54.660 75.570 147.960 76.020 ;
        RECT 54.660 75.530 88.580 75.570 ;
        RECT 54.660 75.210 74.080 75.530 ;
        RECT 54.680 75.170 74.080 75.210 ;
        RECT 75.900 75.170 76.860 75.200 ;
        RECT 54.680 75.150 67.490 75.170 ;
        RECT 55.680 74.790 56.120 75.150 ;
        RECT 57.260 75.040 58.420 75.150 ;
        RECT 57.260 74.790 57.700 75.040 ;
        RECT 58.850 74.790 59.290 75.150 ;
        RECT 60.440 74.790 60.880 75.150 ;
        RECT 54.820 74.740 55.050 74.770 ;
        RECT 55.210 74.740 55.440 74.790 ;
        RECT 54.820 68.850 55.440 74.740 ;
        RECT 54.820 68.570 55.060 68.850 ;
        RECT 55.210 68.790 55.440 68.850 ;
        RECT 55.650 68.850 56.120 74.790 ;
        RECT 56.790 74.720 57.020 74.790 ;
        RECT 56.490 68.870 57.020 74.720 ;
        RECT 56.490 68.850 56.650 68.870 ;
        RECT 55.650 68.790 55.880 68.850 ;
        RECT 56.500 68.610 56.650 68.850 ;
        RECT 56.790 68.790 57.020 68.870 ;
        RECT 57.230 68.870 57.700 74.790 ;
        RECT 58.370 74.720 58.600 74.790 ;
        RECT 58.000 70.130 58.610 74.720 ;
        RECT 57.230 68.790 57.460 68.870 ;
        RECT 57.980 68.840 58.610 70.130 ;
        RECT 58.810 68.880 59.290 74.790 ;
        RECT 59.950 74.740 60.180 74.790 ;
        RECT 54.820 66.140 55.200 68.570 ;
        RECT 55.400 68.560 55.690 68.585 ;
        RECT 55.390 67.830 55.710 68.560 ;
        RECT 55.340 66.830 56.340 67.830 ;
        RECT 55.390 66.140 55.710 66.830 ;
        RECT 54.820 65.830 55.060 66.140 ;
        RECT 55.410 66.100 55.710 66.140 ;
        RECT 55.410 66.090 55.700 66.100 ;
        RECT 56.500 66.080 56.700 68.610 ;
        RECT 56.980 68.580 57.270 68.585 ;
        RECT 56.970 67.880 57.310 68.580 ;
        RECT 56.840 66.880 57.840 67.880 ;
        RECT 56.970 66.110 57.310 66.880 ;
        RECT 56.990 66.090 57.280 66.110 ;
        RECT 55.220 65.830 55.450 65.930 ;
        RECT 54.820 65.820 55.450 65.830 ;
        RECT 54.790 64.020 55.450 65.820 ;
        RECT 54.820 64.000 55.050 64.020 ;
        RECT 55.220 63.930 55.450 64.020 ;
        RECT 55.660 65.860 55.890 65.930 ;
        RECT 55.660 64.050 56.220 65.860 ;
        RECT 56.500 65.820 56.650 66.080 ;
        RECT 56.800 65.820 57.030 65.930 ;
        RECT 56.500 65.810 57.030 65.820 ;
        RECT 55.660 63.930 55.890 64.050 ;
        RECT 56.050 63.730 56.220 64.050 ;
        RECT 56.460 64.010 57.030 65.810 ;
        RECT 56.510 64.000 57.030 64.010 ;
        RECT 56.800 63.930 57.030 64.000 ;
        RECT 57.240 65.880 57.470 65.930 ;
        RECT 57.240 65.850 57.750 65.880 ;
        RECT 57.240 64.040 57.780 65.850 ;
        RECT 57.980 65.830 58.170 68.840 ;
        RECT 58.370 68.790 58.600 68.840 ;
        RECT 58.810 68.790 59.040 68.880 ;
        RECT 59.560 68.840 60.180 74.740 ;
        RECT 58.530 67.880 58.890 68.590 ;
        RECT 58.350 66.880 59.350 67.880 ;
        RECT 58.530 66.090 58.890 66.880 ;
        RECT 58.380 65.830 58.610 65.930 ;
        RECT 57.980 65.160 58.610 65.830 ;
        RECT 57.240 63.930 57.470 64.040 ;
        RECT 57.610 63.810 57.780 64.040 ;
        RECT 58.000 63.960 58.610 65.160 ;
        RECT 58.380 63.930 58.610 63.960 ;
        RECT 58.820 65.880 59.050 65.930 ;
        RECT 58.820 64.000 59.360 65.880 ;
        RECT 59.580 65.860 59.750 68.840 ;
        RECT 59.950 68.790 60.180 68.840 ;
        RECT 60.390 68.870 60.880 74.790 ;
        RECT 61.530 74.710 61.760 74.790 ;
        RECT 60.390 68.790 60.620 68.870 ;
        RECT 61.120 68.830 61.760 74.710 ;
        RECT 60.140 68.580 60.430 68.585 ;
        RECT 60.130 67.910 60.470 68.580 ;
        RECT 59.960 66.910 60.960 67.910 ;
        RECT 60.130 66.100 60.470 66.910 ;
        RECT 60.150 66.090 60.440 66.100 ;
        RECT 59.960 65.860 60.190 65.930 ;
        RECT 59.580 65.820 60.190 65.860 ;
        RECT 59.560 64.020 60.190 65.820 ;
        RECT 59.590 64.000 60.190 64.020 ;
        RECT 58.820 63.930 59.050 64.000 ;
        RECT 54.690 63.590 55.690 63.600 ;
        RECT 55.970 63.590 56.220 63.730 ;
        RECT 57.600 63.590 57.780 63.810 ;
        RECT 59.190 63.760 59.360 64.000 ;
        RECT 59.960 63.930 60.190 64.000 ;
        RECT 60.400 65.860 60.630 65.930 ;
        RECT 60.400 63.980 60.940 65.860 ;
        RECT 61.130 65.850 61.320 68.830 ;
        RECT 61.530 68.790 61.760 68.830 ;
        RECT 61.960 68.820 62.400 75.150 ;
        RECT 63.580 74.790 64.020 75.150 ;
        RECT 65.170 74.790 65.610 75.150 ;
        RECT 66.750 74.790 67.190 75.150 ;
        RECT 63.110 74.770 63.340 74.790 ;
        RECT 62.660 68.840 63.340 74.770 ;
        RECT 61.970 68.790 62.200 68.820 ;
        RECT 61.720 68.580 62.010 68.585 ;
        RECT 61.700 67.880 62.060 68.580 ;
        RECT 61.510 66.880 62.510 67.880 ;
        RECT 61.700 66.090 62.060 66.880 ;
        RECT 61.540 65.850 61.770 65.930 ;
        RECT 61.130 64.000 61.770 65.850 ;
        RECT 60.400 63.930 60.630 63.980 ;
        RECT 59.180 63.590 59.360 63.760 ;
        RECT 60.770 63.590 60.940 63.980 ;
        RECT 61.540 63.930 61.770 64.000 ;
        RECT 61.980 65.880 62.210 65.930 ;
        RECT 62.670 65.890 62.930 68.840 ;
        RECT 63.110 68.790 63.340 68.840 ;
        RECT 63.550 68.850 64.020 74.790 ;
        RECT 64.690 74.750 64.920 74.790 ;
        RECT 63.550 68.790 63.780 68.850 ;
        RECT 64.240 68.840 64.920 74.750 ;
        RECT 63.300 68.580 63.590 68.585 ;
        RECT 63.270 67.910 63.610 68.580 ;
        RECT 63.130 66.910 64.130 67.910 ;
        RECT 63.270 66.090 63.610 66.910 ;
        RECT 63.120 65.890 63.350 65.930 ;
        RECT 61.980 64.000 62.520 65.880 ;
        RECT 61.980 63.930 62.210 64.000 ;
        RECT 62.350 63.590 62.520 64.000 ;
        RECT 62.670 63.970 63.350 65.890 ;
        RECT 63.120 63.930 63.350 63.970 ;
        RECT 63.560 65.870 63.790 65.930 ;
        RECT 63.560 63.990 64.110 65.870 ;
        RECT 64.290 65.850 64.550 68.840 ;
        RECT 64.690 68.790 64.920 68.840 ;
        RECT 65.130 68.830 65.610 74.790 ;
        RECT 66.270 74.750 66.500 74.790 ;
        RECT 65.840 68.860 66.500 74.750 ;
        RECT 65.840 68.840 66.100 68.860 ;
        RECT 65.130 68.790 65.360 68.830 ;
        RECT 65.850 68.630 66.100 68.840 ;
        RECT 66.270 68.790 66.500 68.860 ;
        RECT 66.710 68.880 67.190 74.790 ;
        RECT 73.740 73.530 74.080 75.170 ;
        RECT 75.570 74.970 76.860 75.170 ;
        RECT 75.570 74.730 76.630 74.970 ;
        RECT 77.130 74.765 77.350 75.530 ;
        RECT 82.340 75.200 83.310 75.230 ;
        RECT 78.330 74.970 80.290 75.200 ;
        RECT 81.760 74.970 83.720 75.200 ;
        RECT 85.190 74.970 86.150 75.200 ;
        RECT 73.720 71.890 74.070 72.970 ;
        RECT 73.550 71.030 74.260 71.890 ;
        RECT 66.710 68.790 66.940 68.880 ;
        RECT 64.880 68.580 65.170 68.585 ;
        RECT 64.870 67.880 65.200 68.580 ;
        RECT 64.700 66.880 65.700 67.880 ;
        RECT 64.870 66.090 65.200 66.880 ;
        RECT 65.850 66.530 66.150 68.630 ;
        RECT 66.460 68.580 66.750 68.585 ;
        RECT 66.440 67.900 66.800 68.580 ;
        RECT 66.360 66.900 67.360 67.900 ;
        RECT 73.720 67.540 74.070 71.030 ;
        RECT 75.520 67.620 76.630 74.730 ;
        RECT 65.930 66.080 66.150 66.530 ;
        RECT 66.440 66.090 66.800 66.900 ;
        RECT 73.720 66.540 74.060 66.970 ;
        RECT 75.510 66.560 76.630 67.620 ;
        RECT 76.910 74.560 77.350 74.765 ;
        RECT 78.050 74.740 78.280 74.765 ;
        RECT 78.050 74.730 78.290 74.740 ;
        RECT 76.910 66.820 77.300 74.560 ;
        RECT 77.880 67.670 78.290 74.730 ;
        RECT 78.870 68.380 79.770 74.970 ;
        RECT 80.340 74.720 80.570 74.765 ;
        RECT 81.480 74.740 81.710 74.765 ;
        RECT 77.870 66.850 78.290 67.670 ;
        RECT 78.840 67.370 79.840 68.380 ;
        RECT 76.910 66.765 77.140 66.820 ;
        RECT 77.870 66.765 78.280 66.850 ;
        RECT 64.700 65.850 64.930 65.930 ;
        RECT 64.270 64.000 64.930 65.850 ;
        RECT 63.560 63.930 63.790 63.990 ;
        RECT 63.950 63.590 64.110 63.990 ;
        RECT 64.700 63.930 64.930 64.000 ;
        RECT 65.140 65.870 65.370 65.930 ;
        RECT 65.140 63.980 65.690 65.870 ;
        RECT 65.930 65.840 66.110 66.080 ;
        RECT 66.280 65.840 66.510 65.930 ;
        RECT 65.930 65.690 66.510 65.840 ;
        RECT 65.900 64.020 66.510 65.690 ;
        RECT 65.910 63.990 66.510 64.020 ;
        RECT 65.140 63.930 65.370 63.980 ;
        RECT 65.520 63.590 65.690 63.980 ;
        RECT 66.280 63.930 66.510 63.990 ;
        RECT 66.720 65.870 66.950 65.930 ;
        RECT 66.720 64.020 67.410 65.870 ;
        RECT 73.390 65.430 74.340 66.540 ;
        RECT 75.510 66.330 76.860 66.560 ;
        RECT 75.510 65.690 76.720 66.330 ;
        RECT 66.720 63.930 66.950 64.020 ;
        RECT 67.100 63.770 67.410 64.020 ;
        RECT 67.080 63.730 67.410 63.770 ;
        RECT 67.080 63.590 67.570 63.730 ;
        RECT 54.690 63.560 67.570 63.590 ;
        RECT 54.670 62.570 67.570 63.560 ;
        RECT 54.690 62.530 67.570 62.570 ;
        RECT 55.230 59.850 55.840 62.190 ;
        RECT 56.670 62.000 57.330 62.320 ;
        RECT 56.720 59.880 57.330 62.000 ;
        RECT 57.170 59.850 57.330 59.880 ;
        RECT 58.190 59.840 58.740 62.190 ;
        RECT 59.700 59.820 60.250 62.170 ;
        RECT 61.160 59.850 61.710 62.200 ;
        RECT 62.640 59.880 63.190 62.230 ;
        RECT 64.090 59.870 64.640 62.220 ;
        RECT 65.590 59.880 66.140 62.230 ;
        RECT 67.010 62.090 67.570 62.530 ;
        RECT 67.010 59.930 67.580 62.090 ;
        RECT 73.720 61.550 74.060 65.430 ;
        RECT 75.070 64.440 76.720 65.690 ;
        RECT 67.010 59.920 67.570 59.930 ;
        RECT 73.730 59.570 74.070 60.980 ;
        RECT 72.640 59.540 74.070 59.570 ;
        RECT 72.230 58.830 74.070 59.540 ;
        RECT 54.670 58.670 55.060 58.680 ;
        RECT 54.670 56.510 55.690 58.670 ;
        RECT 54.670 52.690 55.060 56.510 ;
        RECT 56.150 56.270 57.150 58.670 ;
        RECT 57.640 56.540 58.640 58.690 ;
        RECT 55.900 56.040 57.150 56.270 ;
        RECT 55.340 55.880 57.150 56.040 ;
        RECT 57.410 55.900 58.640 56.540 ;
        RECT 59.120 56.530 60.120 58.680 ;
        RECT 60.580 56.530 61.580 58.670 ;
        RECT 55.340 55.580 56.620 55.880 ;
        RECT 55.340 53.700 56.340 55.580 ;
        RECT 57.410 55.430 58.090 55.900 ;
        RECT 58.900 55.890 60.120 56.530 ;
        RECT 58.900 55.430 59.580 55.890 ;
        RECT 60.390 55.880 61.580 56.530 ;
        RECT 62.080 56.500 63.080 58.690 ;
        RECT 65.020 58.670 67.330 58.680 ;
        RECT 61.840 55.900 63.080 56.500 ;
        RECT 63.590 56.490 64.590 58.670 ;
        RECT 65.020 56.500 67.500 58.670 ;
        RECT 60.390 55.430 61.070 55.880 ;
        RECT 61.840 55.430 62.520 55.900 ;
        RECT 56.790 54.960 58.090 55.430 ;
        RECT 56.790 53.790 57.830 54.960 ;
        RECT 58.300 54.950 59.580 55.430 ;
        RECT 59.770 54.950 61.070 55.430 ;
        RECT 58.300 53.790 59.340 54.950 ;
        RECT 59.770 53.790 60.810 54.950 ;
        RECT 61.260 54.920 62.520 55.430 ;
        RECT 63.340 55.880 64.590 56.490 ;
        RECT 64.850 55.890 67.500 56.500 ;
        RECT 63.340 55.420 64.020 55.880 ;
        RECT 64.850 55.430 65.530 55.890 ;
        RECT 66.500 55.880 67.500 55.890 ;
        RECT 72.230 55.590 72.890 58.830 ;
        RECT 74.560 58.770 75.260 64.260 ;
        RECT 75.510 63.780 76.720 64.440 ;
        RECT 77.870 64.550 78.190 66.765 ;
        RECT 78.870 66.560 79.770 67.370 ;
        RECT 80.340 66.830 80.860 74.720 ;
        RECT 80.340 66.765 80.570 66.830 ;
        RECT 81.340 66.820 81.720 74.740 ;
        RECT 82.340 74.300 83.310 74.970 ;
        RECT 83.770 74.720 84.000 74.765 ;
        RECT 84.910 74.720 85.140 74.765 ;
        RECT 82.420 68.340 83.240 74.300 ;
        RECT 82.330 67.340 83.330 68.340 ;
        RECT 81.350 66.765 81.710 66.820 ;
        RECT 78.330 66.330 80.290 66.560 ;
        RECT 81.350 65.200 81.610 66.765 ;
        RECT 82.420 66.560 83.240 67.340 ;
        RECT 83.770 66.850 85.150 74.720 ;
        RECT 85.480 74.600 85.920 74.970 ;
        RECT 86.200 74.720 86.430 74.765 ;
        RECT 86.830 74.720 88.580 75.530 ;
        RECT 90.070 75.560 147.960 75.570 ;
        RECT 90.070 75.510 102.950 75.560 ;
        RECT 105.080 75.540 147.960 75.560 ;
        RECT 105.080 75.510 132.970 75.540 ;
        RECT 135.080 75.510 147.960 75.540 ;
        RECT 90.880 75.150 91.840 75.180 ;
        RECT 85.480 67.230 85.910 74.600 ;
        RECT 86.200 74.410 88.580 74.720 ;
        RECT 90.550 74.950 91.840 75.150 ;
        RECT 90.550 74.710 91.610 74.950 ;
        RECT 92.110 74.745 92.330 75.510 ;
        RECT 97.310 75.180 98.280 75.240 ;
        RECT 93.310 74.950 95.270 75.180 ;
        RECT 96.740 74.950 98.700 75.180 ;
        RECT 100.170 74.950 101.130 75.180 ;
        RECT 86.200 70.740 87.970 74.410 ;
        RECT 86.200 69.740 87.960 70.740 ;
        RECT 83.770 66.765 84.000 66.850 ;
        RECT 84.910 66.765 85.140 66.850 ;
        RECT 85.480 66.560 85.920 67.230 ;
        RECT 86.200 66.860 87.970 69.740 ;
        RECT 90.500 67.600 91.610 74.710 ;
        RECT 86.200 66.765 86.430 66.860 ;
        RECT 81.760 66.330 83.720 66.560 ;
        RECT 85.190 66.330 86.150 66.560 ;
        RECT 85.290 65.450 86.080 66.330 ;
        RECT 86.830 65.850 87.970 66.860 ;
        RECT 81.350 64.580 84.970 65.200 ;
        RECT 85.240 64.690 86.130 65.450 ;
        RECT 75.510 63.550 76.870 63.780 ;
        RECT 75.510 62.380 76.600 63.550 ;
        RECT 77.870 63.390 78.200 64.550 ;
        RECT 78.340 63.550 80.300 63.780 ;
        RECT 75.520 59.430 76.600 62.380 ;
        RECT 75.570 59.230 76.600 59.430 ;
        RECT 76.920 63.380 77.150 63.390 ;
        RECT 76.920 61.070 77.330 63.380 ;
        RECT 77.870 63.370 78.290 63.390 ;
        RECT 77.870 63.320 78.380 63.370 ;
        RECT 78.730 63.320 79.990 63.550 ;
        RECT 81.350 63.390 81.610 64.580 ;
        RECT 84.560 63.930 84.960 64.580 ;
        RECT 86.900 64.530 87.970 65.850 ;
        RECT 90.490 66.540 91.610 67.600 ;
        RECT 91.890 74.540 92.330 74.745 ;
        RECT 93.030 74.720 93.260 74.745 ;
        RECT 93.030 74.710 93.270 74.720 ;
        RECT 91.890 66.800 92.280 74.540 ;
        RECT 92.860 67.650 93.270 74.710 ;
        RECT 93.850 70.220 94.750 74.950 ;
        RECT 95.320 74.700 95.550 74.745 ;
        RECT 96.460 74.720 96.690 74.745 ;
        RECT 93.840 69.110 94.790 70.220 ;
        RECT 93.850 68.360 94.750 69.110 ;
        RECT 92.850 66.830 93.270 67.650 ;
        RECT 93.820 67.350 94.820 68.360 ;
        RECT 91.890 66.745 92.120 66.800 ;
        RECT 92.850 66.745 93.260 66.830 ;
        RECT 90.490 66.310 91.840 66.540 ;
        RECT 90.490 65.670 91.700 66.310 ;
        RECT 86.900 64.030 88.740 64.530 ;
        RECT 90.050 64.420 91.700 65.670 ;
        RECT 85.960 63.930 86.710 63.940 ;
        RECT 84.560 63.880 86.710 63.930 ;
        RECT 84.560 63.840 86.890 63.880 ;
        RECT 81.770 63.550 83.730 63.780 ;
        RECT 84.560 63.590 88.120 63.840 ;
        RECT 84.560 63.580 85.900 63.590 ;
        RECT 85.610 63.560 85.900 63.580 ;
        RECT 76.920 59.390 77.420 61.070 ;
        RECT 77.870 59.460 79.990 63.320 ;
        RECT 77.990 59.450 79.990 59.460 ;
        RECT 78.060 59.390 78.290 59.450 ;
        RECT 75.570 59.050 76.870 59.230 ;
        RECT 75.910 59.000 76.870 59.050 ;
        RECT 77.220 58.770 77.420 59.390 ;
        RECT 78.650 59.230 79.990 59.450 ;
        RECT 80.350 63.350 80.580 63.390 ;
        RECT 81.350 63.360 81.720 63.390 ;
        RECT 81.350 63.350 81.800 63.360 ;
        RECT 80.350 63.340 80.760 63.350 ;
        RECT 80.350 61.120 80.800 63.340 ;
        RECT 80.350 60.630 80.850 61.120 ;
        RECT 80.350 59.960 80.940 60.630 ;
        RECT 80.350 59.710 81.000 59.960 ;
        RECT 80.350 59.680 81.050 59.710 ;
        RECT 80.350 59.390 80.580 59.680 ;
        RECT 80.810 59.310 81.050 59.680 ;
        RECT 81.300 59.450 81.800 63.350 ;
        RECT 81.300 59.440 81.720 59.450 ;
        RECT 81.360 59.430 81.720 59.440 ;
        RECT 81.490 59.390 81.720 59.430 ;
        RECT 78.340 59.000 80.300 59.230 ;
        RECT 80.730 59.070 81.050 59.310 ;
        RECT 82.060 59.230 83.430 63.550 ;
        RECT 86.770 63.500 88.120 63.590 ;
        RECT 87.720 63.495 88.010 63.500 ;
        RECT 83.780 63.210 84.010 63.390 ;
        RECT 85.420 63.340 85.650 63.400 ;
        RECT 85.860 63.340 86.090 63.400 ;
        RECT 84.670 63.330 85.650 63.340 ;
        RECT 84.240 63.210 85.650 63.330 ;
        RECT 83.780 62.460 85.650 63.210 ;
        RECT 85.840 63.200 86.240 63.340 ;
        RECT 88.370 63.290 88.740 64.030 ;
        RECT 87.530 63.200 87.760 63.290 ;
        RECT 85.840 62.470 87.800 63.200 ;
        RECT 85.840 62.460 86.240 62.470 ;
        RECT 83.780 62.000 85.140 62.460 ;
        RECT 85.420 62.400 85.650 62.460 ;
        RECT 85.860 62.400 86.090 62.460 ;
        RECT 83.780 61.730 86.240 62.000 ;
        RECT 83.780 61.690 85.950 61.730 ;
        RECT 83.780 59.940 85.130 61.690 ;
        RECT 86.410 61.510 87.790 62.470 ;
        RECT 86.410 61.380 87.810 61.510 ;
        RECT 85.690 60.380 87.810 61.380 ;
        RECT 86.410 60.350 87.810 60.380 ;
        RECT 87.530 60.340 87.810 60.350 ;
        RECT 87.970 60.350 88.740 63.290 ;
        RECT 90.490 63.760 91.700 64.420 ;
        RECT 92.850 64.530 93.170 66.745 ;
        RECT 93.850 66.540 94.750 67.350 ;
        RECT 95.320 66.810 95.840 74.700 ;
        RECT 95.320 66.745 95.550 66.810 ;
        RECT 96.320 66.800 96.700 74.720 ;
        RECT 97.310 74.310 98.280 74.950 ;
        RECT 98.750 74.700 98.980 74.745 ;
        RECT 99.890 74.700 100.120 74.745 ;
        RECT 97.400 68.320 98.220 74.310 ;
        RECT 97.310 67.320 98.310 68.320 ;
        RECT 96.330 66.745 96.690 66.800 ;
        RECT 93.310 66.310 95.270 66.540 ;
        RECT 96.330 65.180 96.590 66.745 ;
        RECT 97.400 66.540 98.220 67.320 ;
        RECT 98.750 66.830 100.130 74.700 ;
        RECT 100.460 74.580 100.900 74.950 ;
        RECT 101.180 74.700 101.410 74.745 ;
        RECT 101.810 74.700 102.950 75.510 ;
        RECT 105.890 75.150 106.850 75.180 ;
        RECT 105.560 74.950 106.850 75.150 ;
        RECT 105.560 74.710 106.620 74.950 ;
        RECT 107.120 74.745 107.340 75.510 ;
        RECT 116.820 75.500 120.800 75.510 ;
        RECT 112.240 75.180 113.270 75.260 ;
        RECT 108.320 74.950 110.280 75.180 ;
        RECT 111.750 74.950 113.710 75.180 ;
        RECT 115.180 74.950 116.140 75.180 ;
        RECT 100.460 67.210 100.890 74.580 ;
        RECT 101.180 70.720 102.950 74.700 ;
        RECT 101.180 69.720 102.940 70.720 ;
        RECT 98.750 66.745 98.980 66.830 ;
        RECT 99.890 66.745 100.120 66.830 ;
        RECT 100.460 66.540 100.900 67.210 ;
        RECT 101.180 66.840 102.950 69.720 ;
        RECT 105.510 67.600 106.620 74.710 ;
        RECT 101.180 66.745 101.410 66.840 ;
        RECT 96.740 66.310 98.700 66.540 ;
        RECT 100.170 66.310 101.130 66.540 ;
        RECT 100.270 65.430 101.060 66.310 ;
        RECT 101.810 65.830 102.950 66.840 ;
        RECT 96.330 64.560 99.950 65.180 ;
        RECT 100.220 64.670 101.110 65.430 ;
        RECT 90.490 63.530 91.850 63.760 ;
        RECT 90.490 62.360 91.580 63.530 ;
        RECT 92.850 63.370 93.180 64.530 ;
        RECT 93.320 63.530 95.280 63.760 ;
        RECT 87.530 60.290 87.760 60.340 ;
        RECT 87.970 60.290 88.200 60.350 ;
        RECT 83.780 59.620 86.480 59.940 ;
        RECT 83.780 59.390 84.010 59.620 ;
        RECT 80.690 58.770 81.050 59.070 ;
        RECT 81.770 59.000 83.730 59.230 ;
        RECT 84.390 58.770 86.480 59.620 ;
        RECT 90.500 59.410 91.580 62.360 ;
        RECT 90.550 59.210 91.580 59.410 ;
        RECT 91.900 63.360 92.130 63.370 ;
        RECT 91.900 61.050 92.310 63.360 ;
        RECT 92.850 63.350 93.270 63.370 ;
        RECT 92.850 63.300 93.360 63.350 ;
        RECT 93.710 63.300 94.970 63.530 ;
        RECT 96.330 63.370 96.590 64.560 ;
        RECT 99.540 63.910 99.940 64.560 ;
        RECT 101.880 64.510 102.950 65.830 ;
        RECT 105.500 66.540 106.620 67.600 ;
        RECT 106.900 74.540 107.340 74.745 ;
        RECT 108.040 74.720 108.270 74.745 ;
        RECT 108.040 74.710 108.280 74.720 ;
        RECT 106.900 66.800 107.290 74.540 ;
        RECT 107.870 67.650 108.280 74.710 ;
        RECT 108.860 69.950 109.760 74.950 ;
        RECT 110.330 74.700 110.560 74.745 ;
        RECT 111.470 74.720 111.700 74.745 ;
        RECT 108.860 68.840 109.820 69.950 ;
        RECT 108.860 68.360 109.760 68.840 ;
        RECT 107.860 66.830 108.280 67.650 ;
        RECT 108.830 67.350 109.830 68.360 ;
        RECT 106.900 66.745 107.130 66.800 ;
        RECT 107.860 66.745 108.270 66.830 ;
        RECT 105.500 66.310 106.850 66.540 ;
        RECT 105.500 65.670 106.710 66.310 ;
        RECT 101.880 64.010 103.720 64.510 ;
        RECT 105.060 64.420 106.710 65.670 ;
        RECT 100.940 63.910 101.690 63.920 ;
        RECT 99.540 63.860 101.690 63.910 ;
        RECT 99.540 63.820 101.870 63.860 ;
        RECT 96.750 63.530 98.710 63.760 ;
        RECT 99.540 63.570 103.100 63.820 ;
        RECT 99.540 63.560 100.880 63.570 ;
        RECT 100.590 63.540 100.880 63.560 ;
        RECT 91.900 59.370 92.400 61.050 ;
        RECT 92.850 59.440 94.970 63.300 ;
        RECT 92.970 59.430 94.970 59.440 ;
        RECT 93.040 59.370 93.270 59.430 ;
        RECT 90.550 59.030 91.850 59.210 ;
        RECT 90.890 58.980 91.850 59.030 ;
        RECT 74.560 58.730 86.480 58.770 ;
        RECT 87.050 58.730 88.200 58.790 ;
        RECT 92.200 58.750 92.400 59.370 ;
        RECT 93.630 59.210 94.970 59.430 ;
        RECT 95.330 63.330 95.560 63.370 ;
        RECT 96.330 63.340 96.700 63.370 ;
        RECT 96.330 63.330 96.780 63.340 ;
        RECT 95.330 63.320 95.740 63.330 ;
        RECT 95.330 61.100 95.780 63.320 ;
        RECT 95.330 60.610 95.830 61.100 ;
        RECT 95.330 59.940 95.920 60.610 ;
        RECT 95.330 59.690 95.980 59.940 ;
        RECT 95.330 59.660 96.030 59.690 ;
        RECT 95.330 59.370 95.560 59.660 ;
        RECT 95.790 59.290 96.030 59.660 ;
        RECT 96.280 59.430 96.780 63.330 ;
        RECT 96.280 59.420 96.700 59.430 ;
        RECT 96.340 59.410 96.700 59.420 ;
        RECT 96.470 59.370 96.700 59.410 ;
        RECT 93.320 58.980 95.280 59.210 ;
        RECT 95.710 59.050 96.030 59.290 ;
        RECT 97.040 59.210 98.410 63.530 ;
        RECT 101.750 63.480 103.100 63.570 ;
        RECT 102.700 63.475 102.990 63.480 ;
        RECT 98.760 63.190 98.990 63.370 ;
        RECT 100.400 63.320 100.630 63.380 ;
        RECT 100.840 63.320 101.070 63.380 ;
        RECT 99.650 63.310 100.630 63.320 ;
        RECT 99.220 63.190 100.630 63.310 ;
        RECT 98.760 62.440 100.630 63.190 ;
        RECT 100.820 63.180 101.220 63.320 ;
        RECT 103.350 63.270 103.720 64.010 ;
        RECT 102.510 63.180 102.740 63.270 ;
        RECT 100.820 62.450 102.780 63.180 ;
        RECT 100.820 62.440 101.220 62.450 ;
        RECT 98.760 61.980 100.120 62.440 ;
        RECT 100.400 62.380 100.630 62.440 ;
        RECT 100.840 62.380 101.070 62.440 ;
        RECT 98.760 61.710 101.220 61.980 ;
        RECT 98.760 61.670 100.930 61.710 ;
        RECT 98.760 59.920 100.110 61.670 ;
        RECT 101.390 61.490 102.770 62.450 ;
        RECT 101.390 61.360 102.790 61.490 ;
        RECT 100.670 60.360 102.790 61.360 ;
        RECT 101.390 60.330 102.790 60.360 ;
        RECT 102.510 60.320 102.790 60.330 ;
        RECT 102.950 60.330 103.720 63.270 ;
        RECT 105.500 63.760 106.710 64.420 ;
        RECT 107.860 64.530 108.180 66.745 ;
        RECT 108.860 66.540 109.760 67.350 ;
        RECT 110.330 66.810 110.850 74.700 ;
        RECT 110.330 66.745 110.560 66.810 ;
        RECT 111.330 66.800 111.710 74.720 ;
        RECT 112.240 74.270 113.270 74.950 ;
        RECT 113.760 74.700 113.990 74.745 ;
        RECT 114.900 74.700 115.130 74.745 ;
        RECT 112.410 68.320 113.230 74.270 ;
        RECT 112.320 67.320 113.320 68.320 ;
        RECT 111.340 66.745 111.700 66.800 ;
        RECT 108.320 66.310 110.280 66.540 ;
        RECT 111.340 65.180 111.600 66.745 ;
        RECT 112.410 66.540 113.230 67.320 ;
        RECT 113.760 66.830 115.140 74.700 ;
        RECT 115.470 74.580 115.910 74.950 ;
        RECT 116.190 74.700 116.420 74.745 ;
        RECT 116.820 74.700 117.960 75.500 ;
        RECT 120.900 75.150 121.860 75.180 ;
        RECT 120.570 74.950 121.860 75.150 ;
        RECT 120.570 74.710 121.630 74.950 ;
        RECT 122.130 74.745 122.350 75.510 ;
        RECT 127.350 75.180 128.320 75.230 ;
        RECT 123.330 74.950 125.290 75.180 ;
        RECT 126.760 74.950 128.720 75.180 ;
        RECT 130.190 74.950 131.150 75.180 ;
        RECT 115.470 67.210 115.900 74.580 ;
        RECT 116.190 70.720 117.960 74.700 ;
        RECT 116.190 69.720 117.950 70.720 ;
        RECT 113.760 66.745 113.990 66.830 ;
        RECT 114.900 66.745 115.130 66.830 ;
        RECT 115.470 66.540 115.910 67.210 ;
        RECT 116.190 66.840 117.960 69.720 ;
        RECT 120.520 67.600 121.630 74.710 ;
        RECT 116.190 66.745 116.420 66.840 ;
        RECT 111.750 66.310 113.710 66.540 ;
        RECT 115.180 66.310 116.140 66.540 ;
        RECT 115.280 65.430 116.070 66.310 ;
        RECT 116.820 65.830 117.960 66.840 ;
        RECT 111.340 64.560 114.960 65.180 ;
        RECT 115.230 64.670 116.120 65.430 ;
        RECT 105.500 63.530 106.860 63.760 ;
        RECT 105.500 62.360 106.590 63.530 ;
        RECT 107.860 63.370 108.190 64.530 ;
        RECT 108.330 63.530 110.290 63.760 ;
        RECT 102.510 60.270 102.740 60.320 ;
        RECT 102.950 60.270 103.180 60.330 ;
        RECT 98.760 59.600 101.460 59.920 ;
        RECT 98.760 59.370 98.990 59.600 ;
        RECT 95.670 58.750 96.030 59.050 ;
        RECT 96.750 58.980 98.710 59.210 ;
        RECT 99.370 58.750 101.460 59.600 ;
        RECT 105.510 59.410 106.590 62.360 ;
        RECT 105.560 59.210 106.590 59.410 ;
        RECT 106.910 63.360 107.140 63.370 ;
        RECT 106.910 61.050 107.320 63.360 ;
        RECT 107.860 63.350 108.280 63.370 ;
        RECT 107.860 63.300 108.370 63.350 ;
        RECT 108.720 63.300 109.980 63.530 ;
        RECT 111.340 63.370 111.600 64.560 ;
        RECT 114.550 63.910 114.950 64.560 ;
        RECT 116.890 64.510 117.960 65.830 ;
        RECT 120.510 66.540 121.630 67.600 ;
        RECT 121.910 74.540 122.350 74.745 ;
        RECT 123.050 74.720 123.280 74.745 ;
        RECT 123.050 74.710 123.290 74.720 ;
        RECT 121.910 66.800 122.300 74.540 ;
        RECT 122.880 67.650 123.290 74.710 ;
        RECT 123.870 70.310 124.770 74.950 ;
        RECT 125.340 74.700 125.570 74.745 ;
        RECT 126.480 74.720 126.710 74.745 ;
        RECT 123.720 69.010 124.920 70.310 ;
        RECT 123.870 68.360 124.770 69.010 ;
        RECT 122.870 66.830 123.290 67.650 ;
        RECT 123.840 67.350 124.840 68.360 ;
        RECT 121.910 66.745 122.140 66.800 ;
        RECT 122.870 66.745 123.280 66.830 ;
        RECT 120.510 66.310 121.860 66.540 ;
        RECT 120.510 65.670 121.720 66.310 ;
        RECT 116.890 64.010 118.730 64.510 ;
        RECT 120.070 64.420 121.720 65.670 ;
        RECT 115.950 63.910 116.700 63.920 ;
        RECT 114.550 63.860 116.700 63.910 ;
        RECT 114.550 63.820 116.880 63.860 ;
        RECT 111.760 63.530 113.720 63.760 ;
        RECT 114.550 63.570 118.110 63.820 ;
        RECT 114.550 63.560 115.890 63.570 ;
        RECT 115.600 63.540 115.890 63.560 ;
        RECT 106.910 59.370 107.410 61.050 ;
        RECT 107.860 59.440 109.980 63.300 ;
        RECT 107.980 59.430 109.980 59.440 ;
        RECT 108.050 59.370 108.280 59.430 ;
        RECT 105.560 59.030 106.860 59.210 ;
        RECT 105.900 58.980 106.860 59.030 ;
        RECT 107.210 58.750 107.410 59.370 ;
        RECT 108.640 59.210 109.980 59.430 ;
        RECT 110.340 63.330 110.570 63.370 ;
        RECT 111.340 63.340 111.710 63.370 ;
        RECT 111.340 63.330 111.790 63.340 ;
        RECT 110.340 63.320 110.750 63.330 ;
        RECT 110.340 61.100 110.790 63.320 ;
        RECT 110.340 60.610 110.840 61.100 ;
        RECT 110.340 59.940 110.930 60.610 ;
        RECT 110.340 59.690 110.990 59.940 ;
        RECT 110.340 59.660 111.040 59.690 ;
        RECT 110.340 59.370 110.570 59.660 ;
        RECT 110.800 59.290 111.040 59.660 ;
        RECT 111.290 59.430 111.790 63.330 ;
        RECT 111.290 59.420 111.710 59.430 ;
        RECT 111.350 59.410 111.710 59.420 ;
        RECT 111.480 59.370 111.710 59.410 ;
        RECT 108.330 58.980 110.290 59.210 ;
        RECT 110.720 59.050 111.040 59.290 ;
        RECT 112.050 59.210 113.420 63.530 ;
        RECT 116.760 63.480 118.110 63.570 ;
        RECT 117.710 63.475 118.000 63.480 ;
        RECT 113.770 63.190 114.000 63.370 ;
        RECT 115.410 63.320 115.640 63.380 ;
        RECT 115.850 63.320 116.080 63.380 ;
        RECT 114.660 63.310 115.640 63.320 ;
        RECT 114.230 63.190 115.640 63.310 ;
        RECT 113.770 62.440 115.640 63.190 ;
        RECT 115.830 63.180 116.230 63.320 ;
        RECT 118.360 63.270 118.730 64.010 ;
        RECT 117.520 63.180 117.750 63.270 ;
        RECT 115.830 62.450 117.790 63.180 ;
        RECT 115.830 62.440 116.230 62.450 ;
        RECT 113.770 61.980 115.130 62.440 ;
        RECT 115.410 62.380 115.640 62.440 ;
        RECT 115.850 62.380 116.080 62.440 ;
        RECT 113.770 61.710 116.230 61.980 ;
        RECT 113.770 61.670 115.940 61.710 ;
        RECT 113.770 59.920 115.120 61.670 ;
        RECT 116.400 61.490 117.780 62.450 ;
        RECT 116.400 61.360 117.800 61.490 ;
        RECT 115.680 60.360 117.800 61.360 ;
        RECT 116.400 60.330 117.800 60.360 ;
        RECT 117.520 60.320 117.800 60.330 ;
        RECT 117.960 60.330 118.730 63.270 ;
        RECT 120.510 63.760 121.720 64.420 ;
        RECT 122.870 64.530 123.190 66.745 ;
        RECT 123.870 66.540 124.770 67.350 ;
        RECT 125.340 66.810 125.860 74.700 ;
        RECT 125.340 66.745 125.570 66.810 ;
        RECT 126.340 66.800 126.720 74.720 ;
        RECT 127.350 74.380 128.320 74.950 ;
        RECT 128.770 74.700 129.000 74.745 ;
        RECT 129.910 74.700 130.140 74.745 ;
        RECT 127.420 68.320 128.240 74.380 ;
        RECT 127.330 67.320 128.330 68.320 ;
        RECT 126.350 66.745 126.710 66.800 ;
        RECT 123.330 66.310 125.290 66.540 ;
        RECT 126.350 65.180 126.610 66.745 ;
        RECT 127.420 66.540 128.240 67.320 ;
        RECT 128.770 66.830 130.150 74.700 ;
        RECT 130.480 74.580 130.920 74.950 ;
        RECT 131.200 74.700 131.430 74.745 ;
        RECT 131.830 74.700 132.970 75.510 ;
        RECT 135.890 75.150 136.850 75.180 ;
        RECT 135.560 74.950 136.850 75.150 ;
        RECT 135.560 74.710 136.620 74.950 ;
        RECT 137.120 74.745 137.340 75.510 ;
        RECT 142.330 75.180 143.300 75.230 ;
        RECT 138.320 74.950 140.280 75.180 ;
        RECT 141.750 74.950 143.710 75.180 ;
        RECT 145.180 74.950 146.140 75.180 ;
        RECT 130.480 67.210 130.910 74.580 ;
        RECT 131.200 70.720 132.970 74.700 ;
        RECT 131.200 69.720 132.960 70.720 ;
        RECT 128.770 66.745 129.000 66.830 ;
        RECT 129.910 66.745 130.140 66.830 ;
        RECT 130.480 66.540 130.920 67.210 ;
        RECT 131.200 66.840 132.970 69.720 ;
        RECT 135.510 67.600 136.620 74.710 ;
        RECT 131.200 66.745 131.430 66.840 ;
        RECT 126.760 66.310 128.720 66.540 ;
        RECT 130.190 66.310 131.150 66.540 ;
        RECT 130.290 65.430 131.080 66.310 ;
        RECT 131.830 65.830 132.970 66.840 ;
        RECT 126.350 64.560 129.970 65.180 ;
        RECT 130.240 64.670 131.130 65.430 ;
        RECT 120.510 63.530 121.870 63.760 ;
        RECT 120.510 62.360 121.600 63.530 ;
        RECT 122.870 63.370 123.200 64.530 ;
        RECT 123.340 63.530 125.300 63.760 ;
        RECT 117.520 60.270 117.750 60.320 ;
        RECT 117.960 60.270 118.190 60.330 ;
        RECT 113.770 59.600 116.470 59.920 ;
        RECT 113.770 59.370 114.000 59.600 ;
        RECT 110.680 58.750 111.040 59.050 ;
        RECT 111.760 58.980 113.720 59.210 ;
        RECT 114.380 58.750 116.470 59.600 ;
        RECT 120.520 59.410 121.600 62.360 ;
        RECT 120.570 59.210 121.600 59.410 ;
        RECT 121.920 63.360 122.150 63.370 ;
        RECT 121.920 61.050 122.330 63.360 ;
        RECT 122.870 63.350 123.290 63.370 ;
        RECT 122.870 63.300 123.380 63.350 ;
        RECT 123.730 63.300 124.990 63.530 ;
        RECT 126.350 63.370 126.610 64.560 ;
        RECT 129.560 63.910 129.960 64.560 ;
        RECT 131.900 64.510 132.970 65.830 ;
        RECT 135.500 66.540 136.620 67.600 ;
        RECT 136.900 74.540 137.340 74.745 ;
        RECT 138.040 74.720 138.270 74.745 ;
        RECT 138.040 74.710 138.280 74.720 ;
        RECT 136.900 66.800 137.290 74.540 ;
        RECT 137.870 67.650 138.280 74.710 ;
        RECT 138.860 70.290 139.760 74.950 ;
        RECT 140.330 74.700 140.560 74.745 ;
        RECT 141.470 74.720 141.700 74.745 ;
        RECT 138.850 69.210 139.790 70.290 ;
        RECT 138.860 68.360 139.760 69.210 ;
        RECT 137.860 66.830 138.280 67.650 ;
        RECT 138.830 67.350 139.830 68.360 ;
        RECT 136.900 66.745 137.130 66.800 ;
        RECT 137.860 66.745 138.270 66.830 ;
        RECT 135.500 66.310 136.850 66.540 ;
        RECT 135.500 65.670 136.710 66.310 ;
        RECT 131.900 64.010 133.740 64.510 ;
        RECT 135.060 64.420 136.710 65.670 ;
        RECT 130.960 63.910 131.710 63.920 ;
        RECT 129.560 63.860 131.710 63.910 ;
        RECT 129.560 63.820 131.890 63.860 ;
        RECT 126.770 63.530 128.730 63.760 ;
        RECT 129.560 63.570 133.120 63.820 ;
        RECT 129.560 63.560 130.900 63.570 ;
        RECT 130.610 63.540 130.900 63.560 ;
        RECT 121.920 59.370 122.420 61.050 ;
        RECT 122.870 59.440 124.990 63.300 ;
        RECT 122.990 59.430 124.990 59.440 ;
        RECT 123.060 59.370 123.290 59.430 ;
        RECT 120.570 59.030 121.870 59.210 ;
        RECT 120.910 58.980 121.870 59.030 ;
        RECT 122.220 58.750 122.420 59.370 ;
        RECT 123.650 59.210 124.990 59.430 ;
        RECT 125.350 63.330 125.580 63.370 ;
        RECT 126.350 63.340 126.720 63.370 ;
        RECT 126.350 63.330 126.800 63.340 ;
        RECT 125.350 63.320 125.760 63.330 ;
        RECT 125.350 61.100 125.800 63.320 ;
        RECT 125.350 60.610 125.850 61.100 ;
        RECT 125.350 59.940 125.940 60.610 ;
        RECT 125.350 59.690 126.000 59.940 ;
        RECT 125.350 59.660 126.050 59.690 ;
        RECT 125.350 59.370 125.580 59.660 ;
        RECT 125.810 59.290 126.050 59.660 ;
        RECT 126.300 59.430 126.800 63.330 ;
        RECT 126.300 59.420 126.720 59.430 ;
        RECT 126.360 59.410 126.720 59.420 ;
        RECT 126.490 59.370 126.720 59.410 ;
        RECT 123.340 58.980 125.300 59.210 ;
        RECT 125.730 59.050 126.050 59.290 ;
        RECT 127.060 59.210 128.430 63.530 ;
        RECT 131.770 63.480 133.120 63.570 ;
        RECT 132.720 63.475 133.010 63.480 ;
        RECT 128.780 63.190 129.010 63.370 ;
        RECT 130.420 63.320 130.650 63.380 ;
        RECT 130.860 63.320 131.090 63.380 ;
        RECT 129.670 63.310 130.650 63.320 ;
        RECT 129.240 63.190 130.650 63.310 ;
        RECT 128.780 62.440 130.650 63.190 ;
        RECT 130.840 63.180 131.240 63.320 ;
        RECT 133.370 63.270 133.740 64.010 ;
        RECT 132.530 63.180 132.760 63.270 ;
        RECT 130.840 62.450 132.800 63.180 ;
        RECT 130.840 62.440 131.240 62.450 ;
        RECT 128.780 61.980 130.140 62.440 ;
        RECT 130.420 62.380 130.650 62.440 ;
        RECT 130.860 62.380 131.090 62.440 ;
        RECT 128.780 61.710 131.240 61.980 ;
        RECT 128.780 61.670 130.950 61.710 ;
        RECT 128.780 59.920 130.130 61.670 ;
        RECT 131.410 61.490 132.790 62.450 ;
        RECT 131.410 61.360 132.810 61.490 ;
        RECT 130.690 60.360 132.810 61.360 ;
        RECT 131.410 60.330 132.810 60.360 ;
        RECT 132.530 60.320 132.810 60.330 ;
        RECT 132.970 60.330 133.740 63.270 ;
        RECT 135.500 63.760 136.710 64.420 ;
        RECT 137.860 64.530 138.180 66.745 ;
        RECT 138.860 66.540 139.760 67.350 ;
        RECT 140.330 66.810 140.850 74.700 ;
        RECT 140.330 66.745 140.560 66.810 ;
        RECT 141.330 66.800 141.710 74.720 ;
        RECT 142.330 74.380 143.300 74.950 ;
        RECT 143.760 74.700 143.990 74.745 ;
        RECT 144.900 74.700 145.130 74.745 ;
        RECT 142.410 68.320 143.230 74.380 ;
        RECT 142.320 67.320 143.320 68.320 ;
        RECT 141.340 66.745 141.700 66.800 ;
        RECT 138.320 66.310 140.280 66.540 ;
        RECT 141.340 65.180 141.600 66.745 ;
        RECT 142.410 66.540 143.230 67.320 ;
        RECT 143.760 66.830 145.140 74.700 ;
        RECT 145.470 74.580 145.910 74.950 ;
        RECT 146.190 74.700 146.420 74.745 ;
        RECT 146.820 74.700 147.960 75.510 ;
        RECT 145.470 67.210 145.900 74.580 ;
        RECT 146.190 70.720 147.960 74.700 ;
        RECT 146.190 69.720 147.950 70.720 ;
        RECT 143.760 66.745 143.990 66.830 ;
        RECT 144.900 66.745 145.130 66.830 ;
        RECT 145.470 66.540 145.910 67.210 ;
        RECT 146.190 66.840 147.960 69.720 ;
        RECT 146.190 66.745 146.420 66.840 ;
        RECT 141.750 66.310 143.710 66.540 ;
        RECT 145.180 66.310 146.140 66.540 ;
        RECT 145.280 65.430 146.070 66.310 ;
        RECT 146.820 65.830 147.960 66.840 ;
        RECT 141.340 64.560 144.960 65.180 ;
        RECT 145.230 64.670 146.120 65.430 ;
        RECT 135.500 63.530 136.860 63.760 ;
        RECT 135.500 62.360 136.590 63.530 ;
        RECT 137.860 63.370 138.190 64.530 ;
        RECT 138.330 63.530 140.290 63.760 ;
        RECT 132.530 60.270 132.760 60.320 ;
        RECT 132.970 60.270 133.200 60.330 ;
        RECT 128.780 59.600 131.480 59.920 ;
        RECT 128.780 59.370 129.010 59.600 ;
        RECT 125.690 58.750 126.050 59.050 ;
        RECT 126.770 58.980 128.730 59.210 ;
        RECT 129.390 58.750 131.480 59.600 ;
        RECT 135.510 59.410 136.590 62.360 ;
        RECT 135.560 59.210 136.590 59.410 ;
        RECT 136.910 63.360 137.140 63.370 ;
        RECT 136.910 61.050 137.320 63.360 ;
        RECT 137.860 63.350 138.280 63.370 ;
        RECT 137.860 63.300 138.370 63.350 ;
        RECT 138.720 63.300 139.980 63.530 ;
        RECT 141.340 63.370 141.600 64.560 ;
        RECT 144.550 63.910 144.950 64.560 ;
        RECT 146.890 64.510 147.960 65.830 ;
        RECT 146.890 64.010 148.730 64.510 ;
        RECT 145.950 63.910 146.700 63.920 ;
        RECT 144.550 63.860 146.700 63.910 ;
        RECT 144.550 63.820 146.880 63.860 ;
        RECT 141.760 63.530 143.720 63.760 ;
        RECT 144.550 63.570 148.110 63.820 ;
        RECT 144.550 63.560 145.890 63.570 ;
        RECT 145.600 63.540 145.890 63.560 ;
        RECT 136.910 59.370 137.410 61.050 ;
        RECT 137.860 59.440 139.980 63.300 ;
        RECT 137.980 59.430 139.980 59.440 ;
        RECT 138.050 59.370 138.280 59.430 ;
        RECT 135.560 59.030 136.860 59.210 ;
        RECT 135.900 58.980 136.860 59.030 ;
        RECT 137.210 58.750 137.410 59.370 ;
        RECT 138.640 59.210 139.980 59.430 ;
        RECT 140.340 63.330 140.570 63.370 ;
        RECT 141.340 63.340 141.710 63.370 ;
        RECT 141.340 63.330 141.790 63.340 ;
        RECT 140.340 63.320 140.750 63.330 ;
        RECT 140.340 61.100 140.790 63.320 ;
        RECT 140.340 60.610 140.840 61.100 ;
        RECT 140.340 59.940 140.930 60.610 ;
        RECT 140.340 59.690 140.990 59.940 ;
        RECT 140.340 59.660 141.040 59.690 ;
        RECT 140.340 59.370 140.570 59.660 ;
        RECT 140.800 59.290 141.040 59.660 ;
        RECT 141.290 59.430 141.790 63.330 ;
        RECT 141.290 59.420 141.710 59.430 ;
        RECT 141.350 59.410 141.710 59.420 ;
        RECT 141.480 59.370 141.710 59.410 ;
        RECT 138.330 58.980 140.290 59.210 ;
        RECT 140.720 59.050 141.040 59.290 ;
        RECT 142.050 59.210 143.420 63.530 ;
        RECT 146.760 63.480 148.110 63.570 ;
        RECT 147.710 63.475 148.000 63.480 ;
        RECT 143.770 63.190 144.000 63.370 ;
        RECT 145.410 63.320 145.640 63.380 ;
        RECT 145.850 63.320 146.080 63.380 ;
        RECT 144.660 63.310 145.640 63.320 ;
        RECT 144.230 63.190 145.640 63.310 ;
        RECT 143.770 62.440 145.640 63.190 ;
        RECT 145.830 63.180 146.230 63.320 ;
        RECT 148.360 63.270 148.730 64.010 ;
        RECT 147.520 63.180 147.750 63.270 ;
        RECT 145.830 62.450 147.790 63.180 ;
        RECT 145.830 62.440 146.230 62.450 ;
        RECT 143.770 61.980 145.130 62.440 ;
        RECT 145.410 62.380 145.640 62.440 ;
        RECT 145.850 62.380 146.080 62.440 ;
        RECT 143.770 61.710 146.230 61.980 ;
        RECT 143.770 61.670 145.940 61.710 ;
        RECT 143.770 59.920 145.120 61.670 ;
        RECT 146.400 61.490 147.780 62.450 ;
        RECT 146.400 61.360 147.800 61.490 ;
        RECT 145.680 60.360 147.800 61.360 ;
        RECT 146.400 60.330 147.800 60.360 ;
        RECT 147.520 60.320 147.800 60.330 ;
        RECT 147.960 60.330 148.730 63.270 ;
        RECT 147.520 60.270 147.750 60.320 ;
        RECT 147.960 60.270 148.190 60.330 ;
        RECT 143.770 59.600 146.470 59.920 ;
        RECT 143.770 59.370 144.000 59.600 ;
        RECT 140.680 58.750 141.040 59.050 ;
        RECT 141.760 58.980 143.720 59.210 ;
        RECT 144.380 58.750 146.470 59.600 ;
        RECT 90.100 58.730 101.460 58.750 ;
        RECT 74.560 58.710 101.460 58.730 ;
        RECT 105.110 58.710 116.470 58.750 ;
        RECT 74.560 58.680 116.470 58.710 ;
        RECT 120.120 58.720 131.480 58.750 ;
        RECT 135.110 58.720 146.470 58.750 ;
        RECT 120.120 58.680 146.470 58.720 ;
        RECT 74.560 58.070 146.470 58.680 ;
        RECT 75.090 58.000 146.470 58.070 ;
        RECT 75.090 57.940 86.470 58.000 ;
        RECT 90.070 57.990 146.460 58.000 ;
        RECT 90.070 57.980 131.470 57.990 ;
        RECT 90.070 57.920 101.450 57.980 ;
        RECT 105.080 57.950 131.470 57.980 ;
        RECT 105.080 57.920 116.460 57.950 ;
        RECT 120.090 57.920 131.470 57.950 ;
        RECT 135.080 57.920 146.460 57.990 ;
        RECT 73.230 57.100 74.070 57.710 ;
        RECT 132.390 57.500 135.520 57.510 ;
        RECT 75.090 57.430 87.940 57.480 ;
        RECT 117.240 57.470 120.370 57.490 ;
        RECT 132.390 57.470 147.950 57.500 ;
        RECT 90.070 57.430 147.950 57.470 ;
        RECT 75.090 57.370 147.950 57.430 ;
        RECT 73.220 56.420 74.080 57.100 ;
        RECT 75.090 56.560 147.980 57.370 ;
        RECT 75.090 56.540 132.970 56.560 ;
        RECT 135.100 56.540 147.980 56.560 ;
        RECT 75.090 56.520 117.990 56.540 ;
        RECT 73.230 55.870 74.070 56.420 ;
        RECT 75.900 56.160 76.860 56.190 ;
        RECT 72.290 55.575 72.540 55.590 ;
        RECT 55.340 53.250 56.570 53.700 ;
        RECT 56.790 53.250 58.120 53.790 ;
        RECT 58.300 53.250 59.610 53.790 ;
        RECT 59.770 53.250 61.100 53.790 ;
        RECT 61.260 53.780 62.300 54.920 ;
        RECT 62.740 54.910 64.020 55.420 ;
        RECT 64.220 54.920 65.530 55.430 ;
        RECT 73.080 55.560 74.070 55.870 ;
        RECT 75.570 55.960 76.860 56.160 ;
        RECT 75.570 55.720 76.630 55.960 ;
        RECT 77.130 55.755 77.350 56.520 ;
        RECT 86.830 56.510 102.950 56.520 ;
        RECT 105.110 56.510 117.990 56.520 ;
        RECT 120.090 56.510 132.970 56.540 ;
        RECT 86.830 56.480 90.490 56.510 ;
        RECT 78.330 55.960 80.290 56.190 ;
        RECT 81.760 55.960 83.720 56.190 ;
        RECT 85.190 55.960 86.150 56.190 ;
        RECT 72.290 54.970 72.540 54.985 ;
        RECT 73.080 54.970 73.320 55.560 ;
        RECT 62.740 53.780 63.780 54.910 ;
        RECT 61.260 53.250 62.530 53.780 ;
        RECT 55.890 52.690 56.570 53.250 ;
        RECT 57.440 52.700 58.120 53.250 ;
        RECT 58.930 52.710 59.610 53.250 ;
        RECT 60.420 52.710 61.100 53.250 ;
        RECT 61.850 52.710 62.530 53.250 ;
        RECT 62.740 53.240 64.040 53.780 ;
        RECT 64.220 53.250 65.260 54.920 ;
        RECT 72.270 54.680 73.320 54.970 ;
        RECT 63.360 52.710 64.040 53.240 ;
        RECT 72.270 52.890 73.260 54.680 ;
        RECT 73.770 54.240 74.020 54.985 ;
        RECT 73.450 53.160 74.080 54.240 ;
        RECT 72.290 52.880 72.540 52.890 ;
        RECT 54.670 50.540 55.690 52.690 ;
        RECT 55.890 52.120 57.200 52.690 ;
        RECT 57.440 52.210 58.650 52.700 ;
        RECT 58.930 52.210 60.160 52.710 ;
        RECT 60.420 52.210 61.630 52.710 ;
        RECT 54.700 49.525 55.070 50.540 ;
        RECT 56.160 50.530 57.200 52.120 ;
        RECT 57.610 50.520 58.650 52.210 ;
        RECT 59.120 50.530 60.160 52.210 ;
        RECT 60.590 50.530 61.630 52.210 ;
        RECT 61.850 52.200 63.120 52.710 ;
        RECT 63.360 52.200 64.590 52.710 ;
        RECT 73.450 52.480 74.380 53.160 ;
        RECT 73.450 52.400 74.080 52.480 ;
        RECT 72.500 52.370 74.080 52.400 ;
        RECT 62.080 50.530 63.120 52.200 ;
        RECT 63.550 50.530 64.590 52.200 ;
        RECT 72.270 52.100 74.080 52.370 ;
        RECT 72.270 52.020 73.870 52.100 ;
        RECT 72.270 50.070 72.760 52.020 ;
        RECT 73.770 51.590 74.020 51.690 ;
        RECT 73.090 50.920 74.060 51.590 ;
        RECT 73.090 50.240 74.080 50.920 ;
        RECT 72.290 49.585 72.540 50.070 ;
        RECT 73.090 49.810 74.060 50.240 ;
        RECT 72.930 49.660 74.060 49.810 ;
        RECT 54.700 49.155 68.315 49.525 ;
        RECT 54.730 48.340 67.580 48.470 ;
        RECT 54.730 47.510 67.610 48.340 ;
        RECT 55.540 46.950 56.500 47.180 ;
        RECT 55.260 46.710 55.490 46.745 ;
        RECT 55.160 39.600 55.490 46.710 ;
        RECT 55.150 38.745 55.490 39.600 ;
        RECT 55.150 38.740 55.470 38.745 ;
        RECT 55.150 38.160 55.390 38.740 ;
        RECT 55.800 38.540 56.270 46.950 ;
        RECT 56.770 46.745 56.990 47.510 ;
        RECT 57.970 46.950 59.930 47.180 ;
        RECT 61.400 46.950 63.360 47.180 ;
        RECT 64.830 46.950 65.790 47.180 ;
        RECT 56.550 46.540 56.990 46.745 ;
        RECT 57.690 46.720 57.920 46.745 ;
        RECT 57.690 46.710 57.930 46.720 ;
        RECT 56.550 38.800 56.940 46.540 ;
        RECT 57.520 39.650 57.930 46.710 ;
        RECT 58.510 40.360 59.410 46.950 ;
        RECT 59.980 46.700 60.210 46.745 ;
        RECT 61.120 46.720 61.350 46.745 ;
        RECT 57.510 38.830 57.930 39.650 ;
        RECT 58.480 39.350 59.480 40.360 ;
        RECT 56.550 38.745 56.780 38.800 ;
        RECT 57.510 38.745 57.920 38.830 ;
        RECT 55.540 38.310 56.500 38.540 ;
        RECT 55.150 37.670 55.470 38.160 ;
        RECT 54.710 36.420 55.550 37.670 ;
        RECT 55.150 35.370 55.390 36.420 ;
        RECT 55.690 35.760 56.360 38.310 ;
        RECT 57.510 36.530 57.830 38.745 ;
        RECT 58.510 38.540 59.410 39.350 ;
        RECT 59.980 38.810 60.500 46.700 ;
        RECT 59.980 38.745 60.210 38.810 ;
        RECT 60.980 38.800 61.360 46.720 ;
        RECT 62.060 40.320 62.880 46.950 ;
        RECT 63.410 46.700 63.640 46.745 ;
        RECT 64.550 46.700 64.780 46.745 ;
        RECT 61.970 39.320 62.970 40.320 ;
        RECT 60.990 38.745 61.350 38.800 ;
        RECT 57.970 38.310 59.930 38.540 ;
        RECT 60.990 37.180 61.250 38.745 ;
        RECT 62.060 38.540 62.880 39.320 ;
        RECT 63.410 38.830 64.790 46.700 ;
        RECT 65.140 46.580 65.560 46.950 ;
        RECT 65.840 46.700 66.070 46.745 ;
        RECT 66.470 46.700 67.610 47.510 ;
        RECT 65.840 42.720 67.610 46.700 ;
        RECT 65.840 41.720 67.600 42.720 ;
        RECT 63.410 38.745 63.640 38.830 ;
        RECT 64.550 38.745 64.780 38.830 ;
        RECT 65.140 38.540 65.560 39.210 ;
        RECT 65.840 38.840 67.610 41.720 ;
        RECT 65.840 38.745 66.070 38.840 ;
        RECT 61.400 38.310 63.360 38.540 ;
        RECT 64.830 38.310 65.790 38.540 ;
        RECT 64.930 37.430 65.720 38.310 ;
        RECT 66.470 37.830 67.610 38.840 ;
        RECT 60.990 36.560 64.610 37.180 ;
        RECT 64.880 36.670 65.770 37.430 ;
        RECT 55.550 35.530 56.510 35.760 ;
        RECT 55.150 34.360 55.500 35.370 ;
        RECT 55.160 31.410 55.500 34.360 ;
        RECT 55.270 31.370 55.500 31.410 ;
        RECT 55.800 31.210 56.240 35.530 ;
        RECT 57.510 35.370 57.840 36.530 ;
        RECT 57.980 35.530 59.940 35.760 ;
        RECT 56.560 35.360 56.790 35.370 ;
        RECT 56.560 33.050 56.970 35.360 ;
        RECT 57.510 35.330 57.930 35.370 ;
        RECT 58.290 35.330 59.630 35.530 ;
        RECT 60.990 35.370 61.250 36.560 ;
        RECT 64.200 35.910 64.600 36.560 ;
        RECT 66.540 36.280 67.610 37.830 ;
        RECT 67.945 37.475 68.315 49.155 ;
        RECT 72.290 48.990 72.540 48.995 ;
        RECT 72.930 48.990 73.280 49.660 ;
        RECT 73.770 49.585 74.020 49.660 ;
        RECT 72.280 48.760 73.280 48.990 ;
        RECT 72.280 47.200 73.250 48.760 ;
        RECT 73.770 48.630 74.020 48.995 ;
        RECT 73.470 47.750 74.040 48.630 ;
        RECT 75.520 48.610 76.630 55.720 ;
        RECT 72.290 46.890 72.540 47.200 ;
        RECT 73.470 46.940 74.490 47.750 ;
        RECT 75.510 47.550 76.630 48.610 ;
        RECT 76.910 55.550 77.350 55.755 ;
        RECT 78.050 55.730 78.280 55.755 ;
        RECT 78.050 55.720 78.290 55.730 ;
        RECT 76.910 47.810 77.300 55.550 ;
        RECT 77.880 48.660 78.290 55.720 ;
        RECT 78.870 49.370 79.770 55.960 ;
        RECT 80.340 55.710 80.570 55.755 ;
        RECT 81.480 55.730 81.710 55.755 ;
        RECT 77.870 47.840 78.290 48.660 ;
        RECT 78.840 48.360 79.840 49.370 ;
        RECT 76.910 47.755 77.140 47.810 ;
        RECT 77.870 47.755 78.280 47.840 ;
        RECT 75.510 47.320 76.860 47.550 ;
        RECT 73.470 46.420 74.040 46.940 ;
        RECT 75.510 46.680 76.720 47.320 ;
        RECT 72.680 46.350 74.040 46.420 ;
        RECT 72.270 46.120 74.040 46.350 ;
        RECT 72.270 46.010 73.650 46.120 ;
        RECT 72.270 44.330 73.050 46.010 ;
        RECT 73.770 45.690 74.020 45.700 ;
        RECT 73.430 45.020 74.020 45.690 ;
        RECT 75.070 45.430 76.720 46.680 ;
        RECT 72.270 43.580 72.860 44.330 ;
        RECT 73.430 44.210 74.410 45.020 ;
        RECT 73.430 43.930 74.020 44.210 ;
        RECT 73.150 43.590 74.020 43.930 ;
        RECT 73.150 43.200 73.500 43.590 ;
        RECT 72.800 43.120 73.500 43.200 ;
        RECT 72.800 43.070 73.370 43.120 ;
        RECT 72.290 42.970 72.540 43.005 ;
        RECT 72.690 42.970 73.370 43.070 ;
        RECT 72.260 42.900 73.370 42.970 ;
        RECT 72.260 42.810 72.950 42.900 ;
        RECT 72.260 40.870 72.850 42.810 ;
        RECT 73.770 42.550 74.020 43.005 ;
        RECT 73.300 41.300 74.080 42.550 ;
        RECT 73.180 40.840 74.080 41.300 ;
        RECT 73.180 40.390 73.410 40.840 ;
        RECT 72.970 40.310 73.410 40.390 ;
        RECT 72.240 39.850 73.410 40.310 ;
        RECT 72.240 39.600 73.270 39.850 ;
        RECT 74.550 39.760 75.260 45.250 ;
        RECT 75.510 44.770 76.720 45.430 ;
        RECT 77.870 45.540 78.190 47.755 ;
        RECT 78.870 47.550 79.770 48.360 ;
        RECT 80.340 47.820 80.860 55.710 ;
        RECT 80.340 47.755 80.570 47.820 ;
        RECT 81.340 47.810 81.720 55.730 ;
        RECT 82.350 55.280 83.320 55.960 ;
        RECT 82.340 55.260 83.320 55.280 ;
        RECT 83.770 55.710 84.000 55.755 ;
        RECT 84.910 55.710 85.140 55.755 ;
        RECT 82.340 54.350 83.310 55.260 ;
        RECT 82.420 49.330 83.240 54.350 ;
        RECT 82.330 48.330 83.330 49.330 ;
        RECT 81.350 47.755 81.710 47.810 ;
        RECT 78.330 47.320 80.290 47.550 ;
        RECT 81.350 46.190 81.610 47.755 ;
        RECT 82.420 47.550 83.240 48.330 ;
        RECT 83.770 47.840 85.150 55.710 ;
        RECT 85.480 55.590 85.920 55.960 ;
        RECT 86.200 55.710 86.430 55.755 ;
        RECT 86.830 55.710 88.440 56.480 ;
        RECT 90.880 56.150 91.840 56.180 ;
        RECT 90.550 55.950 91.840 56.150 ;
        RECT 90.550 55.710 91.610 55.950 ;
        RECT 92.110 55.745 92.330 56.510 ;
        RECT 93.310 55.950 95.270 56.180 ;
        RECT 96.740 55.950 98.700 56.180 ;
        RECT 100.170 55.950 101.130 56.180 ;
        RECT 85.480 48.220 85.910 55.590 ;
        RECT 86.200 55.510 88.440 55.710 ;
        RECT 86.200 51.730 87.970 55.510 ;
        RECT 86.200 50.730 87.960 51.730 ;
        RECT 83.770 47.755 84.000 47.840 ;
        RECT 84.910 47.755 85.140 47.840 ;
        RECT 85.480 47.550 85.920 48.220 ;
        RECT 86.200 47.850 87.970 50.730 ;
        RECT 90.500 48.600 91.610 55.710 ;
        RECT 86.200 47.755 86.430 47.850 ;
        RECT 81.760 47.320 83.720 47.550 ;
        RECT 85.190 47.320 86.150 47.550 ;
        RECT 85.290 46.440 86.080 47.320 ;
        RECT 86.830 46.840 87.970 47.850 ;
        RECT 81.350 45.570 84.970 46.190 ;
        RECT 85.240 45.680 86.130 46.440 ;
        RECT 75.510 44.540 76.870 44.770 ;
        RECT 75.510 43.370 76.600 44.540 ;
        RECT 77.870 44.380 78.200 45.540 ;
        RECT 78.340 44.540 80.300 44.770 ;
        RECT 75.520 40.420 76.600 43.370 ;
        RECT 75.570 40.220 76.600 40.420 ;
        RECT 76.920 44.370 77.150 44.380 ;
        RECT 76.920 42.060 77.330 44.370 ;
        RECT 77.870 44.360 78.290 44.380 ;
        RECT 77.870 44.310 78.380 44.360 ;
        RECT 78.730 44.310 79.990 44.540 ;
        RECT 81.350 44.380 81.610 45.570 ;
        RECT 84.560 44.920 84.960 45.570 ;
        RECT 86.900 45.520 87.970 46.840 ;
        RECT 90.490 47.540 91.610 48.600 ;
        RECT 91.890 55.540 92.330 55.745 ;
        RECT 93.030 55.720 93.260 55.745 ;
        RECT 93.030 55.710 93.270 55.720 ;
        RECT 91.890 47.800 92.280 55.540 ;
        RECT 92.860 48.650 93.270 55.710 ;
        RECT 93.850 49.360 94.750 55.950 ;
        RECT 95.320 55.700 95.550 55.745 ;
        RECT 96.460 55.720 96.690 55.745 ;
        RECT 92.850 47.830 93.270 48.650 ;
        RECT 93.820 48.350 94.820 49.360 ;
        RECT 91.890 47.745 92.120 47.800 ;
        RECT 92.850 47.745 93.260 47.830 ;
        RECT 90.490 47.310 91.840 47.540 ;
        RECT 90.490 46.670 91.700 47.310 ;
        RECT 86.900 45.020 88.740 45.520 ;
        RECT 90.050 45.420 91.700 46.670 ;
        RECT 85.960 44.920 86.710 44.930 ;
        RECT 84.560 44.870 86.710 44.920 ;
        RECT 84.560 44.830 86.890 44.870 ;
        RECT 81.770 44.540 83.730 44.770 ;
        RECT 84.560 44.580 88.120 44.830 ;
        RECT 84.560 44.570 85.900 44.580 ;
        RECT 85.610 44.550 85.900 44.570 ;
        RECT 76.920 40.380 77.420 42.060 ;
        RECT 77.870 40.450 79.990 44.310 ;
        RECT 77.990 40.440 79.990 40.450 ;
        RECT 78.060 40.380 78.290 40.440 ;
        RECT 75.570 40.040 76.870 40.220 ;
        RECT 75.910 39.990 76.870 40.040 ;
        RECT 77.220 39.760 77.420 40.380 ;
        RECT 78.650 40.220 79.990 40.440 ;
        RECT 80.350 44.340 80.580 44.380 ;
        RECT 81.350 44.350 81.720 44.380 ;
        RECT 81.350 44.340 81.800 44.350 ;
        RECT 80.350 44.330 80.760 44.340 ;
        RECT 80.350 42.110 80.800 44.330 ;
        RECT 80.350 41.620 80.850 42.110 ;
        RECT 80.350 40.950 80.940 41.620 ;
        RECT 80.350 40.700 81.000 40.950 ;
        RECT 80.350 40.670 81.050 40.700 ;
        RECT 80.350 40.380 80.580 40.670 ;
        RECT 80.810 40.300 81.050 40.670 ;
        RECT 81.300 40.440 81.800 44.340 ;
        RECT 81.300 40.430 81.720 40.440 ;
        RECT 81.360 40.420 81.720 40.430 ;
        RECT 81.490 40.380 81.720 40.420 ;
        RECT 78.340 39.990 80.300 40.220 ;
        RECT 80.730 40.060 81.050 40.300 ;
        RECT 82.060 40.220 83.430 44.540 ;
        RECT 86.770 44.490 88.120 44.580 ;
        RECT 87.720 44.485 88.010 44.490 ;
        RECT 83.780 44.200 84.010 44.380 ;
        RECT 85.420 44.330 85.650 44.390 ;
        RECT 85.860 44.330 86.090 44.390 ;
        RECT 84.670 44.320 85.650 44.330 ;
        RECT 84.240 44.200 85.650 44.320 ;
        RECT 83.780 43.450 85.650 44.200 ;
        RECT 85.840 44.190 86.240 44.330 ;
        RECT 88.370 44.280 88.740 45.020 ;
        RECT 87.530 44.190 87.760 44.280 ;
        RECT 85.840 43.460 87.800 44.190 ;
        RECT 85.840 43.450 86.240 43.460 ;
        RECT 83.780 42.990 85.140 43.450 ;
        RECT 85.420 43.390 85.650 43.450 ;
        RECT 85.860 43.390 86.090 43.450 ;
        RECT 83.780 42.720 86.240 42.990 ;
        RECT 83.780 42.680 85.950 42.720 ;
        RECT 83.780 40.930 85.130 42.680 ;
        RECT 86.410 42.500 87.790 43.460 ;
        RECT 86.410 42.370 87.810 42.500 ;
        RECT 85.690 41.370 87.810 42.370 ;
        RECT 86.410 41.340 87.810 41.370 ;
        RECT 87.530 41.330 87.810 41.340 ;
        RECT 87.970 41.340 88.740 44.280 ;
        RECT 90.490 44.760 91.700 45.420 ;
        RECT 92.850 45.530 93.170 47.745 ;
        RECT 93.850 47.540 94.750 48.350 ;
        RECT 95.320 47.810 95.840 55.700 ;
        RECT 95.320 47.745 95.550 47.810 ;
        RECT 96.320 47.800 96.700 55.720 ;
        RECT 97.400 49.320 98.220 55.950 ;
        RECT 98.750 55.700 98.980 55.745 ;
        RECT 99.890 55.700 100.120 55.745 ;
        RECT 97.310 48.320 98.310 49.320 ;
        RECT 96.330 47.745 96.690 47.800 ;
        RECT 93.310 47.310 95.270 47.540 ;
        RECT 96.330 46.180 96.590 47.745 ;
        RECT 97.400 47.540 98.220 48.320 ;
        RECT 98.750 47.830 100.130 55.700 ;
        RECT 100.460 55.580 100.900 55.950 ;
        RECT 101.180 55.700 101.410 55.745 ;
        RECT 101.810 55.700 102.950 56.510 ;
        RECT 105.920 56.150 106.880 56.180 ;
        RECT 105.590 55.950 106.880 56.150 ;
        RECT 105.590 55.710 106.650 55.950 ;
        RECT 107.150 55.745 107.370 56.510 ;
        RECT 108.350 55.950 110.310 56.180 ;
        RECT 111.780 55.950 113.740 56.180 ;
        RECT 115.210 55.950 116.170 56.180 ;
        RECT 100.460 48.210 100.890 55.580 ;
        RECT 101.180 51.720 102.950 55.700 ;
        RECT 101.180 50.720 102.940 51.720 ;
        RECT 98.750 47.745 98.980 47.830 ;
        RECT 99.890 47.745 100.120 47.830 ;
        RECT 100.460 47.540 100.900 48.210 ;
        RECT 101.180 47.840 102.950 50.720 ;
        RECT 105.540 48.600 106.650 55.710 ;
        RECT 101.180 47.745 101.410 47.840 ;
        RECT 96.740 47.310 98.700 47.540 ;
        RECT 100.170 47.310 101.130 47.540 ;
        RECT 100.270 46.430 101.060 47.310 ;
        RECT 101.810 46.830 102.950 47.840 ;
        RECT 96.330 45.560 99.950 46.180 ;
        RECT 100.220 45.670 101.110 46.430 ;
        RECT 90.490 44.530 91.850 44.760 ;
        RECT 90.490 43.360 91.580 44.530 ;
        RECT 92.850 44.370 93.180 45.530 ;
        RECT 93.320 44.530 95.280 44.760 ;
        RECT 87.530 41.280 87.760 41.330 ;
        RECT 87.970 41.280 88.200 41.340 ;
        RECT 83.780 40.610 86.480 40.930 ;
        RECT 83.780 40.380 84.010 40.610 ;
        RECT 80.690 39.760 81.050 40.060 ;
        RECT 81.770 39.990 83.730 40.220 ;
        RECT 84.390 39.760 86.480 40.610 ;
        RECT 90.500 40.410 91.580 43.360 ;
        RECT 90.550 40.210 91.580 40.410 ;
        RECT 91.900 44.360 92.130 44.370 ;
        RECT 91.900 42.050 92.310 44.360 ;
        RECT 92.850 44.350 93.270 44.370 ;
        RECT 92.850 44.300 93.360 44.350 ;
        RECT 93.710 44.300 94.970 44.530 ;
        RECT 96.330 44.370 96.590 45.560 ;
        RECT 99.540 44.910 99.940 45.560 ;
        RECT 101.880 45.510 102.950 46.830 ;
        RECT 105.530 47.540 106.650 48.600 ;
        RECT 106.930 55.540 107.370 55.745 ;
        RECT 108.070 55.720 108.300 55.745 ;
        RECT 108.070 55.710 108.310 55.720 ;
        RECT 106.930 47.800 107.320 55.540 ;
        RECT 107.900 48.650 108.310 55.710 ;
        RECT 108.890 49.360 109.790 55.950 ;
        RECT 110.360 55.700 110.590 55.745 ;
        RECT 111.500 55.720 111.730 55.745 ;
        RECT 107.890 47.830 108.310 48.650 ;
        RECT 108.860 48.350 109.860 49.360 ;
        RECT 106.930 47.745 107.160 47.800 ;
        RECT 107.890 47.745 108.300 47.830 ;
        RECT 105.530 47.310 106.880 47.540 ;
        RECT 105.530 46.670 106.740 47.310 ;
        RECT 101.880 45.010 103.720 45.510 ;
        RECT 105.090 45.420 106.740 46.670 ;
        RECT 100.940 44.910 101.690 44.920 ;
        RECT 99.540 44.860 101.690 44.910 ;
        RECT 99.540 44.820 101.870 44.860 ;
        RECT 96.750 44.530 98.710 44.760 ;
        RECT 99.540 44.570 103.100 44.820 ;
        RECT 99.540 44.560 100.880 44.570 ;
        RECT 100.590 44.540 100.880 44.560 ;
        RECT 91.900 40.370 92.400 42.050 ;
        RECT 92.850 40.440 94.970 44.300 ;
        RECT 92.970 40.430 94.970 40.440 ;
        RECT 93.040 40.370 93.270 40.430 ;
        RECT 90.550 40.030 91.850 40.210 ;
        RECT 90.890 39.980 91.850 40.030 ;
        RECT 74.550 39.710 86.480 39.760 ;
        RECT 92.200 39.750 92.400 40.370 ;
        RECT 93.630 40.210 94.970 40.430 ;
        RECT 95.330 44.330 95.560 44.370 ;
        RECT 96.330 44.340 96.700 44.370 ;
        RECT 96.330 44.330 96.780 44.340 ;
        RECT 95.330 44.320 95.740 44.330 ;
        RECT 95.330 42.100 95.780 44.320 ;
        RECT 95.330 41.610 95.830 42.100 ;
        RECT 95.330 40.940 95.920 41.610 ;
        RECT 95.330 40.690 95.980 40.940 ;
        RECT 95.330 40.660 96.030 40.690 ;
        RECT 95.330 40.370 95.560 40.660 ;
        RECT 95.790 40.290 96.030 40.660 ;
        RECT 96.280 40.430 96.780 44.330 ;
        RECT 96.280 40.420 96.700 40.430 ;
        RECT 96.340 40.410 96.700 40.420 ;
        RECT 96.470 40.370 96.700 40.410 ;
        RECT 93.320 39.980 95.280 40.210 ;
        RECT 95.710 40.050 96.030 40.290 ;
        RECT 97.040 40.210 98.410 44.530 ;
        RECT 101.750 44.480 103.100 44.570 ;
        RECT 102.700 44.475 102.990 44.480 ;
        RECT 98.760 44.190 98.990 44.370 ;
        RECT 100.400 44.320 100.630 44.380 ;
        RECT 100.840 44.320 101.070 44.380 ;
        RECT 99.650 44.310 100.630 44.320 ;
        RECT 99.220 44.190 100.630 44.310 ;
        RECT 98.760 43.440 100.630 44.190 ;
        RECT 100.820 44.180 101.220 44.320 ;
        RECT 103.350 44.270 103.720 45.010 ;
        RECT 102.510 44.180 102.740 44.270 ;
        RECT 100.820 43.450 102.780 44.180 ;
        RECT 100.820 43.440 101.220 43.450 ;
        RECT 98.760 42.980 100.120 43.440 ;
        RECT 100.400 43.380 100.630 43.440 ;
        RECT 100.840 43.380 101.070 43.440 ;
        RECT 98.760 42.710 101.220 42.980 ;
        RECT 98.760 42.670 100.930 42.710 ;
        RECT 98.760 40.920 100.110 42.670 ;
        RECT 101.390 42.490 102.770 43.450 ;
        RECT 101.390 42.360 102.790 42.490 ;
        RECT 100.670 41.360 102.790 42.360 ;
        RECT 101.390 41.330 102.790 41.360 ;
        RECT 102.510 41.320 102.790 41.330 ;
        RECT 102.950 41.330 103.720 44.270 ;
        RECT 105.530 44.760 106.740 45.420 ;
        RECT 107.890 45.530 108.210 47.745 ;
        RECT 108.890 47.540 109.790 48.350 ;
        RECT 110.360 47.810 110.880 55.700 ;
        RECT 110.360 47.745 110.590 47.810 ;
        RECT 111.360 47.800 111.740 55.720 ;
        RECT 112.440 49.320 113.260 55.950 ;
        RECT 113.790 55.700 114.020 55.745 ;
        RECT 114.930 55.700 115.160 55.745 ;
        RECT 112.350 48.320 113.350 49.320 ;
        RECT 111.370 47.745 111.730 47.800 ;
        RECT 108.350 47.310 110.310 47.540 ;
        RECT 111.370 46.180 111.630 47.745 ;
        RECT 112.440 47.540 113.260 48.320 ;
        RECT 113.790 47.830 115.170 55.700 ;
        RECT 115.500 55.580 115.940 55.950 ;
        RECT 116.220 55.700 116.450 55.745 ;
        RECT 116.850 55.700 117.990 56.510 ;
        RECT 120.900 56.150 121.860 56.180 ;
        RECT 120.570 55.950 121.860 56.150 ;
        RECT 120.570 55.710 121.630 55.950 ;
        RECT 122.130 55.745 122.350 56.510 ;
        RECT 123.330 55.950 125.290 56.180 ;
        RECT 126.760 55.950 128.720 56.180 ;
        RECT 130.190 55.950 131.150 56.180 ;
        RECT 115.500 48.210 115.930 55.580 ;
        RECT 116.220 51.720 117.990 55.700 ;
        RECT 116.220 50.720 117.980 51.720 ;
        RECT 113.790 47.745 114.020 47.830 ;
        RECT 114.930 47.745 115.160 47.830 ;
        RECT 115.500 47.540 115.940 48.210 ;
        RECT 116.220 47.840 117.990 50.720 ;
        RECT 120.520 48.600 121.630 55.710 ;
        RECT 116.220 47.745 116.450 47.840 ;
        RECT 111.780 47.310 113.740 47.540 ;
        RECT 115.210 47.310 116.170 47.540 ;
        RECT 115.310 46.430 116.100 47.310 ;
        RECT 116.850 46.830 117.990 47.840 ;
        RECT 111.370 45.560 114.990 46.180 ;
        RECT 115.260 45.670 116.150 46.430 ;
        RECT 105.530 44.530 106.890 44.760 ;
        RECT 105.530 43.360 106.620 44.530 ;
        RECT 107.890 44.370 108.220 45.530 ;
        RECT 108.360 44.530 110.320 44.760 ;
        RECT 102.510 41.270 102.740 41.320 ;
        RECT 102.950 41.270 103.180 41.330 ;
        RECT 98.760 40.600 101.460 40.920 ;
        RECT 98.760 40.370 98.990 40.600 ;
        RECT 95.670 39.750 96.030 40.050 ;
        RECT 96.750 39.980 98.710 40.210 ;
        RECT 99.370 39.750 101.460 40.600 ;
        RECT 105.540 40.410 106.620 43.360 ;
        RECT 105.590 40.210 106.620 40.410 ;
        RECT 106.940 44.360 107.170 44.370 ;
        RECT 106.940 42.050 107.350 44.360 ;
        RECT 107.890 44.350 108.310 44.370 ;
        RECT 107.890 44.300 108.400 44.350 ;
        RECT 108.750 44.300 110.010 44.530 ;
        RECT 111.370 44.370 111.630 45.560 ;
        RECT 114.580 44.910 114.980 45.560 ;
        RECT 116.920 45.510 117.990 46.830 ;
        RECT 120.510 47.540 121.630 48.600 ;
        RECT 121.910 55.540 122.350 55.745 ;
        RECT 123.050 55.720 123.280 55.745 ;
        RECT 123.050 55.710 123.290 55.720 ;
        RECT 121.910 47.800 122.300 55.540 ;
        RECT 122.880 48.650 123.290 55.710 ;
        RECT 123.870 49.360 124.770 55.950 ;
        RECT 125.340 55.700 125.570 55.745 ;
        RECT 126.480 55.720 126.710 55.745 ;
        RECT 122.870 47.830 123.290 48.650 ;
        RECT 123.840 48.350 124.840 49.360 ;
        RECT 121.910 47.745 122.140 47.800 ;
        RECT 122.870 47.745 123.280 47.830 ;
        RECT 120.510 47.310 121.860 47.540 ;
        RECT 120.510 46.670 121.720 47.310 ;
        RECT 116.920 45.010 118.760 45.510 ;
        RECT 120.070 45.420 121.720 46.670 ;
        RECT 115.980 44.910 116.730 44.920 ;
        RECT 114.580 44.860 116.730 44.910 ;
        RECT 114.580 44.820 116.910 44.860 ;
        RECT 111.790 44.530 113.750 44.760 ;
        RECT 114.580 44.570 118.140 44.820 ;
        RECT 114.580 44.560 115.920 44.570 ;
        RECT 115.630 44.540 115.920 44.560 ;
        RECT 106.940 40.370 107.440 42.050 ;
        RECT 107.890 40.440 110.010 44.300 ;
        RECT 108.010 40.430 110.010 40.440 ;
        RECT 108.080 40.370 108.310 40.430 ;
        RECT 105.590 40.030 106.890 40.210 ;
        RECT 105.930 39.980 106.890 40.030 ;
        RECT 107.240 39.750 107.440 40.370 ;
        RECT 108.670 40.210 110.010 40.430 ;
        RECT 110.370 44.330 110.600 44.370 ;
        RECT 111.370 44.340 111.740 44.370 ;
        RECT 111.370 44.330 111.820 44.340 ;
        RECT 110.370 44.320 110.780 44.330 ;
        RECT 110.370 42.100 110.820 44.320 ;
        RECT 110.370 41.610 110.870 42.100 ;
        RECT 110.370 40.940 110.960 41.610 ;
        RECT 110.370 40.690 111.020 40.940 ;
        RECT 110.370 40.660 111.070 40.690 ;
        RECT 110.370 40.370 110.600 40.660 ;
        RECT 110.830 40.290 111.070 40.660 ;
        RECT 111.320 40.430 111.820 44.330 ;
        RECT 111.320 40.420 111.740 40.430 ;
        RECT 111.380 40.410 111.740 40.420 ;
        RECT 111.510 40.370 111.740 40.410 ;
        RECT 108.360 39.980 110.320 40.210 ;
        RECT 110.750 40.050 111.070 40.290 ;
        RECT 112.080 40.210 113.450 44.530 ;
        RECT 116.790 44.480 118.140 44.570 ;
        RECT 117.740 44.475 118.030 44.480 ;
        RECT 113.800 44.190 114.030 44.370 ;
        RECT 115.440 44.320 115.670 44.380 ;
        RECT 115.880 44.320 116.110 44.380 ;
        RECT 114.690 44.310 115.670 44.320 ;
        RECT 114.260 44.190 115.670 44.310 ;
        RECT 113.800 43.440 115.670 44.190 ;
        RECT 115.860 44.180 116.260 44.320 ;
        RECT 118.390 44.270 118.760 45.010 ;
        RECT 117.550 44.180 117.780 44.270 ;
        RECT 115.860 43.450 117.820 44.180 ;
        RECT 115.860 43.440 116.260 43.450 ;
        RECT 113.800 42.980 115.160 43.440 ;
        RECT 115.440 43.380 115.670 43.440 ;
        RECT 115.880 43.380 116.110 43.440 ;
        RECT 113.800 42.710 116.260 42.980 ;
        RECT 113.800 42.670 115.970 42.710 ;
        RECT 113.800 40.920 115.150 42.670 ;
        RECT 116.430 42.490 117.810 43.450 ;
        RECT 116.430 42.360 117.830 42.490 ;
        RECT 115.710 41.360 117.830 42.360 ;
        RECT 116.430 41.330 117.830 41.360 ;
        RECT 117.550 41.320 117.830 41.330 ;
        RECT 117.990 41.330 118.760 44.270 ;
        RECT 120.510 44.760 121.720 45.420 ;
        RECT 122.870 45.530 123.190 47.745 ;
        RECT 123.870 47.540 124.770 48.350 ;
        RECT 125.340 47.810 125.860 55.700 ;
        RECT 125.340 47.745 125.570 47.810 ;
        RECT 126.340 47.800 126.720 55.720 ;
        RECT 127.420 49.320 128.240 55.950 ;
        RECT 128.770 55.700 129.000 55.745 ;
        RECT 129.910 55.700 130.140 55.745 ;
        RECT 127.330 48.320 128.330 49.320 ;
        RECT 126.350 47.745 126.710 47.800 ;
        RECT 123.330 47.310 125.290 47.540 ;
        RECT 126.350 46.180 126.610 47.745 ;
        RECT 127.420 47.540 128.240 48.320 ;
        RECT 128.770 47.830 130.150 55.700 ;
        RECT 130.480 55.580 130.920 55.950 ;
        RECT 131.200 55.700 131.430 55.745 ;
        RECT 131.830 55.700 132.970 56.510 ;
        RECT 135.910 56.180 136.870 56.210 ;
        RECT 135.580 55.980 136.870 56.180 ;
        RECT 135.580 55.740 136.640 55.980 ;
        RECT 137.140 55.775 137.360 56.540 ;
        RECT 138.340 55.980 140.300 56.210 ;
        RECT 141.770 55.980 143.730 56.210 ;
        RECT 145.200 55.980 146.160 56.210 ;
        RECT 130.480 48.210 130.910 55.580 ;
        RECT 131.200 51.720 132.970 55.700 ;
        RECT 131.200 50.720 132.960 51.720 ;
        RECT 128.770 47.745 129.000 47.830 ;
        RECT 129.910 47.745 130.140 47.830 ;
        RECT 130.480 47.540 130.920 48.210 ;
        RECT 131.200 47.840 132.970 50.720 ;
        RECT 135.530 48.630 136.640 55.740 ;
        RECT 131.200 47.745 131.430 47.840 ;
        RECT 126.760 47.310 128.720 47.540 ;
        RECT 130.190 47.310 131.150 47.540 ;
        RECT 130.290 46.430 131.080 47.310 ;
        RECT 131.830 46.830 132.970 47.840 ;
        RECT 126.350 45.560 129.970 46.180 ;
        RECT 130.240 45.670 131.130 46.430 ;
        RECT 120.510 44.530 121.870 44.760 ;
        RECT 120.510 43.360 121.600 44.530 ;
        RECT 122.870 44.370 123.200 45.530 ;
        RECT 123.340 44.530 125.300 44.760 ;
        RECT 117.550 41.270 117.780 41.320 ;
        RECT 117.990 41.270 118.220 41.330 ;
        RECT 113.800 40.600 116.500 40.920 ;
        RECT 113.800 40.370 114.030 40.600 ;
        RECT 110.710 39.750 111.070 40.050 ;
        RECT 111.790 39.980 113.750 40.210 ;
        RECT 114.410 39.750 116.500 40.600 ;
        RECT 120.520 40.410 121.600 43.360 ;
        RECT 120.570 40.210 121.600 40.410 ;
        RECT 121.920 44.360 122.150 44.370 ;
        RECT 121.920 42.050 122.330 44.360 ;
        RECT 122.870 44.350 123.290 44.370 ;
        RECT 122.870 44.300 123.380 44.350 ;
        RECT 123.730 44.300 124.990 44.530 ;
        RECT 126.350 44.370 126.610 45.560 ;
        RECT 129.560 44.910 129.960 45.560 ;
        RECT 131.900 45.510 132.970 46.830 ;
        RECT 135.520 47.570 136.640 48.630 ;
        RECT 136.920 55.570 137.360 55.775 ;
        RECT 138.060 55.750 138.290 55.775 ;
        RECT 138.060 55.740 138.300 55.750 ;
        RECT 136.920 47.830 137.310 55.570 ;
        RECT 137.890 48.680 138.300 55.740 ;
        RECT 138.880 49.390 139.780 55.980 ;
        RECT 140.350 55.730 140.580 55.775 ;
        RECT 141.490 55.750 141.720 55.775 ;
        RECT 137.880 47.860 138.300 48.680 ;
        RECT 138.850 48.380 139.850 49.390 ;
        RECT 136.920 47.775 137.150 47.830 ;
        RECT 137.880 47.775 138.290 47.860 ;
        RECT 135.520 47.340 136.870 47.570 ;
        RECT 135.520 46.700 136.730 47.340 ;
        RECT 131.900 45.010 133.740 45.510 ;
        RECT 135.080 45.450 136.730 46.700 ;
        RECT 130.960 44.910 131.710 44.920 ;
        RECT 129.560 44.860 131.710 44.910 ;
        RECT 129.560 44.820 131.890 44.860 ;
        RECT 126.770 44.530 128.730 44.760 ;
        RECT 129.560 44.570 133.120 44.820 ;
        RECT 129.560 44.560 130.900 44.570 ;
        RECT 130.610 44.540 130.900 44.560 ;
        RECT 121.920 40.370 122.420 42.050 ;
        RECT 122.870 40.440 124.990 44.300 ;
        RECT 122.990 40.430 124.990 40.440 ;
        RECT 123.060 40.370 123.290 40.430 ;
        RECT 120.570 40.030 121.870 40.210 ;
        RECT 120.910 39.980 121.870 40.030 ;
        RECT 122.220 39.750 122.420 40.370 ;
        RECT 123.650 40.210 124.990 40.430 ;
        RECT 125.350 44.330 125.580 44.370 ;
        RECT 126.350 44.340 126.720 44.370 ;
        RECT 126.350 44.330 126.800 44.340 ;
        RECT 125.350 44.320 125.760 44.330 ;
        RECT 125.350 42.100 125.800 44.320 ;
        RECT 125.350 41.610 125.850 42.100 ;
        RECT 125.350 40.940 125.940 41.610 ;
        RECT 125.350 40.690 126.000 40.940 ;
        RECT 125.350 40.660 126.050 40.690 ;
        RECT 125.350 40.370 125.580 40.660 ;
        RECT 125.810 40.290 126.050 40.660 ;
        RECT 126.300 40.430 126.800 44.330 ;
        RECT 126.300 40.420 126.720 40.430 ;
        RECT 126.360 40.410 126.720 40.420 ;
        RECT 126.490 40.370 126.720 40.410 ;
        RECT 123.340 39.980 125.300 40.210 ;
        RECT 125.730 40.050 126.050 40.290 ;
        RECT 127.060 40.210 128.430 44.530 ;
        RECT 131.770 44.480 133.120 44.570 ;
        RECT 132.720 44.475 133.010 44.480 ;
        RECT 128.780 44.190 129.010 44.370 ;
        RECT 130.420 44.320 130.650 44.380 ;
        RECT 130.860 44.320 131.090 44.380 ;
        RECT 129.670 44.310 130.650 44.320 ;
        RECT 129.240 44.190 130.650 44.310 ;
        RECT 128.780 43.440 130.650 44.190 ;
        RECT 130.840 44.180 131.240 44.320 ;
        RECT 133.370 44.270 133.740 45.010 ;
        RECT 132.530 44.180 132.760 44.270 ;
        RECT 130.840 43.450 132.800 44.180 ;
        RECT 130.840 43.440 131.240 43.450 ;
        RECT 128.780 42.980 130.140 43.440 ;
        RECT 130.420 43.380 130.650 43.440 ;
        RECT 130.860 43.380 131.090 43.440 ;
        RECT 128.780 42.710 131.240 42.980 ;
        RECT 128.780 42.670 130.950 42.710 ;
        RECT 128.780 40.920 130.130 42.670 ;
        RECT 131.410 42.490 132.790 43.450 ;
        RECT 131.410 42.360 132.810 42.490 ;
        RECT 130.690 41.360 132.810 42.360 ;
        RECT 131.410 41.330 132.810 41.360 ;
        RECT 132.530 41.320 132.810 41.330 ;
        RECT 132.970 41.330 133.740 44.270 ;
        RECT 135.520 44.790 136.730 45.450 ;
        RECT 137.880 45.560 138.200 47.775 ;
        RECT 138.880 47.570 139.780 48.380 ;
        RECT 140.350 47.840 140.870 55.730 ;
        RECT 140.350 47.775 140.580 47.840 ;
        RECT 141.350 47.830 141.730 55.750 ;
        RECT 142.430 49.350 143.250 55.980 ;
        RECT 143.780 55.730 144.010 55.775 ;
        RECT 144.920 55.730 145.150 55.775 ;
        RECT 142.340 48.350 143.340 49.350 ;
        RECT 141.360 47.775 141.720 47.830 ;
        RECT 138.340 47.340 140.300 47.570 ;
        RECT 141.360 46.210 141.620 47.775 ;
        RECT 142.430 47.570 143.250 48.350 ;
        RECT 143.780 47.860 145.160 55.730 ;
        RECT 145.490 55.610 145.930 55.980 ;
        RECT 146.210 55.730 146.440 55.775 ;
        RECT 146.840 55.730 147.980 56.540 ;
        RECT 145.490 48.240 145.920 55.610 ;
        RECT 146.210 51.750 147.980 55.730 ;
        RECT 146.210 50.750 147.970 51.750 ;
        RECT 143.780 47.775 144.010 47.860 ;
        RECT 144.920 47.775 145.150 47.860 ;
        RECT 145.490 47.570 145.930 48.240 ;
        RECT 146.210 47.870 147.980 50.750 ;
        RECT 146.210 47.775 146.440 47.870 ;
        RECT 141.770 47.340 143.730 47.570 ;
        RECT 145.200 47.340 146.160 47.570 ;
        RECT 145.300 46.460 146.090 47.340 ;
        RECT 146.840 46.860 147.980 47.870 ;
        RECT 141.360 45.590 144.980 46.210 ;
        RECT 145.250 45.700 146.140 46.460 ;
        RECT 135.520 44.560 136.880 44.790 ;
        RECT 135.520 43.390 136.610 44.560 ;
        RECT 137.880 44.400 138.210 45.560 ;
        RECT 138.350 44.560 140.310 44.790 ;
        RECT 132.530 41.270 132.760 41.320 ;
        RECT 132.970 41.270 133.200 41.330 ;
        RECT 128.780 40.600 131.480 40.920 ;
        RECT 128.780 40.370 129.010 40.600 ;
        RECT 125.690 39.750 126.050 40.050 ;
        RECT 126.770 39.980 128.730 40.210 ;
        RECT 129.390 39.750 131.480 40.600 ;
        RECT 135.530 40.440 136.610 43.390 ;
        RECT 135.580 40.240 136.610 40.440 ;
        RECT 136.930 44.390 137.160 44.400 ;
        RECT 136.930 42.080 137.340 44.390 ;
        RECT 137.880 44.380 138.300 44.400 ;
        RECT 137.880 44.330 138.390 44.380 ;
        RECT 138.740 44.330 140.000 44.560 ;
        RECT 141.360 44.400 141.620 45.590 ;
        RECT 144.570 44.940 144.970 45.590 ;
        RECT 146.910 45.540 147.980 46.860 ;
        RECT 146.910 45.040 148.750 45.540 ;
        RECT 145.970 44.940 146.720 44.950 ;
        RECT 144.570 44.890 146.720 44.940 ;
        RECT 144.570 44.850 146.900 44.890 ;
        RECT 141.780 44.560 143.740 44.790 ;
        RECT 144.570 44.600 148.130 44.850 ;
        RECT 144.570 44.590 145.910 44.600 ;
        RECT 145.620 44.570 145.910 44.590 ;
        RECT 136.930 40.400 137.430 42.080 ;
        RECT 137.880 40.470 140.000 44.330 ;
        RECT 138.000 40.460 140.000 40.470 ;
        RECT 138.070 40.400 138.300 40.460 ;
        RECT 135.580 40.060 136.880 40.240 ;
        RECT 135.920 40.010 136.880 40.060 ;
        RECT 137.230 39.780 137.430 40.400 ;
        RECT 138.660 40.240 140.000 40.460 ;
        RECT 140.360 44.360 140.590 44.400 ;
        RECT 141.360 44.370 141.730 44.400 ;
        RECT 141.360 44.360 141.810 44.370 ;
        RECT 140.360 44.350 140.770 44.360 ;
        RECT 140.360 42.130 140.810 44.350 ;
        RECT 140.360 41.640 140.860 42.130 ;
        RECT 140.360 40.970 140.950 41.640 ;
        RECT 140.360 40.720 141.010 40.970 ;
        RECT 140.360 40.690 141.060 40.720 ;
        RECT 140.360 40.400 140.590 40.690 ;
        RECT 140.820 40.320 141.060 40.690 ;
        RECT 141.310 40.460 141.810 44.360 ;
        RECT 141.310 40.450 141.730 40.460 ;
        RECT 141.370 40.440 141.730 40.450 ;
        RECT 141.500 40.400 141.730 40.440 ;
        RECT 138.350 40.010 140.310 40.240 ;
        RECT 140.740 40.080 141.060 40.320 ;
        RECT 142.070 40.240 143.440 44.560 ;
        RECT 146.780 44.510 148.130 44.600 ;
        RECT 147.730 44.505 148.020 44.510 ;
        RECT 143.790 44.220 144.020 44.400 ;
        RECT 145.430 44.350 145.660 44.410 ;
        RECT 145.870 44.350 146.100 44.410 ;
        RECT 144.680 44.340 145.660 44.350 ;
        RECT 144.250 44.220 145.660 44.340 ;
        RECT 143.790 43.470 145.660 44.220 ;
        RECT 145.850 44.210 146.250 44.350 ;
        RECT 148.380 44.300 148.750 45.040 ;
        RECT 147.540 44.210 147.770 44.300 ;
        RECT 145.850 43.480 147.810 44.210 ;
        RECT 145.850 43.470 146.250 43.480 ;
        RECT 143.790 43.010 145.150 43.470 ;
        RECT 145.430 43.410 145.660 43.470 ;
        RECT 145.870 43.410 146.100 43.470 ;
        RECT 143.790 42.740 146.250 43.010 ;
        RECT 143.790 42.700 145.960 42.740 ;
        RECT 143.790 40.950 145.140 42.700 ;
        RECT 146.420 42.520 147.800 43.480 ;
        RECT 146.420 42.390 147.820 42.520 ;
        RECT 145.700 41.390 147.820 42.390 ;
        RECT 146.420 41.360 147.820 41.390 ;
        RECT 147.540 41.350 147.820 41.360 ;
        RECT 147.980 41.360 148.750 44.300 ;
        RECT 147.540 41.300 147.770 41.350 ;
        RECT 147.980 41.300 148.210 41.360 ;
        RECT 143.790 40.630 146.490 40.950 ;
        RECT 143.790 40.400 144.020 40.630 ;
        RECT 140.700 39.780 141.060 40.080 ;
        RECT 141.780 40.010 143.740 40.240 ;
        RECT 144.400 39.780 146.490 40.630 ;
        RECT 90.100 39.730 101.460 39.750 ;
        RECT 105.140 39.730 116.500 39.750 ;
        RECT 90.100 39.710 116.500 39.730 ;
        RECT 72.240 38.240 73.080 39.600 ;
        RECT 73.770 39.400 74.020 39.710 ;
        RECT 74.550 39.690 116.500 39.710 ;
        RECT 120.120 39.690 131.480 39.750 ;
        RECT 74.550 39.680 131.480 39.690 ;
        RECT 135.130 39.680 146.490 39.780 ;
        RECT 72.240 37.690 72.870 38.240 ;
        RECT 73.360 37.870 74.070 39.400 ;
        RECT 74.550 39.030 146.490 39.680 ;
        RECT 74.550 39.000 146.480 39.030 ;
        RECT 74.550 38.980 101.450 39.000 ;
        RECT 74.550 38.930 86.470 38.980 ;
        RECT 74.550 38.900 75.260 38.930 ;
        RECT 90.070 38.920 101.450 38.980 ;
        RECT 105.110 38.960 146.480 39.000 ;
        RECT 105.110 38.920 116.490 38.960 ;
        RECT 120.090 38.950 146.480 38.960 ;
        RECT 120.090 38.920 131.470 38.950 ;
        RECT 117.460 38.470 120.590 38.490 ;
        RECT 72.290 37.605 72.540 37.690 ;
        RECT 73.130 37.650 74.070 37.870 ;
        RECT 75.130 38.440 87.980 38.470 ;
        RECT 90.070 38.440 102.920 38.470 ;
        RECT 75.130 38.430 102.920 38.440 ;
        RECT 105.080 38.430 132.970 38.470 ;
        RECT 135.080 38.430 147.930 38.470 ;
        RECT 75.130 38.340 147.930 38.430 ;
        RECT 67.945 37.105 69.195 37.475 ;
        RECT 73.130 37.200 73.430 37.650 ;
        RECT 73.770 37.605 74.020 37.650 ;
        RECT 75.130 37.540 147.960 38.340 ;
        RECT 75.130 37.510 117.960 37.540 ;
        RECT 120.120 37.510 147.960 37.540 ;
        RECT 66.540 36.010 67.600 36.280 ;
        RECT 65.600 35.910 66.350 35.920 ;
        RECT 64.200 35.860 66.350 35.910 ;
        RECT 64.200 35.820 66.530 35.860 ;
        RECT 61.410 35.530 63.370 35.760 ;
        RECT 64.200 35.570 67.760 35.820 ;
        RECT 64.200 35.560 65.540 35.570 ;
        RECT 65.250 35.540 65.540 35.560 ;
        RECT 57.510 34.400 59.630 35.330 ;
        RECT 56.560 31.370 57.060 33.050 ;
        RECT 57.630 31.430 59.630 34.400 ;
        RECT 57.700 31.370 57.930 31.430 ;
        RECT 55.550 30.980 56.510 31.210 ;
        RECT 56.860 30.750 57.060 31.370 ;
        RECT 58.290 31.210 59.630 31.430 ;
        RECT 59.990 35.320 60.220 35.370 ;
        RECT 60.990 35.320 61.360 35.370 ;
        RECT 61.700 35.320 63.070 35.530 ;
        RECT 66.410 35.480 67.760 35.570 ;
        RECT 67.360 35.475 67.650 35.480 ;
        RECT 59.990 33.100 60.440 35.320 ;
        RECT 60.990 35.030 63.070 35.320 ;
        RECT 59.990 32.610 60.490 33.100 ;
        RECT 59.990 31.940 60.580 32.610 ;
        RECT 59.990 31.690 60.640 31.940 ;
        RECT 59.990 31.660 60.690 31.690 ;
        RECT 59.990 31.370 60.220 31.660 ;
        RECT 60.450 31.290 60.690 31.660 ;
        RECT 61.000 31.430 63.070 35.030 ;
        RECT 61.000 31.410 61.360 31.430 ;
        RECT 61.130 31.370 61.360 31.410 ;
        RECT 57.980 30.980 59.940 31.210 ;
        RECT 60.370 31.050 60.690 31.290 ;
        RECT 61.700 31.210 63.070 31.430 ;
        RECT 63.420 35.190 63.650 35.370 ;
        RECT 65.060 35.320 65.290 35.380 ;
        RECT 65.500 35.320 65.730 35.380 ;
        RECT 64.310 35.310 65.290 35.320 ;
        RECT 63.880 35.190 65.290 35.310 ;
        RECT 63.420 34.440 65.290 35.190 ;
        RECT 65.480 35.180 65.880 35.320 ;
        RECT 67.170 35.180 67.400 35.270 ;
        RECT 65.480 34.450 67.440 35.180 ;
        RECT 65.480 34.440 65.880 34.450 ;
        RECT 63.420 33.980 64.780 34.440 ;
        RECT 65.060 34.380 65.290 34.440 ;
        RECT 65.500 34.380 65.730 34.440 ;
        RECT 63.420 33.710 65.880 33.980 ;
        RECT 63.420 33.670 65.590 33.710 ;
        RECT 63.420 31.920 64.770 33.670 ;
        RECT 66.050 33.490 67.430 34.450 ;
        RECT 66.050 33.360 67.450 33.490 ;
        RECT 65.330 32.360 67.450 33.360 ;
        RECT 66.050 32.330 67.450 32.360 ;
        RECT 67.170 32.320 67.450 32.330 ;
        RECT 67.170 32.270 67.400 32.320 ;
        RECT 67.610 32.270 67.840 35.270 ;
        RECT 63.420 31.620 66.120 31.920 ;
        RECT 63.420 31.370 63.650 31.620 ;
        RECT 60.330 30.750 60.690 31.050 ;
        RECT 61.410 30.980 63.370 31.210 ;
        RECT 64.030 30.750 66.120 31.620 ;
        RECT 54.760 30.180 66.120 30.750 ;
        RECT 54.730 30.000 66.120 30.180 ;
        RECT 54.730 29.920 66.110 30.000 ;
        RECT 54.055 29.505 61.125 29.655 ;
        RECT 53.625 29.065 60.725 29.275 ;
        RECT 53.035 28.675 60.235 28.890 ;
        RECT 60.020 17.620 60.235 28.675 ;
        RECT 60.515 18.085 60.725 29.065 ;
        RECT 60.975 22.235 61.125 29.505 ;
        RECT 61.490 28.980 66.810 29.180 ;
        RECT 61.440 28.570 66.810 28.980 ;
        RECT 61.440 28.490 63.410 28.570 ;
        RECT 61.440 28.210 63.240 28.490 ;
        RECT 61.490 28.160 63.240 28.210 ;
        RECT 61.490 27.370 61.840 28.160 ;
        RECT 63.990 28.140 66.790 28.390 ;
        RECT 62.230 27.920 62.520 27.950 ;
        RECT 62.220 27.670 62.540 27.920 ;
        RECT 63.990 27.515 64.150 28.140 ;
        RECT 64.290 27.670 64.620 28.000 ;
        RECT 64.900 27.870 65.110 28.140 ;
        RECT 64.970 27.530 65.110 27.870 ;
        RECT 65.250 27.670 65.580 28.000 ;
        RECT 66.050 27.660 66.790 28.140 ;
        RECT 64.970 27.515 65.260 27.530 ;
        RECT 66.050 27.515 66.220 27.660 ;
        RECT 66.400 27.580 66.790 27.660 ;
        RECT 62.040 27.370 62.270 27.515 ;
        RECT 61.490 23.515 62.270 27.370 ;
        RECT 62.480 27.460 62.710 27.515 ;
        RECT 62.480 24.280 63.120 27.460 ;
        RECT 62.480 23.570 63.130 24.280 ;
        RECT 63.620 23.750 63.850 27.515 ;
        RECT 63.990 27.370 64.330 27.515 ;
        RECT 62.480 23.515 62.710 23.570 ;
        RECT 61.490 23.500 62.240 23.515 ;
        RECT 61.490 23.490 61.840 23.500 ;
        RECT 62.230 23.210 62.520 23.310 ;
        RECT 61.990 22.700 62.670 23.210 ;
        RECT 61.490 22.235 62.670 22.700 ;
        RECT 60.975 22.085 62.670 22.235 ;
        RECT 61.490 21.700 62.670 22.085 ;
        RECT 61.990 21.210 62.670 21.700 ;
        RECT 62.220 21.170 62.510 21.210 ;
        RECT 62.030 20.960 62.260 21.010 ;
        RECT 61.490 20.080 62.260 20.960 ;
        RECT 61.490 19.860 61.890 20.080 ;
        RECT 62.030 20.010 62.260 20.080 ;
        RECT 62.470 20.950 62.700 21.010 ;
        RECT 62.910 20.950 63.130 23.570 ;
        RECT 63.410 23.515 63.850 23.750 ;
        RECT 64.100 23.515 64.330 27.370 ;
        RECT 64.580 23.690 64.810 27.515 ;
        RECT 64.970 27.380 65.290 27.515 ;
        RECT 64.470 23.515 64.810 23.690 ;
        RECT 65.060 23.515 65.290 27.380 ;
        RECT 65.540 23.710 65.770 27.515 ;
        RECT 65.460 23.660 65.770 23.710 ;
        RECT 65.430 23.515 65.770 23.660 ;
        RECT 66.020 23.515 66.250 27.515 ;
        RECT 63.410 23.500 63.700 23.515 ;
        RECT 64.470 23.510 64.680 23.515 ;
        RECT 65.430 23.510 65.630 23.515 ;
        RECT 63.410 22.820 63.670 23.500 ;
        RECT 63.810 23.030 64.140 23.360 ;
        RECT 64.470 22.850 64.630 23.510 ;
        RECT 64.770 23.030 65.100 23.360 ;
        RECT 65.430 22.880 65.590 23.510 ;
        RECT 65.730 23.030 66.060 23.360 ;
        RECT 63.410 22.810 63.700 22.820 ;
        RECT 64.470 22.810 64.680 22.850 ;
        RECT 65.430 22.810 65.630 22.880 ;
        RECT 63.410 22.670 65.630 22.810 ;
        RECT 66.490 22.760 66.780 27.580 ;
        RECT 62.470 20.670 63.130 20.950 ;
        RECT 63.400 22.640 65.630 22.670 ;
        RECT 63.400 22.160 65.600 22.640 ;
        RECT 66.020 22.475 67.020 22.760 ;
        RECT 68.825 22.475 69.195 37.105 ;
        RECT 72.290 36.990 72.540 37.015 ;
        RECT 72.910 37.000 73.430 37.200 ;
        RECT 75.940 37.150 76.900 37.180 ;
        RECT 73.770 37.010 74.020 37.015 ;
        RECT 72.910 36.990 73.260 37.000 ;
        RECT 72.260 36.530 73.260 36.990 ;
        RECT 72.260 34.890 73.080 36.530 ;
        RECT 73.720 36.290 74.070 37.010 ;
        RECT 75.610 36.950 76.900 37.150 ;
        RECT 75.610 36.710 76.670 36.950 ;
        RECT 77.170 36.745 77.390 37.510 ;
        RECT 86.870 37.490 90.420 37.510 ;
        RECT 78.370 36.950 80.330 37.180 ;
        RECT 81.800 36.950 83.760 37.180 ;
        RECT 85.230 36.950 86.190 37.180 ;
        RECT 73.340 34.900 74.070 36.290 ;
        RECT 73.340 34.590 74.050 34.900 ;
        RECT 72.630 34.440 74.050 34.590 ;
        RECT 72.630 34.390 73.610 34.440 ;
        RECT 72.250 34.120 73.610 34.390 ;
        RECT 72.250 31.590 72.760 34.120 ;
        RECT 73.250 31.900 74.060 33.740 ;
        RECT 73.000 31.590 74.060 31.900 ;
        RECT 73.000 31.210 73.310 31.590 ;
        RECT 72.770 31.030 73.310 31.210 ;
        RECT 72.250 30.930 73.310 31.030 ;
        RECT 72.250 30.690 73.110 30.930 ;
        RECT 72.250 28.900 72.910 30.690 ;
        RECT 73.720 29.770 74.090 31.040 ;
        RECT 73.390 29.730 74.090 29.770 ;
        RECT 73.320 28.870 74.090 29.730 ;
        RECT 75.560 29.600 76.670 36.710 ;
        RECT 73.320 28.600 73.900 28.870 ;
        RECT 70.760 28.420 73.900 28.600 ;
        RECT 70.740 28.350 73.900 28.420 ;
        RECT 75.550 28.540 76.670 29.600 ;
        RECT 76.950 36.540 77.390 36.745 ;
        RECT 78.090 36.720 78.320 36.745 ;
        RECT 78.090 36.710 78.330 36.720 ;
        RECT 76.950 28.800 77.340 36.540 ;
        RECT 77.920 29.650 78.330 36.710 ;
        RECT 78.910 30.360 79.810 36.950 ;
        RECT 80.380 36.700 80.610 36.745 ;
        RECT 81.520 36.720 81.750 36.745 ;
        RECT 77.910 28.830 78.330 29.650 ;
        RECT 78.880 29.350 79.880 30.360 ;
        RECT 76.950 28.745 77.180 28.800 ;
        RECT 77.910 28.745 78.320 28.830 ;
        RECT 70.740 28.190 73.890 28.350 ;
        RECT 75.550 28.310 76.900 28.540 ;
        RECT 70.740 25.610 71.130 28.190 ;
        RECT 72.240 27.760 72.660 27.770 ;
        RECT 71.710 27.750 72.660 27.760 ;
        RECT 71.420 25.610 72.660 27.750 ;
        RECT 73.260 25.850 74.090 27.770 ;
        RECT 75.550 27.670 76.760 28.310 ;
        RECT 75.110 26.420 76.760 27.670 ;
        RECT 73.150 25.610 74.090 25.850 ;
        RECT 71.420 25.590 72.580 25.610 ;
        RECT 71.420 25.050 71.880 25.590 ;
        RECT 73.150 25.170 73.380 25.610 ;
        RECT 72.750 25.070 73.380 25.170 ;
        RECT 70.770 24.850 71.880 25.050 ;
        RECT 72.260 24.870 73.380 25.070 ;
        RECT 73.710 25.040 74.120 25.050 ;
        RECT 74.550 25.040 75.280 26.250 ;
        RECT 70.770 22.930 71.810 24.850 ;
        RECT 72.260 24.710 73.230 24.870 ;
        RECT 72.260 22.920 72.890 24.710 ;
        RECT 73.710 22.900 75.280 25.040 ;
        RECT 75.550 25.760 76.760 26.420 ;
        RECT 77.910 26.530 78.230 28.745 ;
        RECT 78.910 28.540 79.810 29.350 ;
        RECT 80.380 28.810 80.900 36.700 ;
        RECT 80.380 28.745 80.610 28.810 ;
        RECT 81.380 28.800 81.760 36.720 ;
        RECT 82.460 30.320 83.280 36.950 ;
        RECT 83.810 36.700 84.040 36.745 ;
        RECT 84.950 36.700 85.180 36.745 ;
        RECT 82.370 29.320 83.370 30.320 ;
        RECT 81.390 28.745 81.750 28.800 ;
        RECT 78.370 28.310 80.330 28.540 ;
        RECT 81.390 27.180 81.650 28.745 ;
        RECT 82.460 28.540 83.280 29.320 ;
        RECT 83.810 28.830 85.190 36.700 ;
        RECT 85.520 36.580 85.960 36.950 ;
        RECT 86.240 36.700 86.470 36.745 ;
        RECT 86.870 36.700 88.010 37.490 ;
        RECT 88.340 36.880 89.740 37.490 ;
        RECT 90.880 37.150 91.840 37.180 ;
        RECT 90.550 36.950 91.840 37.150 ;
        RECT 90.550 36.710 91.610 36.950 ;
        RECT 92.110 36.745 92.330 37.510 ;
        RECT 101.810 37.480 105.800 37.510 ;
        RECT 93.310 36.950 95.270 37.180 ;
        RECT 96.740 36.950 98.700 37.180 ;
        RECT 100.170 36.950 101.130 37.180 ;
        RECT 85.520 29.210 85.950 36.580 ;
        RECT 86.240 32.720 88.010 36.700 ;
        RECT 86.240 31.720 88.000 32.720 ;
        RECT 83.810 28.745 84.040 28.830 ;
        RECT 84.950 28.745 85.180 28.830 ;
        RECT 85.520 28.540 85.960 29.210 ;
        RECT 86.240 28.840 88.010 31.720 ;
        RECT 90.500 29.600 91.610 36.710 ;
        RECT 86.240 28.745 86.470 28.840 ;
        RECT 81.800 28.310 83.760 28.540 ;
        RECT 85.230 28.310 86.190 28.540 ;
        RECT 85.330 27.430 86.120 28.310 ;
        RECT 86.870 27.830 88.010 28.840 ;
        RECT 81.390 26.560 85.010 27.180 ;
        RECT 85.280 26.670 86.170 27.430 ;
        RECT 75.550 25.530 76.910 25.760 ;
        RECT 75.550 24.360 76.640 25.530 ;
        RECT 77.910 25.370 78.240 26.530 ;
        RECT 78.380 25.530 80.340 25.760 ;
        RECT 73.710 22.890 74.120 22.900 ;
        RECT 74.570 22.730 75.280 22.900 ;
        RECT 63.400 21.810 65.870 22.160 ;
        RECT 66.020 22.105 69.195 22.475 ;
        RECT 74.550 22.260 75.300 22.730 ;
        RECT 63.400 21.720 65.880 21.810 ;
        RECT 66.020 21.760 67.020 22.105 ;
        RECT 63.400 21.010 63.810 21.720 ;
        RECT 64.280 21.170 64.610 21.500 ;
        RECT 64.760 21.150 64.930 21.720 ;
        RECT 65.550 21.710 65.880 21.720 ;
        RECT 65.240 21.170 65.570 21.500 ;
        RECT 65.730 21.150 65.880 21.710 ;
        RECT 64.760 21.010 64.900 21.150 ;
        RECT 65.730 21.010 65.870 21.150 ;
        RECT 63.400 20.770 63.840 21.010 ;
        RECT 62.470 20.070 63.100 20.670 ;
        RECT 62.470 20.010 62.700 20.070 ;
        RECT 63.610 20.010 63.840 20.770 ;
        RECT 64.090 20.180 64.320 21.010 ;
        RECT 64.570 20.780 64.900 21.010 ;
        RECT 64.090 20.010 64.420 20.180 ;
        RECT 64.570 20.010 64.800 20.780 ;
        RECT 65.050 20.240 65.280 21.010 ;
        RECT 65.530 20.790 65.870 21.010 ;
        RECT 66.010 20.930 66.240 21.010 ;
        RECT 66.490 20.930 66.780 21.760 ;
        RECT 65.050 20.010 65.390 20.240 ;
        RECT 65.530 20.010 65.760 20.790 ;
        RECT 66.010 20.010 66.780 20.930 ;
        RECT 61.490 19.320 61.980 19.860 ;
        RECT 62.190 19.640 62.540 19.850 ;
        RECT 62.200 19.580 62.540 19.640 ;
        RECT 63.800 19.530 64.130 19.860 ;
        RECT 64.280 19.370 64.420 20.010 ;
        RECT 65.230 19.860 65.390 20.010 ;
        RECT 64.760 19.530 65.090 19.860 ;
        RECT 65.230 19.370 65.400 19.860 ;
        RECT 65.720 19.530 66.050 19.860 ;
        RECT 66.190 19.370 66.780 20.010 ;
        RECT 74.560 20.750 75.300 22.260 ;
        RECT 75.560 21.410 76.640 24.360 ;
        RECT 75.610 21.210 76.640 21.410 ;
        RECT 76.960 25.360 77.190 25.370 ;
        RECT 76.960 23.050 77.370 25.360 ;
        RECT 77.910 25.350 78.330 25.370 ;
        RECT 77.910 25.300 78.420 25.350 ;
        RECT 78.770 25.300 80.030 25.530 ;
        RECT 81.390 25.370 81.650 26.560 ;
        RECT 84.600 25.910 85.000 26.560 ;
        RECT 86.940 26.510 88.010 27.830 ;
        RECT 90.490 28.540 91.610 29.600 ;
        RECT 91.890 36.540 92.330 36.745 ;
        RECT 93.030 36.720 93.260 36.745 ;
        RECT 93.030 36.710 93.270 36.720 ;
        RECT 91.890 28.800 92.280 36.540 ;
        RECT 92.860 29.650 93.270 36.710 ;
        RECT 93.850 30.360 94.750 36.950 ;
        RECT 95.320 36.700 95.550 36.745 ;
        RECT 96.460 36.720 96.690 36.745 ;
        RECT 92.850 28.830 93.270 29.650 ;
        RECT 93.820 29.350 94.820 30.360 ;
        RECT 91.890 28.745 92.120 28.800 ;
        RECT 92.850 28.745 93.260 28.830 ;
        RECT 90.490 28.310 91.840 28.540 ;
        RECT 90.490 27.670 91.700 28.310 ;
        RECT 86.940 26.010 88.780 26.510 ;
        RECT 90.050 26.420 91.700 27.670 ;
        RECT 86.000 25.910 86.750 25.920 ;
        RECT 84.600 25.860 86.750 25.910 ;
        RECT 84.600 25.820 86.930 25.860 ;
        RECT 81.810 25.530 83.770 25.760 ;
        RECT 84.600 25.570 88.160 25.820 ;
        RECT 84.600 25.560 85.940 25.570 ;
        RECT 85.650 25.540 85.940 25.560 ;
        RECT 76.960 21.370 77.460 23.050 ;
        RECT 77.910 21.440 80.030 25.300 ;
        RECT 78.030 21.430 80.030 21.440 ;
        RECT 78.100 21.370 78.330 21.430 ;
        RECT 75.610 21.030 76.910 21.210 ;
        RECT 75.950 20.980 76.910 21.030 ;
        RECT 77.260 20.750 77.460 21.370 ;
        RECT 78.690 21.210 80.030 21.430 ;
        RECT 80.390 25.330 80.620 25.370 ;
        RECT 81.390 25.340 81.760 25.370 ;
        RECT 81.390 25.330 81.840 25.340 ;
        RECT 80.390 25.320 80.800 25.330 ;
        RECT 80.390 23.100 80.840 25.320 ;
        RECT 80.390 22.610 80.890 23.100 ;
        RECT 80.390 21.940 80.980 22.610 ;
        RECT 80.390 21.690 81.040 21.940 ;
        RECT 80.390 21.660 81.090 21.690 ;
        RECT 80.390 21.370 80.620 21.660 ;
        RECT 80.850 21.290 81.090 21.660 ;
        RECT 81.340 21.430 81.840 25.330 ;
        RECT 81.340 21.420 81.760 21.430 ;
        RECT 81.400 21.410 81.760 21.420 ;
        RECT 81.530 21.370 81.760 21.410 ;
        RECT 78.380 20.980 80.340 21.210 ;
        RECT 80.770 21.050 81.090 21.290 ;
        RECT 82.100 21.210 83.470 25.530 ;
        RECT 86.810 25.480 88.160 25.570 ;
        RECT 87.760 25.475 88.050 25.480 ;
        RECT 83.820 25.190 84.050 25.370 ;
        RECT 85.460 25.320 85.690 25.380 ;
        RECT 85.900 25.320 86.130 25.380 ;
        RECT 84.710 25.310 85.690 25.320 ;
        RECT 84.280 25.190 85.690 25.310 ;
        RECT 83.820 24.440 85.690 25.190 ;
        RECT 85.880 25.180 86.280 25.320 ;
        RECT 88.410 25.270 88.780 26.010 ;
        RECT 87.570 25.180 87.800 25.270 ;
        RECT 85.880 24.450 87.840 25.180 ;
        RECT 85.880 24.440 86.280 24.450 ;
        RECT 83.820 23.980 85.180 24.440 ;
        RECT 85.460 24.380 85.690 24.440 ;
        RECT 85.900 24.380 86.130 24.440 ;
        RECT 83.820 23.710 86.280 23.980 ;
        RECT 83.820 23.670 85.990 23.710 ;
        RECT 83.820 21.920 85.170 23.670 ;
        RECT 86.450 23.490 87.830 24.450 ;
        RECT 86.450 23.360 87.850 23.490 ;
        RECT 85.730 22.360 87.850 23.360 ;
        RECT 86.450 22.330 87.850 22.360 ;
        RECT 87.570 22.320 87.850 22.330 ;
        RECT 88.010 22.330 88.780 25.270 ;
        RECT 90.490 25.760 91.700 26.420 ;
        RECT 92.850 26.530 93.170 28.745 ;
        RECT 93.850 28.540 94.750 29.350 ;
        RECT 95.320 28.810 95.840 36.700 ;
        RECT 95.320 28.745 95.550 28.810 ;
        RECT 96.320 28.800 96.700 36.720 ;
        RECT 97.400 30.320 98.220 36.950 ;
        RECT 98.750 36.700 98.980 36.745 ;
        RECT 99.890 36.700 100.120 36.745 ;
        RECT 97.310 29.320 98.310 30.320 ;
        RECT 96.330 28.745 96.690 28.800 ;
        RECT 93.310 28.310 95.270 28.540 ;
        RECT 96.330 27.180 96.590 28.745 ;
        RECT 97.400 28.540 98.220 29.320 ;
        RECT 98.750 28.830 100.130 36.700 ;
        RECT 100.460 36.580 100.900 36.950 ;
        RECT 101.180 36.700 101.410 36.745 ;
        RECT 101.810 36.700 102.950 37.480 ;
        RECT 105.890 37.150 106.850 37.180 ;
        RECT 105.560 36.950 106.850 37.150 ;
        RECT 105.560 36.710 106.620 36.950 ;
        RECT 107.120 36.745 107.340 37.510 ;
        RECT 108.320 36.950 110.280 37.180 ;
        RECT 111.750 36.950 113.710 37.180 ;
        RECT 115.180 36.950 116.140 37.180 ;
        RECT 100.460 29.210 100.890 36.580 ;
        RECT 101.180 32.720 102.950 36.700 ;
        RECT 101.180 31.720 102.940 32.720 ;
        RECT 98.750 28.745 98.980 28.830 ;
        RECT 99.890 28.745 100.120 28.830 ;
        RECT 100.460 28.540 100.900 29.210 ;
        RECT 101.180 28.840 102.950 31.720 ;
        RECT 105.510 29.600 106.620 36.710 ;
        RECT 101.180 28.745 101.410 28.840 ;
        RECT 96.740 28.310 98.700 28.540 ;
        RECT 100.170 28.310 101.130 28.540 ;
        RECT 100.270 27.430 101.060 28.310 ;
        RECT 101.810 27.830 102.950 28.840 ;
        RECT 96.330 26.560 99.950 27.180 ;
        RECT 100.220 26.670 101.110 27.430 ;
        RECT 90.490 25.530 91.850 25.760 ;
        RECT 90.490 24.360 91.580 25.530 ;
        RECT 92.850 25.370 93.180 26.530 ;
        RECT 93.320 25.530 95.280 25.760 ;
        RECT 87.570 22.270 87.800 22.320 ;
        RECT 88.010 22.270 88.240 22.330 ;
        RECT 83.820 21.600 86.520 21.920 ;
        RECT 83.820 21.370 84.050 21.600 ;
        RECT 80.730 20.750 81.090 21.050 ;
        RECT 81.810 20.980 83.770 21.210 ;
        RECT 84.430 20.750 86.520 21.600 ;
        RECT 90.500 21.410 91.580 24.360 ;
        RECT 90.550 21.210 91.580 21.410 ;
        RECT 91.900 25.360 92.130 25.370 ;
        RECT 91.900 23.050 92.310 25.360 ;
        RECT 92.850 25.350 93.270 25.370 ;
        RECT 92.850 25.300 93.360 25.350 ;
        RECT 93.710 25.300 94.970 25.530 ;
        RECT 96.330 25.370 96.590 26.560 ;
        RECT 99.540 25.910 99.940 26.560 ;
        RECT 101.880 26.510 102.950 27.830 ;
        RECT 105.500 28.540 106.620 29.600 ;
        RECT 106.900 36.540 107.340 36.745 ;
        RECT 108.040 36.720 108.270 36.745 ;
        RECT 108.040 36.710 108.280 36.720 ;
        RECT 106.900 28.800 107.290 36.540 ;
        RECT 107.870 29.650 108.280 36.710 ;
        RECT 108.860 30.360 109.760 36.950 ;
        RECT 110.330 36.700 110.560 36.745 ;
        RECT 111.470 36.720 111.700 36.745 ;
        RECT 107.860 28.830 108.280 29.650 ;
        RECT 108.830 29.350 109.830 30.360 ;
        RECT 106.900 28.745 107.130 28.800 ;
        RECT 107.860 28.745 108.270 28.830 ;
        RECT 105.500 28.310 106.850 28.540 ;
        RECT 105.500 27.670 106.710 28.310 ;
        RECT 101.880 26.010 103.720 26.510 ;
        RECT 105.060 26.420 106.710 27.670 ;
        RECT 100.940 25.910 101.690 25.920 ;
        RECT 99.540 25.860 101.690 25.910 ;
        RECT 99.540 25.820 101.870 25.860 ;
        RECT 96.750 25.530 98.710 25.760 ;
        RECT 99.540 25.570 103.100 25.820 ;
        RECT 99.540 25.560 100.880 25.570 ;
        RECT 100.590 25.540 100.880 25.560 ;
        RECT 91.900 21.370 92.400 23.050 ;
        RECT 92.850 21.440 94.970 25.300 ;
        RECT 92.970 21.430 94.970 21.440 ;
        RECT 93.040 21.370 93.270 21.430 ;
        RECT 90.550 21.030 91.850 21.210 ;
        RECT 90.890 20.980 91.850 21.030 ;
        RECT 92.200 20.750 92.400 21.370 ;
        RECT 93.630 21.210 94.970 21.430 ;
        RECT 95.330 25.330 95.560 25.370 ;
        RECT 96.330 25.340 96.700 25.370 ;
        RECT 96.330 25.330 96.780 25.340 ;
        RECT 95.330 25.320 95.740 25.330 ;
        RECT 95.330 23.100 95.780 25.320 ;
        RECT 95.330 22.610 95.830 23.100 ;
        RECT 95.330 21.940 95.920 22.610 ;
        RECT 95.330 21.690 95.980 21.940 ;
        RECT 95.330 21.660 96.030 21.690 ;
        RECT 95.330 21.370 95.560 21.660 ;
        RECT 95.790 21.290 96.030 21.660 ;
        RECT 96.280 21.430 96.780 25.330 ;
        RECT 96.280 21.420 96.700 21.430 ;
        RECT 96.340 21.410 96.700 21.420 ;
        RECT 96.470 21.370 96.700 21.410 ;
        RECT 93.320 20.980 95.280 21.210 ;
        RECT 95.710 21.050 96.030 21.290 ;
        RECT 97.040 21.210 98.410 25.530 ;
        RECT 101.750 25.480 103.100 25.570 ;
        RECT 102.700 25.475 102.990 25.480 ;
        RECT 98.760 25.190 98.990 25.370 ;
        RECT 100.400 25.320 100.630 25.380 ;
        RECT 100.840 25.320 101.070 25.380 ;
        RECT 99.650 25.310 100.630 25.320 ;
        RECT 99.220 25.190 100.630 25.310 ;
        RECT 98.760 24.440 100.630 25.190 ;
        RECT 100.820 25.180 101.220 25.320 ;
        RECT 103.350 25.270 103.720 26.010 ;
        RECT 102.510 25.180 102.740 25.270 ;
        RECT 100.820 24.450 102.780 25.180 ;
        RECT 100.820 24.440 101.220 24.450 ;
        RECT 98.760 23.980 100.120 24.440 ;
        RECT 100.400 24.380 100.630 24.440 ;
        RECT 100.840 24.380 101.070 24.440 ;
        RECT 98.760 23.710 101.220 23.980 ;
        RECT 98.760 23.670 100.930 23.710 ;
        RECT 98.760 21.920 100.110 23.670 ;
        RECT 101.390 23.490 102.770 24.450 ;
        RECT 101.390 23.360 102.790 23.490 ;
        RECT 100.670 22.360 102.790 23.360 ;
        RECT 101.390 22.330 102.790 22.360 ;
        RECT 102.510 22.320 102.790 22.330 ;
        RECT 102.950 22.330 103.720 25.270 ;
        RECT 105.500 25.760 106.710 26.420 ;
        RECT 107.860 26.530 108.180 28.745 ;
        RECT 108.860 28.540 109.760 29.350 ;
        RECT 110.330 28.810 110.850 36.700 ;
        RECT 110.330 28.745 110.560 28.810 ;
        RECT 111.330 28.800 111.710 36.720 ;
        RECT 112.410 30.320 113.230 36.950 ;
        RECT 113.760 36.700 113.990 36.745 ;
        RECT 114.900 36.700 115.130 36.745 ;
        RECT 112.320 29.320 113.320 30.320 ;
        RECT 111.340 28.745 111.700 28.800 ;
        RECT 108.320 28.310 110.280 28.540 ;
        RECT 111.340 27.180 111.600 28.745 ;
        RECT 112.410 28.540 113.230 29.320 ;
        RECT 113.760 28.830 115.140 36.700 ;
        RECT 115.470 36.580 115.910 36.950 ;
        RECT 116.190 36.700 116.420 36.745 ;
        RECT 116.820 36.700 117.960 37.510 ;
        RECT 120.930 37.150 121.890 37.180 ;
        RECT 120.600 36.950 121.890 37.150 ;
        RECT 120.600 36.710 121.660 36.950 ;
        RECT 122.160 36.745 122.380 37.510 ;
        RECT 131.860 37.480 135.350 37.510 ;
        RECT 123.360 36.950 125.320 37.180 ;
        RECT 126.790 36.950 128.750 37.180 ;
        RECT 130.220 36.950 131.180 37.180 ;
        RECT 115.470 29.210 115.900 36.580 ;
        RECT 116.190 32.720 117.960 36.700 ;
        RECT 116.190 31.720 117.950 32.720 ;
        RECT 113.760 28.745 113.990 28.830 ;
        RECT 114.900 28.745 115.130 28.830 ;
        RECT 115.470 28.540 115.910 29.210 ;
        RECT 116.190 28.840 117.960 31.720 ;
        RECT 120.550 29.600 121.660 36.710 ;
        RECT 116.190 28.745 116.420 28.840 ;
        RECT 111.750 28.310 113.710 28.540 ;
        RECT 115.180 28.310 116.140 28.540 ;
        RECT 115.280 27.430 116.070 28.310 ;
        RECT 116.820 27.830 117.960 28.840 ;
        RECT 111.340 26.560 114.960 27.180 ;
        RECT 115.230 26.670 116.120 27.430 ;
        RECT 105.500 25.530 106.860 25.760 ;
        RECT 105.500 24.360 106.590 25.530 ;
        RECT 107.860 25.370 108.190 26.530 ;
        RECT 108.330 25.530 110.290 25.760 ;
        RECT 102.510 22.270 102.740 22.320 ;
        RECT 102.950 22.270 103.180 22.330 ;
        RECT 98.760 21.600 101.460 21.920 ;
        RECT 98.760 21.370 98.990 21.600 ;
        RECT 95.670 20.750 96.030 21.050 ;
        RECT 96.750 20.980 98.710 21.210 ;
        RECT 99.370 20.750 101.460 21.600 ;
        RECT 105.510 21.410 106.590 24.360 ;
        RECT 105.560 21.210 106.590 21.410 ;
        RECT 106.910 25.360 107.140 25.370 ;
        RECT 106.910 23.050 107.320 25.360 ;
        RECT 107.860 25.350 108.280 25.370 ;
        RECT 107.860 25.300 108.370 25.350 ;
        RECT 108.720 25.300 109.980 25.530 ;
        RECT 111.340 25.370 111.600 26.560 ;
        RECT 114.550 25.910 114.950 26.560 ;
        RECT 116.890 26.510 117.960 27.830 ;
        RECT 120.540 28.540 121.660 29.600 ;
        RECT 121.940 36.540 122.380 36.745 ;
        RECT 123.080 36.720 123.310 36.745 ;
        RECT 123.080 36.710 123.320 36.720 ;
        RECT 121.940 28.800 122.330 36.540 ;
        RECT 122.910 29.650 123.320 36.710 ;
        RECT 123.900 30.360 124.800 36.950 ;
        RECT 125.370 36.700 125.600 36.745 ;
        RECT 126.510 36.720 126.740 36.745 ;
        RECT 122.900 28.830 123.320 29.650 ;
        RECT 123.870 29.350 124.870 30.360 ;
        RECT 121.940 28.745 122.170 28.800 ;
        RECT 122.900 28.745 123.310 28.830 ;
        RECT 120.540 28.310 121.890 28.540 ;
        RECT 120.540 27.670 121.750 28.310 ;
        RECT 116.890 26.010 118.730 26.510 ;
        RECT 120.100 26.420 121.750 27.670 ;
        RECT 115.950 25.910 116.700 25.920 ;
        RECT 114.550 25.860 116.700 25.910 ;
        RECT 114.550 25.820 116.880 25.860 ;
        RECT 111.760 25.530 113.720 25.760 ;
        RECT 114.550 25.570 118.110 25.820 ;
        RECT 114.550 25.560 115.890 25.570 ;
        RECT 115.600 25.540 115.890 25.560 ;
        RECT 106.910 21.370 107.410 23.050 ;
        RECT 107.860 21.440 109.980 25.300 ;
        RECT 107.980 21.430 109.980 21.440 ;
        RECT 108.050 21.370 108.280 21.430 ;
        RECT 105.560 21.030 106.860 21.210 ;
        RECT 105.900 20.980 106.860 21.030 ;
        RECT 107.210 20.750 107.410 21.370 ;
        RECT 108.640 21.210 109.980 21.430 ;
        RECT 110.340 25.330 110.570 25.370 ;
        RECT 111.340 25.340 111.710 25.370 ;
        RECT 111.340 25.330 111.790 25.340 ;
        RECT 110.340 25.320 110.750 25.330 ;
        RECT 110.340 23.100 110.790 25.320 ;
        RECT 110.340 22.610 110.840 23.100 ;
        RECT 110.340 21.940 110.930 22.610 ;
        RECT 110.340 21.690 110.990 21.940 ;
        RECT 110.340 21.660 111.040 21.690 ;
        RECT 110.340 21.370 110.570 21.660 ;
        RECT 110.800 21.290 111.040 21.660 ;
        RECT 111.290 21.430 111.790 25.330 ;
        RECT 111.290 21.420 111.710 21.430 ;
        RECT 111.350 21.410 111.710 21.420 ;
        RECT 111.480 21.370 111.710 21.410 ;
        RECT 108.330 20.980 110.290 21.210 ;
        RECT 110.720 21.050 111.040 21.290 ;
        RECT 112.050 21.210 113.420 25.530 ;
        RECT 116.760 25.480 118.110 25.570 ;
        RECT 117.710 25.475 118.000 25.480 ;
        RECT 113.770 25.190 114.000 25.370 ;
        RECT 115.410 25.320 115.640 25.380 ;
        RECT 115.850 25.320 116.080 25.380 ;
        RECT 114.660 25.310 115.640 25.320 ;
        RECT 114.230 25.190 115.640 25.310 ;
        RECT 113.770 24.440 115.640 25.190 ;
        RECT 115.830 25.180 116.230 25.320 ;
        RECT 118.360 25.270 118.730 26.010 ;
        RECT 117.520 25.180 117.750 25.270 ;
        RECT 115.830 24.450 117.790 25.180 ;
        RECT 115.830 24.440 116.230 24.450 ;
        RECT 113.770 23.980 115.130 24.440 ;
        RECT 115.410 24.380 115.640 24.440 ;
        RECT 115.850 24.380 116.080 24.440 ;
        RECT 113.770 23.710 116.230 23.980 ;
        RECT 113.770 23.670 115.940 23.710 ;
        RECT 113.770 21.920 115.120 23.670 ;
        RECT 116.400 23.490 117.780 24.450 ;
        RECT 116.400 23.360 117.800 23.490 ;
        RECT 115.680 22.360 117.800 23.360 ;
        RECT 116.400 22.330 117.800 22.360 ;
        RECT 117.520 22.320 117.800 22.330 ;
        RECT 117.960 22.330 118.730 25.270 ;
        RECT 120.540 25.760 121.750 26.420 ;
        RECT 122.900 26.530 123.220 28.745 ;
        RECT 123.900 28.540 124.800 29.350 ;
        RECT 125.370 28.810 125.890 36.700 ;
        RECT 125.370 28.745 125.600 28.810 ;
        RECT 126.370 28.800 126.750 36.720 ;
        RECT 127.450 30.320 128.270 36.950 ;
        RECT 128.800 36.700 129.030 36.745 ;
        RECT 129.940 36.700 130.170 36.745 ;
        RECT 127.360 29.320 128.360 30.320 ;
        RECT 126.380 28.745 126.740 28.800 ;
        RECT 123.360 28.310 125.320 28.540 ;
        RECT 126.380 27.180 126.640 28.745 ;
        RECT 127.450 28.540 128.270 29.320 ;
        RECT 128.800 28.830 130.180 36.700 ;
        RECT 130.510 36.580 130.950 36.950 ;
        RECT 131.230 36.700 131.460 36.745 ;
        RECT 131.860 36.700 133.000 37.480 ;
        RECT 135.890 37.150 136.850 37.180 ;
        RECT 135.560 36.950 136.850 37.150 ;
        RECT 135.560 36.710 136.620 36.950 ;
        RECT 137.120 36.745 137.340 37.510 ;
        RECT 138.320 36.950 140.280 37.180 ;
        RECT 141.750 36.950 143.710 37.180 ;
        RECT 145.180 36.950 146.140 37.180 ;
        RECT 130.510 29.210 130.940 36.580 ;
        RECT 131.230 32.720 133.000 36.700 ;
        RECT 131.230 31.720 132.990 32.720 ;
        RECT 128.800 28.745 129.030 28.830 ;
        RECT 129.940 28.745 130.170 28.830 ;
        RECT 130.510 28.540 130.950 29.210 ;
        RECT 131.230 28.840 133.000 31.720 ;
        RECT 135.510 29.600 136.620 36.710 ;
        RECT 131.230 28.745 131.460 28.840 ;
        RECT 126.790 28.310 128.750 28.540 ;
        RECT 130.220 28.310 131.180 28.540 ;
        RECT 130.320 27.430 131.110 28.310 ;
        RECT 131.860 27.830 133.000 28.840 ;
        RECT 126.380 26.560 130.000 27.180 ;
        RECT 130.270 26.670 131.160 27.430 ;
        RECT 120.540 25.530 121.900 25.760 ;
        RECT 120.540 24.360 121.630 25.530 ;
        RECT 122.900 25.370 123.230 26.530 ;
        RECT 123.370 25.530 125.330 25.760 ;
        RECT 117.520 22.270 117.750 22.320 ;
        RECT 117.960 22.270 118.190 22.330 ;
        RECT 113.770 21.600 116.470 21.920 ;
        RECT 113.770 21.370 114.000 21.600 ;
        RECT 110.680 20.750 111.040 21.050 ;
        RECT 111.760 20.980 113.720 21.210 ;
        RECT 114.380 20.750 116.470 21.600 ;
        RECT 120.550 21.410 121.630 24.360 ;
        RECT 120.600 21.210 121.630 21.410 ;
        RECT 121.950 25.360 122.180 25.370 ;
        RECT 121.950 23.050 122.360 25.360 ;
        RECT 122.900 25.350 123.320 25.370 ;
        RECT 122.900 25.300 123.410 25.350 ;
        RECT 123.760 25.300 125.020 25.530 ;
        RECT 126.380 25.370 126.640 26.560 ;
        RECT 129.590 25.910 129.990 26.560 ;
        RECT 131.930 26.510 133.000 27.830 ;
        RECT 135.500 28.540 136.620 29.600 ;
        RECT 136.900 36.540 137.340 36.745 ;
        RECT 138.040 36.720 138.270 36.745 ;
        RECT 138.040 36.710 138.280 36.720 ;
        RECT 136.900 28.800 137.290 36.540 ;
        RECT 137.870 29.650 138.280 36.710 ;
        RECT 138.860 30.360 139.760 36.950 ;
        RECT 140.330 36.700 140.560 36.745 ;
        RECT 141.470 36.720 141.700 36.745 ;
        RECT 137.860 28.830 138.280 29.650 ;
        RECT 138.830 29.350 139.830 30.360 ;
        RECT 136.900 28.745 137.130 28.800 ;
        RECT 137.860 28.745 138.270 28.830 ;
        RECT 135.500 28.310 136.850 28.540 ;
        RECT 135.500 27.670 136.710 28.310 ;
        RECT 131.930 26.010 133.770 26.510 ;
        RECT 135.060 26.420 136.710 27.670 ;
        RECT 130.990 25.910 131.740 25.920 ;
        RECT 129.590 25.860 131.740 25.910 ;
        RECT 129.590 25.820 131.920 25.860 ;
        RECT 126.800 25.530 128.760 25.760 ;
        RECT 129.590 25.570 133.150 25.820 ;
        RECT 129.590 25.560 130.930 25.570 ;
        RECT 130.640 25.540 130.930 25.560 ;
        RECT 121.950 21.370 122.450 23.050 ;
        RECT 122.900 21.440 125.020 25.300 ;
        RECT 123.020 21.430 125.020 21.440 ;
        RECT 123.090 21.370 123.320 21.430 ;
        RECT 120.600 21.030 121.900 21.210 ;
        RECT 120.940 20.980 121.900 21.030 ;
        RECT 122.250 20.750 122.450 21.370 ;
        RECT 123.680 21.210 125.020 21.430 ;
        RECT 125.380 25.330 125.610 25.370 ;
        RECT 126.380 25.340 126.750 25.370 ;
        RECT 126.380 25.330 126.830 25.340 ;
        RECT 125.380 25.320 125.790 25.330 ;
        RECT 125.380 23.100 125.830 25.320 ;
        RECT 125.380 22.610 125.880 23.100 ;
        RECT 125.380 21.940 125.970 22.610 ;
        RECT 125.380 21.690 126.030 21.940 ;
        RECT 125.380 21.660 126.080 21.690 ;
        RECT 125.380 21.370 125.610 21.660 ;
        RECT 125.840 21.290 126.080 21.660 ;
        RECT 126.330 21.430 126.830 25.330 ;
        RECT 126.330 21.420 126.750 21.430 ;
        RECT 126.390 21.410 126.750 21.420 ;
        RECT 126.520 21.370 126.750 21.410 ;
        RECT 123.370 20.980 125.330 21.210 ;
        RECT 125.760 21.050 126.080 21.290 ;
        RECT 127.090 21.210 128.460 25.530 ;
        RECT 131.800 25.480 133.150 25.570 ;
        RECT 132.750 25.475 133.040 25.480 ;
        RECT 128.810 25.190 129.040 25.370 ;
        RECT 130.450 25.320 130.680 25.380 ;
        RECT 130.890 25.320 131.120 25.380 ;
        RECT 129.700 25.310 130.680 25.320 ;
        RECT 129.270 25.190 130.680 25.310 ;
        RECT 128.810 24.440 130.680 25.190 ;
        RECT 130.870 25.180 131.270 25.320 ;
        RECT 133.400 25.270 133.770 26.010 ;
        RECT 132.560 25.180 132.790 25.270 ;
        RECT 130.870 24.450 132.830 25.180 ;
        RECT 130.870 24.440 131.270 24.450 ;
        RECT 128.810 23.980 130.170 24.440 ;
        RECT 130.450 24.380 130.680 24.440 ;
        RECT 130.890 24.380 131.120 24.440 ;
        RECT 128.810 23.710 131.270 23.980 ;
        RECT 128.810 23.670 130.980 23.710 ;
        RECT 128.810 21.920 130.160 23.670 ;
        RECT 131.440 23.490 132.820 24.450 ;
        RECT 131.440 23.360 132.840 23.490 ;
        RECT 130.720 22.360 132.840 23.360 ;
        RECT 131.440 22.330 132.840 22.360 ;
        RECT 132.560 22.320 132.840 22.330 ;
        RECT 133.000 22.330 133.770 25.270 ;
        RECT 135.500 25.760 136.710 26.420 ;
        RECT 137.860 26.530 138.180 28.745 ;
        RECT 138.860 28.540 139.760 29.350 ;
        RECT 140.330 28.810 140.850 36.700 ;
        RECT 140.330 28.745 140.560 28.810 ;
        RECT 141.330 28.800 141.710 36.720 ;
        RECT 142.410 30.320 143.230 36.950 ;
        RECT 143.760 36.700 143.990 36.745 ;
        RECT 144.900 36.700 145.130 36.745 ;
        RECT 142.320 29.320 143.320 30.320 ;
        RECT 141.340 28.745 141.700 28.800 ;
        RECT 138.320 28.310 140.280 28.540 ;
        RECT 141.340 27.180 141.600 28.745 ;
        RECT 142.410 28.540 143.230 29.320 ;
        RECT 143.760 28.830 145.140 36.700 ;
        RECT 145.470 36.580 145.910 36.950 ;
        RECT 146.190 36.700 146.420 36.745 ;
        RECT 146.820 36.700 147.960 37.510 ;
        RECT 145.470 29.210 145.900 36.580 ;
        RECT 146.190 32.720 147.960 36.700 ;
        RECT 146.190 31.720 147.950 32.720 ;
        RECT 143.760 28.745 143.990 28.830 ;
        RECT 144.900 28.745 145.130 28.830 ;
        RECT 145.470 28.540 145.910 29.210 ;
        RECT 146.190 28.840 147.960 31.720 ;
        RECT 146.190 28.745 146.420 28.840 ;
        RECT 141.750 28.310 143.710 28.540 ;
        RECT 145.180 28.310 146.140 28.540 ;
        RECT 145.280 27.430 146.070 28.310 ;
        RECT 146.820 27.830 147.960 28.840 ;
        RECT 141.340 26.560 144.960 27.180 ;
        RECT 145.230 26.670 146.120 27.430 ;
        RECT 135.500 25.530 136.860 25.760 ;
        RECT 135.500 24.360 136.590 25.530 ;
        RECT 137.860 25.370 138.190 26.530 ;
        RECT 138.330 25.530 140.290 25.760 ;
        RECT 132.560 22.270 132.790 22.320 ;
        RECT 133.000 22.270 133.230 22.330 ;
        RECT 128.810 21.600 131.510 21.920 ;
        RECT 128.810 21.370 129.040 21.600 ;
        RECT 125.720 20.750 126.080 21.050 ;
        RECT 126.800 20.980 128.760 21.210 ;
        RECT 129.420 20.750 131.510 21.600 ;
        RECT 135.510 21.410 136.590 24.360 ;
        RECT 135.560 21.210 136.590 21.410 ;
        RECT 136.910 25.360 137.140 25.370 ;
        RECT 136.910 23.050 137.320 25.360 ;
        RECT 137.860 25.350 138.280 25.370 ;
        RECT 137.860 25.300 138.370 25.350 ;
        RECT 138.720 25.300 139.980 25.530 ;
        RECT 141.340 25.370 141.600 26.560 ;
        RECT 144.550 25.910 144.950 26.560 ;
        RECT 146.890 26.510 147.960 27.830 ;
        RECT 146.890 26.010 148.730 26.510 ;
        RECT 145.950 25.910 146.700 25.920 ;
        RECT 144.550 25.860 146.700 25.910 ;
        RECT 144.550 25.820 146.880 25.860 ;
        RECT 141.760 25.530 143.720 25.760 ;
        RECT 144.550 25.570 148.110 25.820 ;
        RECT 144.550 25.560 145.890 25.570 ;
        RECT 145.600 25.540 145.890 25.560 ;
        RECT 136.910 21.370 137.410 23.050 ;
        RECT 137.860 21.440 139.980 25.300 ;
        RECT 137.980 21.430 139.980 21.440 ;
        RECT 138.050 21.370 138.280 21.430 ;
        RECT 135.560 21.030 136.860 21.210 ;
        RECT 135.900 20.980 136.860 21.030 ;
        RECT 137.210 20.750 137.410 21.370 ;
        RECT 138.640 21.210 139.980 21.430 ;
        RECT 140.340 25.330 140.570 25.370 ;
        RECT 141.340 25.340 141.710 25.370 ;
        RECT 141.340 25.330 141.790 25.340 ;
        RECT 140.340 25.320 140.750 25.330 ;
        RECT 140.340 23.100 140.790 25.320 ;
        RECT 140.340 22.610 140.840 23.100 ;
        RECT 140.340 21.940 140.930 22.610 ;
        RECT 140.340 21.690 140.990 21.940 ;
        RECT 140.340 21.660 141.040 21.690 ;
        RECT 140.340 21.370 140.570 21.660 ;
        RECT 140.800 21.290 141.040 21.660 ;
        RECT 141.290 21.430 141.790 25.330 ;
        RECT 141.290 21.420 141.710 21.430 ;
        RECT 141.350 21.410 141.710 21.420 ;
        RECT 141.480 21.370 141.710 21.410 ;
        RECT 138.330 20.980 140.290 21.210 ;
        RECT 140.720 21.050 141.040 21.290 ;
        RECT 142.050 21.210 143.420 25.530 ;
        RECT 146.760 25.480 148.110 25.570 ;
        RECT 147.710 25.475 148.000 25.480 ;
        RECT 143.770 25.190 144.000 25.370 ;
        RECT 145.410 25.320 145.640 25.380 ;
        RECT 145.850 25.320 146.080 25.380 ;
        RECT 144.660 25.310 145.640 25.320 ;
        RECT 144.230 25.190 145.640 25.310 ;
        RECT 143.770 24.440 145.640 25.190 ;
        RECT 145.830 25.180 146.230 25.320 ;
        RECT 148.360 25.270 148.730 26.010 ;
        RECT 147.520 25.180 147.750 25.270 ;
        RECT 145.830 24.450 147.790 25.180 ;
        RECT 145.830 24.440 146.230 24.450 ;
        RECT 143.770 23.980 145.130 24.440 ;
        RECT 145.410 24.380 145.640 24.440 ;
        RECT 145.850 24.380 146.080 24.440 ;
        RECT 143.770 23.710 146.230 23.980 ;
        RECT 143.770 23.670 145.940 23.710 ;
        RECT 143.770 21.920 145.120 23.670 ;
        RECT 146.400 23.490 147.780 24.450 ;
        RECT 146.400 23.360 147.800 23.490 ;
        RECT 145.680 22.360 147.800 23.360 ;
        RECT 146.400 22.330 147.800 22.360 ;
        RECT 143.770 21.600 146.470 21.920 ;
        RECT 143.770 21.370 144.000 21.600 ;
        RECT 140.680 20.750 141.040 21.050 ;
        RECT 141.760 20.980 143.720 21.210 ;
        RECT 144.380 20.750 146.470 21.600 ;
        RECT 74.560 20.720 86.520 20.750 ;
        RECT 90.100 20.730 101.460 20.750 ;
        RECT 105.110 20.730 116.470 20.750 ;
        RECT 120.150 20.730 131.510 20.750 ;
        RECT 90.100 20.720 131.510 20.730 ;
        RECT 74.560 20.670 131.510 20.720 ;
        RECT 135.110 20.670 146.470 20.750 ;
        RECT 74.560 20.000 146.470 20.670 ;
        RECT 74.560 19.990 101.450 20.000 ;
        RECT 74.560 19.920 86.510 19.990 ;
        RECT 90.070 19.920 101.450 19.990 ;
        RECT 105.080 19.920 116.460 20.000 ;
        RECT 120.120 19.940 146.460 20.000 ;
        RECT 120.120 19.920 131.500 19.940 ;
        RECT 135.080 19.920 146.460 19.940 ;
        RECT 74.560 19.910 75.300 19.920 ;
        RECT 61.490 19.300 62.490 19.320 ;
        RECT 61.490 18.870 63.290 19.300 ;
        RECT 63.510 19.170 66.780 19.370 ;
        RECT 63.510 19.160 66.340 19.170 ;
        RECT 63.510 19.010 66.260 19.160 ;
        RECT 66.520 18.870 66.780 18.910 ;
        RECT 61.490 18.320 66.780 18.870 ;
        RECT 61.500 18.310 66.780 18.320 ;
        RECT 116.010 18.085 116.410 18.180 ;
        RECT 60.515 17.875 116.410 18.085 ;
        RECT 116.010 17.780 116.410 17.875 ;
        RECT 146.830 17.620 147.045 22.330 ;
        RECT 147.520 22.320 147.800 22.330 ;
        RECT 147.960 22.330 148.730 25.270 ;
        RECT 147.520 22.270 147.750 22.320 ;
        RECT 147.960 22.270 148.190 22.330 ;
        RECT 60.020 17.405 147.045 17.620 ;
      LAYER met2 ;
        RECT 33.300 224.810 33.870 225.380 ;
        RECT 63.670 225.040 64.140 225.560 ;
        RECT 63.830 224.310 63.970 225.040 ;
        RECT 71.910 224.880 72.380 225.650 ;
        RECT 74.640 224.940 75.350 225.590 ;
        RECT 57.290 224.170 63.970 224.310 ;
        RECT 57.290 223.370 57.430 224.170 ;
        RECT 72.035 223.895 72.305 224.880 ;
        RECT 77.450 224.860 78.030 225.470 ;
        RECT 80.190 224.880 80.730 225.500 ;
        RECT 82.970 224.880 83.500 225.440 ;
        RECT 83.135 224.055 83.340 224.880 ;
        RECT 85.640 224.780 86.400 225.570 ;
        RECT 88.520 225.060 89.040 225.620 ;
        RECT 91.220 224.940 91.850 225.620 ;
        RECT 93.980 224.910 94.550 225.440 ;
        RECT 85.820 224.125 86.095 224.780 ;
        RECT 132.450 224.710 133.340 225.530 ;
        RECT 135.310 224.910 136.020 225.580 ;
        RECT 137.980 224.970 138.430 225.420 ;
        RECT 140.930 224.920 141.430 225.440 ;
        RECT 11.990 223.230 57.430 223.370 ;
        RECT 58.065 223.625 72.305 223.895 ;
        RECT 75.030 223.850 83.340 224.055 ;
        RECT 83.840 223.920 86.095 224.125 ;
        RECT 125.800 223.980 126.280 224.400 ;
        RECT 11.990 138.470 12.130 223.230 ;
        RECT 58.065 222.855 58.335 223.625 ;
        RECT 75.030 223.320 75.235 223.850 ;
        RECT 83.900 223.675 84.105 223.920 ;
        RECT 84.260 223.850 86.095 223.920 ;
        RECT 75.530 223.510 84.105 223.675 ;
        RECT 132.580 223.670 133.040 224.710 ;
        RECT 75.530 223.470 79.300 223.510 ;
        RECT 79.900 223.470 84.105 223.510 ;
        RECT 12.465 222.585 58.335 222.855 ;
        RECT 58.715 223.115 75.270 223.320 ;
        RECT 12.465 139.685 12.735 222.585 ;
        RECT 58.715 222.360 58.920 223.115 ;
        RECT 14.575 222.155 58.920 222.360 ;
        RECT 59.325 222.905 75.270 222.910 ;
        RECT 75.530 222.905 75.735 223.470 ;
        RECT 79.450 222.975 79.750 223.365 ;
        RECT 84.540 223.210 133.040 223.670 ;
        RECT 59.325 222.700 75.735 222.905 ;
        RECT 59.325 222.645 75.270 222.700 ;
        RECT 13.500 143.750 14.200 144.420 ;
        RECT 13.150 140.350 14.220 141.070 ;
        RECT 12.465 139.415 14.005 139.685 ;
        RECT 11.990 138.330 13.230 138.470 ;
        RECT 12.295 135.665 12.595 136.055 ;
        RECT 12.345 119.425 12.540 135.665 ;
        RECT 13.090 129.350 13.230 138.330 ;
        RECT 13.735 130.565 14.005 139.415 ;
        RECT 14.575 131.415 14.890 222.155 ;
        RECT 59.325 221.900 59.590 222.645 ;
        RECT 63.800 222.300 64.270 222.390 ;
        RECT 60.740 222.290 64.270 222.300 ;
        RECT 15.350 221.635 59.590 221.900 ;
        RECT 60.210 222.020 64.270 222.290 ;
        RECT 79.530 222.140 79.670 222.975 ;
        RECT 84.540 222.230 85.000 223.210 ;
        RECT 135.500 222.660 135.780 224.910 ;
        RECT 136.550 223.930 137.150 224.410 ;
        RECT 94.890 222.410 135.780 222.660 ;
        RECT 94.890 222.380 95.820 222.410 ;
        RECT 96.450 222.380 135.780 222.410 ;
        RECT 15.350 132.210 15.615 221.635 ;
        RECT 32.820 221.085 34.360 221.455 ;
        RECT 15.970 220.585 16.360 220.620 ;
        RECT 15.970 220.350 16.905 220.585 ;
        RECT 15.970 220.320 16.360 220.350 ;
        RECT 15.990 162.800 16.250 163.120 ;
        RECT 16.050 161.955 16.190 162.800 ;
        RECT 15.980 161.585 16.260 161.955 ;
        RECT 16.670 159.575 16.905 220.350 ;
        RECT 60.210 219.900 60.350 222.020 ;
        RECT 63.800 221.910 64.270 222.020 ;
        RECT 75.670 221.860 79.670 222.140 ;
        RECT 79.530 220.580 79.670 221.860 ;
        RECT 80.850 222.220 82.590 222.230 ;
        RECT 83.080 222.220 85.170 222.230 ;
        RECT 80.850 221.770 85.170 222.220 ;
        RECT 85.960 221.920 89.960 222.160 ;
        RECT 94.890 221.920 95.170 222.380 ;
        RECT 95.960 222.160 96.290 222.270 ;
        RECT 96.750 222.160 99.610 222.180 ;
        RECT 85.960 221.880 95.170 221.920 ;
        RECT 95.610 221.900 99.610 222.160 ;
        RECT 82.740 221.600 82.920 221.770 ;
        RECT 79.470 220.260 79.730 220.580 ;
        RECT 82.750 219.900 82.890 221.600 ;
        RECT 85.970 220.240 86.110 221.880 ;
        RECT 89.660 221.640 95.170 221.880 ;
        RECT 95.630 220.580 95.770 221.900 ;
        RECT 141.110 221.850 141.250 224.920 ;
        RECT 141.110 221.710 147.570 221.850 ;
        RECT 87.750 220.260 88.010 220.580 ;
        RECT 95.570 220.260 95.830 220.580 ;
        RECT 85.910 219.920 86.170 220.240 ;
        RECT 60.150 219.580 60.410 219.900 ;
        RECT 82.690 219.580 82.950 219.900 ;
        RECT 87.290 219.580 87.550 219.900 ;
        RECT 51.870 219.240 52.130 219.560 ;
        RECT 84.530 219.240 84.790 219.560 ;
        RECT 36.120 218.365 37.660 218.735 ;
        RECT 32.820 215.645 34.360 216.015 ;
        RECT 50.950 214.820 51.210 215.140 ;
        RECT 49.110 213.460 49.370 213.780 ;
        RECT 36.120 212.925 37.660 213.295 ;
        RECT 49.170 212.760 49.310 213.460 ;
        RECT 49.110 212.440 49.370 212.760 ;
        RECT 45.430 212.100 45.690 212.420 ;
        RECT 32.820 210.205 34.360 210.575 ;
        RECT 45.490 209.360 45.630 212.100 ;
        RECT 50.490 211.760 50.750 212.080 ;
        RECT 45.890 210.740 46.150 211.060 ;
        RECT 43.590 209.040 43.850 209.360 ;
        RECT 45.430 209.040 45.690 209.360 ;
        RECT 36.120 207.485 37.660 207.855 ;
        RECT 32.820 204.765 34.360 205.135 ;
        RECT 42.670 203.940 42.930 204.260 ;
        RECT 21.510 203.260 21.770 203.580 ;
        RECT 26.110 203.260 26.370 203.580 ;
        RECT 32.090 203.260 32.350 203.580 ;
        RECT 21.570 201.540 21.710 203.260 ;
        RECT 21.510 201.220 21.770 201.540 ;
        RECT 18.750 200.880 19.010 201.200 ;
        RECT 18.810 198.675 18.950 200.880 ;
        RECT 18.740 198.305 19.020 198.675 ;
        RECT 21.570 196.440 21.710 201.220 ;
        RECT 25.190 200.880 25.450 201.200 ;
        RECT 25.650 200.880 25.910 201.200 ;
        RECT 24.730 200.200 24.990 200.520 ;
        RECT 23.810 199.860 24.070 200.180 ;
        RECT 22.890 197.480 23.150 197.800 ;
        RECT 21.510 196.120 21.770 196.440 ;
        RECT 22.950 193.720 23.090 197.480 ;
        RECT 23.870 196.100 24.010 199.860 ;
        RECT 23.810 195.780 24.070 196.100 ;
        RECT 22.890 193.400 23.150 193.720 ;
        RECT 24.790 192.360 24.930 200.200 ;
        RECT 25.250 198.140 25.390 200.880 ;
        RECT 25.190 197.820 25.450 198.140 ;
        RECT 25.250 196.440 25.390 197.820 ;
        RECT 25.190 196.120 25.450 196.440 ;
        RECT 24.730 192.040 24.990 192.360 ;
        RECT 24.790 187.940 24.930 192.040 ;
        RECT 25.710 192.020 25.850 200.880 ;
        RECT 26.170 197.800 26.310 203.260 ;
        RECT 28.870 202.920 29.130 203.240 ;
        RECT 27.030 202.580 27.290 202.900 ;
        RECT 26.110 197.480 26.370 197.800 ;
        RECT 26.110 194.420 26.370 194.740 ;
        RECT 26.170 193.040 26.310 194.420 ;
        RECT 27.090 193.720 27.230 202.580 ;
        RECT 28.930 198.140 29.070 202.920 ;
        RECT 32.150 200.520 32.290 203.260 ;
        RECT 39.450 202.920 39.710 203.240 ;
        RECT 36.120 202.045 37.660 202.415 ;
        RECT 39.510 201.880 39.650 202.920 ;
        RECT 39.910 202.580 40.170 202.900 ;
        RECT 39.450 201.560 39.710 201.880 ;
        RECT 35.770 200.880 36.030 201.200 ;
        RECT 32.090 200.430 32.350 200.520 ;
        RECT 31.690 200.290 32.350 200.430 ;
        RECT 31.690 198.140 31.830 200.290 ;
        RECT 32.090 200.200 32.350 200.290 ;
        RECT 32.820 199.325 34.360 199.695 ;
        RECT 35.830 199.160 35.970 200.880 ;
        RECT 39.970 200.600 40.110 202.580 ;
        RECT 40.830 200.880 41.090 201.200 ;
        RECT 39.510 200.460 40.110 200.600 ;
        RECT 39.510 200.430 39.650 200.460 ;
        RECT 39.050 200.290 39.650 200.430 ;
        RECT 39.050 200.035 39.190 200.290 ;
        RECT 40.370 200.200 40.630 200.520 ;
        RECT 39.910 200.090 40.170 200.180 ;
        RECT 38.980 199.665 39.260 200.035 ;
        RECT 39.510 199.950 40.170 200.090 ;
        RECT 35.770 198.840 36.030 199.160 ;
        RECT 39.050 198.140 39.190 199.665 ;
        RECT 28.870 197.820 29.130 198.140 ;
        RECT 31.630 197.820 31.890 198.140 ;
        RECT 32.550 197.880 32.810 198.140 ;
        RECT 33.930 197.880 34.190 198.140 ;
        RECT 32.550 197.820 34.190 197.880 ;
        RECT 38.990 197.820 39.250 198.140 ;
        RECT 28.410 197.140 28.670 197.460 ;
        RECT 28.470 195.760 28.610 197.140 ;
        RECT 28.930 196.440 29.070 197.820 ;
        RECT 30.710 197.140 30.970 197.460 ;
        RECT 28.870 196.120 29.130 196.440 ;
        RECT 28.410 195.440 28.670 195.760 ;
        RECT 28.930 195.420 29.070 196.120 ;
        RECT 28.870 195.100 29.130 195.420 ;
        RECT 27.490 194.420 27.750 194.740 ;
        RECT 27.030 193.400 27.290 193.720 ;
        RECT 26.110 192.720 26.370 193.040 ;
        RECT 25.650 191.700 25.910 192.020 ;
        RECT 25.650 190.000 25.910 190.320 ;
        RECT 24.730 187.620 24.990 187.940 ;
        RECT 25.710 186.920 25.850 190.000 ;
        RECT 26.170 189.980 26.310 192.720 ;
        RECT 27.550 192.700 27.690 194.420 ;
        RECT 27.490 192.380 27.750 192.700 ;
        RECT 30.770 192.020 30.910 197.140 ;
        RECT 31.690 196.100 31.830 197.820 ;
        RECT 32.090 197.480 32.350 197.800 ;
        RECT 32.610 197.740 34.130 197.820 ;
        RECT 31.630 196.010 31.890 196.100 ;
        RECT 31.230 195.870 31.890 196.010 ;
        RECT 31.230 195.420 31.370 195.870 ;
        RECT 31.630 195.780 31.890 195.870 ;
        RECT 31.170 195.100 31.430 195.420 ;
        RECT 31.230 194.740 31.370 195.100 ;
        RECT 31.170 194.420 31.430 194.740 ;
        RECT 32.150 192.360 32.290 197.480 ;
        RECT 32.610 197.460 32.750 197.740 ;
        RECT 32.550 197.140 32.810 197.460 ;
        RECT 32.610 195.080 32.750 197.140 ;
        RECT 36.120 196.605 37.660 196.975 ;
        RECT 35.770 195.440 36.030 195.760 ;
        RECT 37.150 195.440 37.410 195.760 ;
        RECT 38.530 195.440 38.790 195.760 ;
        RECT 32.550 194.760 32.810 195.080 ;
        RECT 34.850 194.760 35.110 195.080 ;
        RECT 32.820 193.885 34.360 194.255 ;
        RECT 32.090 192.040 32.350 192.360 ;
        RECT 30.710 191.700 30.970 192.020 ;
        RECT 26.110 189.660 26.370 189.980 ;
        RECT 26.170 187.260 26.310 189.660 ;
        RECT 34.910 189.640 35.050 194.760 ;
        RECT 35.310 193.400 35.570 193.720 ;
        RECT 35.370 191.000 35.510 193.400 ;
        RECT 35.830 192.700 35.970 195.440 ;
        RECT 37.210 194.740 37.350 195.440 ;
        RECT 37.150 194.420 37.410 194.740 ;
        RECT 35.770 192.380 36.030 192.700 ;
        RECT 35.310 190.680 35.570 191.000 ;
        RECT 35.830 190.660 35.970 192.380 ;
        RECT 37.210 192.360 37.350 194.420 ;
        RECT 38.590 192.700 38.730 195.440 ;
        RECT 39.050 193.720 39.190 197.820 ;
        RECT 39.510 195.760 39.650 199.950 ;
        RECT 39.910 199.860 40.170 199.950 ;
        RECT 40.430 198.820 40.570 200.200 ;
        RECT 40.370 198.500 40.630 198.820 ;
        RECT 40.430 195.760 40.570 198.500 ;
        RECT 40.890 198.140 41.030 200.880 ;
        RECT 42.730 200.180 42.870 203.940 ;
        RECT 43.650 201.540 43.790 209.040 ;
        RECT 45.950 208.680 46.090 210.740 ;
        RECT 45.890 208.360 46.150 208.680 ;
        RECT 50.550 207.320 50.690 211.760 ;
        RECT 50.490 207.000 50.750 207.320 ;
        RECT 51.010 206.640 51.150 214.820 ;
        RECT 50.950 206.320 51.210 206.640 ;
        RECT 50.490 205.640 50.750 205.960 ;
        RECT 43.590 201.220 43.850 201.540 ;
        RECT 46.350 201.220 46.610 201.540 ;
        RECT 43.130 200.540 43.390 200.860 ;
        RECT 42.670 199.860 42.930 200.180 ;
        RECT 40.830 197.820 41.090 198.140 ;
        RECT 41.290 197.480 41.550 197.800 ;
        RECT 41.350 195.760 41.490 197.480 ;
        RECT 42.730 195.840 42.870 199.860 ;
        RECT 43.190 198.140 43.330 200.540 ;
        RECT 43.130 197.820 43.390 198.140 ;
        RECT 43.190 196.440 43.330 197.820 ;
        RECT 43.130 196.120 43.390 196.440 ;
        RECT 39.450 195.440 39.710 195.760 ;
        RECT 40.370 195.440 40.630 195.760 ;
        RECT 41.290 195.440 41.550 195.760 ;
        RECT 42.730 195.700 43.330 195.840 ;
        RECT 43.190 195.420 43.330 195.700 ;
        RECT 39.910 195.100 40.170 195.420 ;
        RECT 43.130 195.100 43.390 195.420 ;
        RECT 38.990 193.400 39.250 193.720 ;
        RECT 38.530 192.380 38.790 192.700 ;
        RECT 39.450 192.380 39.710 192.700 ;
        RECT 37.150 192.040 37.410 192.360 ;
        RECT 36.120 191.165 37.660 191.535 ;
        RECT 36.230 190.680 36.490 191.000 ;
        RECT 35.770 190.340 36.030 190.660 ;
        RECT 35.310 190.000 35.570 190.320 ;
        RECT 34.850 189.320 35.110 189.640 ;
        RECT 29.330 188.980 29.590 189.300 ;
        RECT 27.950 187.620 28.210 187.940 ;
        RECT 26.110 186.940 26.370 187.260 ;
        RECT 27.030 186.940 27.290 187.260 ;
        RECT 25.650 186.600 25.910 186.920 ;
        RECT 22.430 186.260 22.690 186.580 ;
        RECT 22.490 185.220 22.630 186.260 ;
        RECT 22.430 184.900 22.690 185.220 ;
        RECT 25.710 183.860 25.850 186.600 ;
        RECT 26.170 184.880 26.310 186.940 ;
        RECT 27.090 185.220 27.230 186.940 ;
        RECT 27.030 184.900 27.290 185.220 ;
        RECT 26.110 184.560 26.370 184.880 ;
        RECT 26.570 183.880 26.830 184.200 ;
        RECT 25.190 183.540 25.450 183.860 ;
        RECT 25.650 183.540 25.910 183.860 ;
        RECT 25.250 181.820 25.390 183.540 ;
        RECT 25.710 182.840 25.850 183.540 ;
        RECT 25.650 182.520 25.910 182.840 ;
        RECT 25.190 181.500 25.450 181.820 ;
        RECT 21.050 175.380 21.310 175.700 ;
        RECT 19.210 170.620 19.470 170.940 ;
        RECT 19.270 168.560 19.410 170.620 ;
        RECT 20.130 169.940 20.390 170.260 ;
        RECT 20.190 169.240 20.330 169.940 ;
        RECT 20.130 168.920 20.390 169.240 ;
        RECT 19.210 168.240 19.470 168.560 ;
        RECT 21.110 167.540 21.250 175.380 ;
        RECT 21.970 174.020 22.230 174.340 ;
        RECT 21.510 172.660 21.770 172.980 ;
        RECT 21.570 169.240 21.710 172.660 ;
        RECT 22.030 170.260 22.170 174.020 ;
        RECT 23.350 172.890 23.610 172.980 ;
        RECT 23.350 172.750 24.010 172.890 ;
        RECT 23.350 172.660 23.610 172.750 ;
        RECT 21.970 169.940 22.230 170.260 ;
        RECT 21.510 168.920 21.770 169.240 ;
        RECT 22.030 168.900 22.170 169.940 ;
        RECT 23.870 168.900 24.010 172.750 ;
        RECT 25.250 169.240 25.390 181.500 ;
        RECT 26.630 176.380 26.770 183.880 ;
        RECT 26.570 176.060 26.830 176.380 ;
        RECT 26.630 174.340 26.770 176.060 ;
        RECT 27.490 175.720 27.750 176.040 ;
        RECT 26.570 174.020 26.830 174.340 ;
        RECT 27.550 174.000 27.690 175.720 ;
        RECT 27.490 173.680 27.750 174.000 ;
        RECT 26.110 173.000 26.370 173.320 ;
        RECT 26.170 171.960 26.310 173.000 ;
        RECT 27.030 172.660 27.290 172.980 ;
        RECT 27.090 171.960 27.230 172.660 ;
        RECT 26.110 171.640 26.370 171.960 ;
        RECT 27.030 171.640 27.290 171.960 ;
        RECT 27.550 170.940 27.690 173.680 ;
        RECT 27.490 170.620 27.750 170.940 ;
        RECT 27.490 170.000 27.750 170.260 ;
        RECT 28.010 170.000 28.150 187.620 ;
        RECT 29.390 187.260 29.530 188.980 ;
        RECT 32.820 188.445 34.360 188.815 ;
        RECT 32.090 187.960 32.350 188.280 ;
        RECT 31.170 187.620 31.430 187.940 ;
        RECT 30.250 187.280 30.510 187.600 ;
        RECT 29.330 186.940 29.590 187.260 ;
        RECT 29.390 184.280 29.530 186.940 ;
        RECT 30.310 185.560 30.450 187.280 ;
        RECT 30.250 185.240 30.510 185.560 ;
        RECT 31.230 185.220 31.370 187.620 ;
        RECT 32.150 185.560 32.290 187.960 ;
        RECT 35.370 187.260 35.510 190.000 ;
        RECT 35.770 189.660 36.030 189.980 ;
        RECT 35.830 187.260 35.970 189.660 ;
        RECT 35.310 186.940 35.570 187.260 ;
        RECT 35.770 186.940 36.030 187.260 ;
        RECT 36.290 186.490 36.430 190.680 ;
        RECT 39.510 189.980 39.650 192.380 ;
        RECT 39.970 190.320 40.110 195.100 ;
        RECT 40.830 194.760 41.090 195.080 ;
        RECT 40.370 194.420 40.630 194.740 ;
        RECT 40.430 192.700 40.570 194.420 ;
        RECT 40.370 192.380 40.630 192.700 ;
        RECT 40.890 192.360 41.030 194.760 ;
        RECT 42.670 194.420 42.930 194.740 ;
        RECT 42.210 192.440 42.470 192.700 ;
        RECT 42.730 192.440 42.870 194.420 ;
        RECT 43.190 193.380 43.330 195.100 ;
        RECT 43.130 193.060 43.390 193.380 ;
        RECT 42.210 192.380 42.870 192.440 ;
        RECT 40.830 192.040 41.090 192.360 ;
        RECT 42.270 192.300 42.870 192.380 ;
        RECT 41.290 191.700 41.550 192.020 ;
        RECT 41.750 191.700 42.010 192.020 ;
        RECT 41.350 190.320 41.490 191.700 ;
        RECT 41.810 190.660 41.950 191.700 ;
        RECT 41.750 190.340 42.010 190.660 ;
        RECT 39.910 190.000 40.170 190.320 ;
        RECT 41.290 190.000 41.550 190.320 ;
        RECT 39.450 189.660 39.710 189.980 ;
        RECT 36.690 189.320 36.950 189.640 ;
        RECT 36.750 187.260 36.890 189.320 ;
        RECT 39.450 188.980 39.710 189.300 ;
        RECT 36.690 186.940 36.950 187.260 ;
        RECT 37.610 186.940 37.870 187.260 ;
        RECT 38.530 186.940 38.790 187.260 ;
        RECT 37.670 186.580 37.810 186.940 ;
        RECT 35.830 186.350 36.430 186.490 ;
        RECT 32.090 185.240 32.350 185.560 ;
        RECT 31.170 184.900 31.430 185.220 ;
        RECT 29.390 184.140 29.990 184.280 ;
        RECT 34.850 184.220 35.110 184.540 ;
        RECT 29.850 183.860 29.990 184.140 ;
        RECT 29.330 183.540 29.590 183.860 ;
        RECT 29.790 183.540 30.050 183.860 ;
        RECT 29.390 181.480 29.530 183.540 ;
        RECT 32.820 183.005 34.360 183.375 ;
        RECT 29.330 181.160 29.590 181.480 ;
        RECT 34.910 179.440 35.050 184.220 ;
        RECT 34.850 179.120 35.110 179.440 ;
        RECT 32.820 177.565 34.360 177.935 ;
        RECT 29.330 176.740 29.590 177.060 ;
        RECT 28.870 175.380 29.130 175.700 ;
        RECT 28.930 174.000 29.070 175.380 ;
        RECT 29.390 174.000 29.530 176.740 ;
        RECT 33.930 176.060 34.190 176.380 ;
        RECT 31.630 175.720 31.890 176.040 ;
        RECT 28.870 173.680 29.130 174.000 ;
        RECT 29.330 173.680 29.590 174.000 ;
        RECT 28.410 173.340 28.670 173.660 ;
        RECT 28.470 170.260 28.610 173.340 ;
        RECT 28.930 171.960 29.070 173.680 ;
        RECT 31.690 173.660 31.830 175.720 ;
        RECT 33.990 174.680 34.130 176.060 ;
        RECT 33.930 174.360 34.190 174.680 ;
        RECT 32.090 173.680 32.350 174.000 ;
        RECT 31.630 173.340 31.890 173.660 ;
        RECT 30.710 172.660 30.970 172.980 ;
        RECT 31.630 172.660 31.890 172.980 ;
        RECT 28.870 171.640 29.130 171.960 ;
        RECT 27.490 169.940 28.150 170.000 ;
        RECT 28.410 169.940 28.670 170.260 ;
        RECT 27.550 169.860 28.150 169.940 ;
        RECT 25.190 168.920 25.450 169.240 ;
        RECT 28.010 168.900 28.150 169.860 ;
        RECT 21.970 168.580 22.230 168.900 ;
        RECT 23.810 168.580 24.070 168.900 ;
        RECT 27.950 168.580 28.210 168.900 ;
        RECT 28.930 167.880 29.070 171.640 ;
        RECT 30.250 170.620 30.510 170.940 ;
        RECT 29.790 170.280 30.050 170.600 ;
        RECT 29.850 168.900 29.990 170.280 ;
        RECT 30.310 169.240 30.450 170.620 ;
        RECT 30.770 169.240 30.910 172.660 ;
        RECT 30.250 168.920 30.510 169.240 ;
        RECT 30.710 168.920 30.970 169.240 ;
        RECT 29.790 168.580 30.050 168.900 ;
        RECT 28.870 167.560 29.130 167.880 ;
        RECT 31.690 167.540 31.830 172.660 ;
        RECT 32.150 171.960 32.290 173.680 ;
        RECT 34.910 173.320 35.050 179.120 ;
        RECT 35.310 175.720 35.570 176.040 ;
        RECT 35.370 173.660 35.510 175.720 ;
        RECT 35.830 174.680 35.970 186.350 ;
        RECT 37.610 186.260 37.870 186.580 ;
        RECT 38.070 186.260 38.330 186.580 ;
        RECT 36.120 185.725 37.660 186.095 ;
        RECT 38.130 184.960 38.270 186.260 ;
        RECT 38.590 185.220 38.730 186.940 ;
        RECT 38.990 185.240 39.250 185.560 ;
        RECT 37.670 184.880 38.270 184.960 ;
        RECT 38.530 184.900 38.790 185.220 ;
        RECT 37.610 184.820 38.270 184.880 ;
        RECT 37.610 184.560 37.870 184.820 ;
        RECT 38.530 183.540 38.790 183.860 ;
        RECT 38.590 182.500 38.730 183.540 ;
        RECT 38.530 182.180 38.790 182.500 ;
        RECT 38.070 181.500 38.330 181.820 ;
        RECT 36.120 180.285 37.660 180.655 ;
        RECT 38.130 180.120 38.270 181.500 ;
        RECT 37.150 179.800 37.410 180.120 ;
        RECT 38.070 179.800 38.330 180.120 ;
        RECT 36.230 179.120 36.490 179.440 ;
        RECT 36.290 177.400 36.430 179.120 ;
        RECT 37.210 177.400 37.350 179.800 ;
        RECT 38.530 179.120 38.790 179.440 ;
        RECT 36.230 177.080 36.490 177.400 ;
        RECT 37.150 177.080 37.410 177.400 ;
        RECT 38.590 177.060 38.730 179.120 ;
        RECT 39.050 178.420 39.190 185.240 ;
        RECT 39.510 181.820 39.650 188.980 ;
        RECT 42.270 188.280 42.410 192.300 ;
        RECT 42.670 190.000 42.930 190.320 ;
        RECT 42.210 187.960 42.470 188.280 ;
        RECT 39.910 186.940 40.170 187.260 ;
        RECT 39.970 185.560 40.110 186.940 ;
        RECT 40.370 186.600 40.630 186.920 ;
        RECT 39.910 185.240 40.170 185.560 ;
        RECT 40.430 184.540 40.570 186.600 ;
        RECT 42.730 184.880 42.870 190.000 ;
        RECT 42.670 184.560 42.930 184.880 ;
        RECT 40.370 184.220 40.630 184.540 ;
        RECT 39.910 183.880 40.170 184.200 ;
        RECT 39.970 182.500 40.110 183.880 ;
        RECT 39.910 182.180 40.170 182.500 ;
        RECT 39.450 181.500 39.710 181.820 ;
        RECT 39.970 180.120 40.110 182.180 ;
        RECT 43.190 181.820 43.330 193.060 ;
        RECT 43.650 187.600 43.790 201.220 ;
        RECT 44.970 200.880 45.230 201.200 ;
        RECT 45.430 200.880 45.690 201.200 ;
        RECT 45.030 195.760 45.170 200.880 ;
        RECT 45.490 197.800 45.630 200.880 ;
        RECT 46.410 198.820 46.550 201.220 ;
        RECT 46.350 198.500 46.610 198.820 ;
        RECT 45.890 198.160 46.150 198.480 ;
        RECT 45.430 197.480 45.690 197.800 ;
        RECT 44.970 195.440 45.230 195.760 ;
        RECT 45.030 195.160 45.170 195.440 ;
        RECT 44.110 195.020 45.170 195.160 ;
        RECT 44.110 191.000 44.250 195.020 ;
        RECT 45.490 193.020 45.630 197.480 ;
        RECT 45.950 193.380 46.090 198.160 ;
        RECT 46.410 197.800 46.550 198.500 ;
        RECT 50.550 198.480 50.690 205.640 ;
        RECT 51.410 205.300 51.670 205.620 ;
        RECT 51.470 201.880 51.610 205.300 ;
        RECT 51.410 201.560 51.670 201.880 ;
        RECT 51.930 201.540 52.070 219.240 ;
        RECT 55.090 217.880 55.350 218.200 ;
        RECT 55.150 217.520 55.290 217.880 ;
        RECT 64.290 217.540 64.550 217.860 ;
        RECT 53.710 217.200 53.970 217.520 ;
        RECT 55.090 217.200 55.350 217.520 ;
        RECT 60.610 217.200 60.870 217.520 ;
        RECT 52.330 216.860 52.590 217.180 ;
        RECT 52.390 206.640 52.530 216.860 ;
        RECT 53.250 214.480 53.510 214.800 ;
        RECT 53.310 211.060 53.450 214.480 ;
        RECT 53.250 210.740 53.510 211.060 ;
        RECT 53.310 209.020 53.450 210.740 ;
        RECT 53.770 210.040 53.910 217.200 ;
        RECT 54.170 216.180 54.430 216.500 ;
        RECT 54.230 212.080 54.370 216.180 ;
        RECT 54.630 214.140 54.890 214.460 ;
        RECT 54.170 211.760 54.430 212.080 ;
        RECT 53.710 209.720 53.970 210.040 ;
        RECT 53.250 208.700 53.510 209.020 ;
        RECT 54.170 208.700 54.430 209.020 ;
        RECT 52.330 206.320 52.590 206.640 ;
        RECT 52.790 203.600 53.050 203.920 ;
        RECT 52.850 201.880 52.990 203.600 ;
        RECT 54.230 203.580 54.370 208.700 ;
        RECT 54.690 208.680 54.830 214.140 ;
        RECT 55.150 211.060 55.290 217.200 ;
        RECT 56.930 216.860 57.190 217.180 ;
        RECT 55.550 216.180 55.810 216.500 ;
        RECT 55.610 214.460 55.750 216.180 ;
        RECT 56.990 215.480 57.130 216.860 ;
        RECT 60.150 216.520 60.410 216.840 ;
        RECT 56.930 215.160 57.190 215.480 ;
        RECT 55.550 214.140 55.810 214.460 ;
        RECT 55.090 210.740 55.350 211.060 ;
        RECT 56.990 208.680 57.130 215.160 ;
        RECT 59.690 211.080 59.950 211.400 ;
        RECT 59.750 209.700 59.890 211.080 ;
        RECT 59.690 209.610 59.950 209.700 ;
        RECT 59.290 209.470 59.950 209.610 ;
        RECT 59.290 208.680 59.430 209.470 ;
        RECT 59.690 209.380 59.950 209.470 ;
        RECT 60.210 209.360 60.350 216.520 ;
        RECT 60.670 210.040 60.810 217.200 ;
        RECT 64.350 213.780 64.490 217.540 ;
        RECT 68.430 217.200 68.690 217.520 ;
        RECT 68.890 217.200 69.150 217.520 ;
        RECT 70.730 217.200 70.990 217.520 ;
        RECT 65.210 216.180 65.470 216.500 ;
        RECT 64.290 213.460 64.550 213.780 ;
        RECT 61.070 210.740 61.330 211.060 ;
        RECT 60.610 209.720 60.870 210.040 ;
        RECT 60.150 209.040 60.410 209.360 ;
        RECT 61.130 209.020 61.270 210.740 ;
        RECT 62.910 209.040 63.170 209.360 ;
        RECT 61.070 208.700 61.330 209.020 ;
        RECT 61.530 208.700 61.790 209.020 ;
        RECT 54.630 208.360 54.890 208.680 ;
        RECT 56.470 208.360 56.730 208.680 ;
        RECT 56.930 208.360 57.190 208.680 ;
        RECT 59.230 208.360 59.490 208.680 ;
        RECT 59.690 208.360 59.950 208.680 ;
        RECT 56.530 206.640 56.670 208.360 ;
        RECT 56.470 206.320 56.730 206.640 ;
        RECT 56.990 204.000 57.130 208.360 ;
        RECT 58.310 208.020 58.570 208.340 ;
        RECT 56.530 203.860 57.130 204.000 ;
        RECT 54.170 203.260 54.430 203.580 ;
        RECT 56.530 203.320 56.670 203.860 ;
        RECT 53.710 202.920 53.970 203.240 ;
        RECT 52.790 201.560 53.050 201.880 ;
        RECT 51.870 201.220 52.130 201.540 ;
        RECT 51.870 200.540 52.130 200.860 ;
        RECT 50.490 198.160 50.750 198.480 ;
        RECT 46.350 197.480 46.610 197.800 ;
        RECT 46.410 195.420 46.550 197.480 ;
        RECT 46.810 197.140 47.070 197.460 ;
        RECT 46.870 196.100 47.010 197.140 ;
        RECT 46.810 195.780 47.070 196.100 ;
        RECT 46.350 195.100 46.610 195.420 ;
        RECT 45.890 193.060 46.150 193.380 ;
        RECT 45.030 192.880 45.630 193.020 ;
        RECT 45.030 192.020 45.170 192.880 ;
        RECT 45.950 192.360 46.090 193.060 ;
        RECT 46.410 192.700 46.550 195.100 ;
        RECT 50.550 194.740 50.690 198.160 ;
        RECT 51.930 196.440 52.070 200.540 ;
        RECT 52.330 200.035 52.590 200.180 ;
        RECT 52.320 199.665 52.600 200.035 ;
        RECT 53.250 199.860 53.510 200.180 ;
        RECT 52.330 197.820 52.590 198.140 ;
        RECT 51.870 196.120 52.130 196.440 ;
        RECT 52.390 195.760 52.530 197.820 ;
        RECT 53.310 197.460 53.450 199.860 ;
        RECT 53.250 197.140 53.510 197.460 ;
        RECT 53.770 196.100 53.910 202.920 ;
        RECT 54.230 201.200 54.370 203.260 ;
        RECT 56.070 203.240 56.670 203.320 ;
        RECT 56.010 203.180 56.670 203.240 ;
        RECT 56.010 202.920 56.270 203.180 ;
        RECT 55.090 202.580 55.350 202.900 ;
        RECT 55.150 201.880 55.290 202.580 ;
        RECT 55.090 201.560 55.350 201.880 ;
        RECT 54.170 200.880 54.430 201.200 ;
        RECT 54.630 200.200 54.890 200.520 ;
        RECT 54.170 197.820 54.430 198.140 ;
        RECT 54.230 196.440 54.370 197.820 ;
        RECT 54.690 196.440 54.830 200.200 ;
        RECT 55.150 198.560 55.290 201.560 ;
        RECT 55.150 198.480 55.750 198.560 ;
        RECT 55.150 198.420 55.810 198.480 ;
        RECT 55.550 198.160 55.810 198.420 ;
        RECT 55.090 197.820 55.350 198.140 ;
        RECT 55.150 196.440 55.290 197.820 ;
        RECT 54.170 196.120 54.430 196.440 ;
        RECT 54.630 196.120 54.890 196.440 ;
        RECT 55.090 196.120 55.350 196.440 ;
        RECT 53.710 195.780 53.970 196.100 ;
        RECT 50.950 195.440 51.210 195.760 ;
        RECT 52.330 195.440 52.590 195.760 ;
        RECT 50.490 194.420 50.750 194.740 ;
        RECT 51.010 193.380 51.150 195.440 ;
        RECT 50.950 193.060 51.210 193.380 ;
        RECT 52.330 193.060 52.590 193.380 ;
        RECT 46.350 192.380 46.610 192.700 ;
        RECT 45.890 192.040 46.150 192.360 ;
        RECT 44.970 191.700 45.230 192.020 ;
        RECT 44.050 190.680 44.310 191.000 ;
        RECT 43.590 187.280 43.850 187.600 ;
        RECT 43.590 183.540 43.850 183.860 ;
        RECT 43.650 182.160 43.790 183.540 ;
        RECT 43.590 181.840 43.850 182.160 ;
        RECT 43.130 181.500 43.390 181.820 ;
        RECT 43.590 181.160 43.850 181.480 ;
        RECT 40.370 180.820 40.630 181.140 ;
        RECT 41.290 180.820 41.550 181.140 ;
        RECT 39.910 179.800 40.170 180.120 ;
        RECT 40.430 179.440 40.570 180.820 ;
        RECT 40.370 179.120 40.630 179.440 ;
        RECT 38.990 178.100 39.250 178.420 ;
        RECT 39.450 177.080 39.710 177.400 ;
        RECT 38.530 176.740 38.790 177.060 ;
        RECT 36.120 174.845 37.660 175.215 ;
        RECT 35.770 174.360 36.030 174.680 ;
        RECT 39.510 174.000 39.650 177.080 ;
        RECT 39.450 173.680 39.710 174.000 ;
        RECT 40.370 173.680 40.630 174.000 ;
        RECT 35.310 173.340 35.570 173.660 ;
        RECT 39.510 173.400 39.650 173.680 ;
        RECT 34.850 173.000 35.110 173.320 ;
        RECT 39.510 173.260 40.110 173.400 ;
        RECT 32.820 172.125 34.360 172.495 ;
        RECT 32.090 171.640 32.350 171.960 ;
        RECT 32.090 170.280 32.350 170.600 ;
        RECT 32.150 169.240 32.290 170.280 ;
        RECT 34.910 170.260 35.050 173.000 ;
        RECT 38.070 172.660 38.330 172.980 ;
        RECT 39.450 172.660 39.710 172.980 ;
        RECT 34.850 169.940 35.110 170.260 ;
        RECT 36.120 169.405 37.660 169.775 ;
        RECT 32.090 168.920 32.350 169.240 ;
        RECT 36.690 168.240 36.950 168.560 ;
        RECT 21.050 167.220 21.310 167.540 ;
        RECT 31.630 167.220 31.890 167.540 ;
        RECT 32.820 166.685 34.360 167.055 ;
        RECT 36.750 166.520 36.890 168.240 ;
        RECT 36.690 166.200 36.950 166.520 ;
        RECT 38.130 165.160 38.270 172.660 ;
        RECT 38.530 169.940 38.790 170.260 ;
        RECT 38.590 165.160 38.730 169.940 ;
        RECT 39.510 166.520 39.650 172.660 ;
        RECT 39.970 170.940 40.110 173.260 ;
        RECT 40.430 171.960 40.570 173.680 ;
        RECT 40.370 171.640 40.630 171.960 ;
        RECT 40.430 170.940 40.570 171.640 ;
        RECT 39.910 170.620 40.170 170.940 ;
        RECT 40.370 170.620 40.630 170.940 ;
        RECT 39.970 169.240 40.110 170.620 ;
        RECT 41.350 170.600 41.490 180.820 ;
        RECT 43.650 180.120 43.790 181.160 ;
        RECT 43.590 179.800 43.850 180.120 ;
        RECT 43.590 175.720 43.850 176.040 ;
        RECT 43.650 174.680 43.790 175.720 ;
        RECT 41.750 174.360 42.010 174.680 ;
        RECT 43.590 174.360 43.850 174.680 ;
        RECT 41.290 170.280 41.550 170.600 ;
        RECT 39.910 168.920 40.170 169.240 ;
        RECT 39.450 166.200 39.710 166.520 ;
        RECT 38.070 164.840 38.330 165.160 ;
        RECT 38.530 164.840 38.790 165.160 ;
        RECT 36.120 163.965 37.660 164.335 ;
        RECT 32.820 161.245 34.360 161.615 ;
        RECT 35.310 160.760 35.570 161.080 ;
        RECT 32.550 159.740 32.810 160.060 ;
        RECT 16.485 159.340 16.905 159.575 ;
        RECT 15.840 158.400 16.260 158.410 ;
        RECT 16.485 158.400 16.720 159.340 ;
        RECT 15.840 158.060 16.860 158.400 ;
        RECT 15.840 157.960 16.260 158.060 ;
        RECT 32.610 157.680 32.750 159.740 ;
        RECT 33.470 159.400 33.730 159.720 ;
        RECT 29.330 157.360 29.590 157.680 ;
        RECT 32.550 157.360 32.810 157.680 ;
        RECT 29.390 151.900 29.530 157.360 ;
        RECT 32.610 157.080 32.750 157.360 ;
        RECT 33.530 157.340 33.670 159.400 ;
        RECT 33.930 159.060 34.190 159.380 ;
        RECT 33.990 158.020 34.130 159.060 ;
        RECT 35.370 158.270 35.510 160.760 ;
        RECT 35.770 160.420 36.030 160.740 ;
        RECT 34.450 158.130 35.510 158.270 ;
        RECT 33.930 157.700 34.190 158.020 ;
        RECT 32.150 156.940 32.750 157.080 ;
        RECT 33.470 157.020 33.730 157.340 ;
        RECT 34.450 157.000 34.590 158.130 ;
        RECT 34.850 157.360 35.110 157.680 ;
        RECT 32.150 155.640 32.290 156.940 ;
        RECT 34.390 156.680 34.650 157.000 ;
        RECT 32.820 155.805 34.360 156.175 ;
        RECT 32.090 155.320 32.350 155.640 ;
        RECT 34.910 154.620 35.050 157.360 ;
        RECT 34.850 154.300 35.110 154.620 ;
        RECT 29.330 151.580 29.590 151.900 ;
        RECT 29.390 147.480 29.530 151.580 ;
        RECT 32.090 150.900 32.350 151.220 ;
        RECT 32.150 148.840 32.290 150.900 ;
        RECT 32.820 150.365 34.360 150.735 ;
        RECT 34.910 149.520 35.050 154.300 ;
        RECT 35.370 151.900 35.510 158.130 ;
        RECT 35.830 157.680 35.970 160.420 ;
        RECT 38.990 160.080 39.250 160.400 ;
        RECT 38.530 159.740 38.790 160.060 ;
        RECT 38.070 159.400 38.330 159.720 ;
        RECT 36.120 158.525 37.660 158.895 ;
        RECT 35.770 157.360 36.030 157.680 ;
        RECT 36.230 156.340 36.490 156.660 ;
        RECT 36.290 154.280 36.430 156.340 ;
        RECT 38.130 155.300 38.270 159.400 ;
        RECT 38.070 154.980 38.330 155.300 ;
        RECT 36.230 153.960 36.490 154.280 ;
        RECT 35.770 153.620 36.030 153.940 ;
        RECT 35.310 151.580 35.570 151.900 ;
        RECT 35.310 150.900 35.570 151.220 ;
        RECT 34.850 149.200 35.110 149.520 ;
        RECT 32.090 148.520 32.350 148.840 ;
        RECT 34.850 148.520 35.110 148.840 ;
        RECT 29.330 147.160 29.590 147.480 ;
        RECT 22.890 146.480 23.150 146.800 ;
        RECT 19.210 145.460 19.470 145.780 ;
        RECT 19.270 144.275 19.410 145.460 ;
        RECT 19.200 143.905 19.480 144.275 ;
        RECT 20.590 143.420 20.850 143.740 ;
        RECT 15.990 142.740 16.250 143.060 ;
        RECT 16.050 141.555 16.190 142.740 ;
        RECT 15.980 141.185 16.260 141.555 ;
        RECT 18.750 141.040 19.010 141.360 ;
        RECT 18.810 139.320 18.950 141.040 ;
        RECT 19.210 140.700 19.470 141.020 ;
        RECT 18.750 139.000 19.010 139.320 ;
        RECT 16.440 137.105 16.720 137.475 ;
        RECT 16.510 136.260 16.650 137.105 ;
        RECT 16.450 135.940 16.710 136.260 ;
        RECT 15.990 134.755 16.250 134.900 ;
        RECT 15.980 134.385 16.260 134.755 ;
        RECT 19.270 133.280 19.410 140.700 ;
        RECT 20.650 140.340 20.790 143.420 ;
        RECT 22.950 141.700 23.090 146.480 ;
        RECT 32.820 144.925 34.360 145.295 ;
        RECT 34.910 143.400 35.050 148.520 ;
        RECT 35.370 147.480 35.510 150.900 ;
        RECT 35.830 150.200 35.970 153.620 ;
        RECT 36.120 153.085 37.660 153.455 ;
        RECT 38.130 152.920 38.270 154.980 ;
        RECT 38.590 154.620 38.730 159.740 ;
        RECT 39.050 154.620 39.190 160.080 ;
        RECT 41.810 160.060 41.950 174.360 ;
        RECT 44.110 174.000 44.250 190.680 ;
        RECT 44.510 186.940 44.770 187.260 ;
        RECT 44.570 179.100 44.710 186.940 ;
        RECT 45.030 185.220 45.170 191.700 ;
        RECT 46.410 189.640 46.550 192.380 ;
        RECT 47.730 190.000 47.990 190.320 ;
        RECT 46.350 189.320 46.610 189.640 ;
        RECT 47.790 187.260 47.930 190.000 ;
        RECT 47.730 186.940 47.990 187.260 ;
        RECT 45.430 186.260 45.690 186.580 ;
        RECT 44.970 184.900 45.230 185.220 ;
        RECT 45.490 184.880 45.630 186.260 ;
        RECT 45.430 184.560 45.690 184.880 ;
        RECT 45.890 184.560 46.150 184.880 ;
        RECT 45.950 182.840 46.090 184.560 ;
        RECT 45.890 182.520 46.150 182.840 ;
        RECT 48.190 181.500 48.450 181.820 ;
        RECT 48.250 179.440 48.390 181.500 ;
        RECT 48.190 179.120 48.450 179.440 ;
        RECT 44.510 178.780 44.770 179.100 ;
        RECT 45.430 178.780 45.690 179.100 ;
        RECT 46.810 178.780 47.070 179.100 ;
        RECT 48.650 178.780 48.910 179.100 ;
        RECT 50.490 178.780 50.750 179.100 ;
        RECT 44.570 177.400 44.710 178.780 ;
        RECT 44.510 177.080 44.770 177.400 ;
        RECT 45.490 176.720 45.630 178.780 ;
        RECT 45.890 178.100 46.150 178.420 ;
        RECT 45.430 176.400 45.690 176.720 ;
        RECT 44.970 175.380 45.230 175.700 ;
        RECT 45.030 174.000 45.170 175.380 ;
        RECT 45.490 174.680 45.630 176.400 ;
        RECT 45.430 174.360 45.690 174.680 ;
        RECT 45.950 174.000 46.090 178.100 ;
        RECT 46.870 177.060 47.010 178.780 ;
        RECT 48.710 177.400 48.850 178.780 ;
        RECT 47.730 177.080 47.990 177.400 ;
        RECT 48.650 177.080 48.910 177.400 ;
        RECT 46.810 176.740 47.070 177.060 ;
        RECT 47.790 176.380 47.930 177.080 ;
        RECT 50.550 176.380 50.690 178.780 ;
        RECT 47.730 176.060 47.990 176.380 ;
        RECT 50.490 176.060 50.750 176.380 ;
        RECT 47.270 175.380 47.530 175.700 ;
        RECT 47.330 174.000 47.470 175.380 ;
        RECT 44.050 173.680 44.310 174.000 ;
        RECT 44.970 173.680 45.230 174.000 ;
        RECT 45.890 173.680 46.150 174.000 ;
        RECT 46.350 173.680 46.610 174.000 ;
        RECT 47.270 173.680 47.530 174.000 ;
        RECT 43.130 173.340 43.390 173.660 ;
        RECT 43.190 170.600 43.330 173.340 ;
        RECT 45.950 172.040 46.090 173.680 ;
        RECT 46.410 172.980 46.550 173.680 ;
        RECT 47.790 172.980 47.930 176.060 ;
        RECT 46.350 172.660 46.610 172.980 ;
        RECT 47.270 172.660 47.530 172.980 ;
        RECT 47.730 172.660 47.990 172.980 ;
        RECT 45.950 171.900 47.010 172.040 ;
        RECT 47.330 171.960 47.470 172.660 ;
        RECT 43.130 170.280 43.390 170.600 ;
        RECT 43.190 169.240 43.330 170.280 ;
        RECT 46.350 169.940 46.610 170.260 ;
        RECT 43.130 168.920 43.390 169.240 ;
        RECT 46.410 168.560 46.550 169.940 ;
        RECT 46.350 168.240 46.610 168.560 ;
        RECT 41.750 159.970 42.010 160.060 ;
        RECT 41.750 159.830 42.870 159.970 ;
        RECT 41.750 159.740 42.010 159.830 ;
        RECT 39.450 159.400 39.710 159.720 ;
        RECT 39.510 159.120 39.650 159.400 ;
        RECT 39.510 158.980 40.110 159.120 ;
        RECT 39.970 156.660 40.110 158.980 ;
        RECT 39.910 156.340 40.170 156.660 ;
        RECT 39.970 154.620 40.110 156.340 ;
        RECT 42.730 154.620 42.870 159.830 ;
        RECT 46.870 159.720 47.010 171.900 ;
        RECT 47.270 171.640 47.530 171.960 ;
        RECT 47.330 171.280 47.470 171.640 ;
        RECT 47.270 170.960 47.530 171.280 ;
        RECT 47.790 170.940 47.930 172.660 ;
        RECT 50.550 170.940 50.690 176.060 ;
        RECT 47.730 170.620 47.990 170.940 ;
        RECT 50.490 170.620 50.750 170.940 ;
        RECT 47.730 160.760 47.990 161.080 ;
        RECT 46.810 159.400 47.070 159.720 ;
        RECT 46.350 159.060 46.610 159.380 ;
        RECT 47.270 159.060 47.530 159.380 ;
        RECT 46.410 157.680 46.550 159.060 ;
        RECT 47.330 158.020 47.470 159.060 ;
        RECT 47.790 158.020 47.930 160.760 ;
        RECT 50.490 159.060 50.750 159.380 ;
        RECT 47.270 157.700 47.530 158.020 ;
        RECT 47.730 157.700 47.990 158.020 ;
        RECT 46.350 157.360 46.610 157.680 ;
        RECT 46.810 157.360 47.070 157.680 ;
        RECT 46.870 154.620 47.010 157.360 ;
        RECT 47.790 155.300 47.930 157.700 ;
        RECT 50.550 157.680 50.690 159.060 ;
        RECT 50.030 157.360 50.290 157.680 ;
        RECT 50.490 157.360 50.750 157.680 ;
        RECT 50.090 156.660 50.230 157.360 ;
        RECT 51.010 157.340 51.150 193.060 ;
        RECT 51.870 181.160 52.130 181.480 ;
        RECT 51.930 180.120 52.070 181.160 ;
        RECT 51.870 179.800 52.130 180.120 ;
        RECT 52.390 176.720 52.530 193.060 ;
        RECT 54.690 192.360 54.830 196.120 ;
        RECT 55.550 195.440 55.810 195.760 ;
        RECT 55.610 193.380 55.750 195.440 ;
        RECT 56.070 195.080 56.210 202.920 ;
        RECT 58.370 202.900 58.510 208.020 ;
        RECT 59.290 205.960 59.430 208.360 ;
        RECT 59.750 206.640 59.890 208.360 ;
        RECT 59.690 206.320 59.950 206.640 ;
        RECT 59.230 205.640 59.490 205.960 ;
        RECT 58.770 203.600 59.030 203.920 ;
        RECT 58.310 202.580 58.570 202.900 ;
        RECT 58.830 201.200 58.970 203.600 ;
        RECT 58.770 200.880 59.030 201.200 ;
        RECT 59.230 200.880 59.490 201.200 ;
        RECT 57.390 200.770 57.650 200.860 ;
        RECT 56.990 200.630 57.650 200.770 ;
        RECT 56.990 200.180 57.130 200.630 ;
        RECT 57.390 200.540 57.650 200.630 ;
        RECT 56.930 199.860 57.190 200.180 ;
        RECT 57.390 199.860 57.650 200.180 ;
        RECT 57.450 199.160 57.590 199.860 ;
        RECT 57.390 198.840 57.650 199.160 ;
        RECT 57.850 198.500 58.110 198.820 ;
        RECT 57.390 197.820 57.650 198.140 ;
        RECT 56.470 197.140 56.730 197.460 ;
        RECT 56.010 194.760 56.270 195.080 ;
        RECT 55.550 193.060 55.810 193.380 ;
        RECT 56.530 192.700 56.670 197.140 ;
        RECT 57.450 196.350 57.590 197.820 ;
        RECT 56.990 196.210 57.590 196.350 ;
        RECT 56.990 195.760 57.130 196.210 ;
        RECT 56.930 195.440 57.190 195.760 ;
        RECT 57.390 195.440 57.650 195.760 ;
        RECT 56.990 192.700 57.130 195.440 ;
        RECT 57.450 193.040 57.590 195.440 ;
        RECT 57.910 195.080 58.050 198.500 ;
        RECT 59.290 198.140 59.430 200.880 ;
        RECT 59.230 197.820 59.490 198.140 ;
        RECT 59.750 195.760 59.890 206.320 ;
        RECT 61.590 204.600 61.730 208.700 ;
        RECT 62.970 207.320 63.110 209.040 ;
        RECT 64.350 209.020 64.490 213.460 ;
        RECT 64.290 208.700 64.550 209.020 ;
        RECT 62.910 207.000 63.170 207.320 ;
        RECT 65.270 206.640 65.410 216.180 ;
        RECT 65.670 214.140 65.930 214.460 ;
        RECT 65.730 211.740 65.870 214.140 ;
        RECT 68.490 212.760 68.630 217.200 ;
        RECT 68.430 212.440 68.690 212.760 ;
        RECT 66.130 211.760 66.390 212.080 ;
        RECT 65.670 211.420 65.930 211.740 ;
        RECT 65.730 209.360 65.870 211.420 ;
        RECT 65.670 209.040 65.930 209.360 ;
        RECT 66.190 208.340 66.330 211.760 ;
        RECT 68.950 210.040 69.090 217.200 ;
        RECT 69.350 216.180 69.610 216.500 ;
        RECT 69.410 214.120 69.550 216.180 ;
        RECT 69.350 213.800 69.610 214.120 ;
        RECT 69.350 211.760 69.610 212.080 ;
        RECT 69.410 210.040 69.550 211.760 ;
        RECT 68.890 209.720 69.150 210.040 ;
        RECT 69.350 209.720 69.610 210.040 ;
        RECT 67.050 208.360 67.310 208.680 ;
        RECT 66.130 208.020 66.390 208.340 ;
        RECT 65.210 206.320 65.470 206.640 ;
        RECT 61.530 204.280 61.790 204.600 ;
        RECT 60.610 203.940 60.870 204.260 ;
        RECT 60.150 199.860 60.410 200.180 ;
        RECT 60.210 196.100 60.350 199.860 ;
        RECT 60.670 198.480 60.810 203.940 ;
        RECT 61.590 201.200 61.730 204.280 ;
        RECT 62.450 203.260 62.710 203.580 ;
        RECT 61.530 200.880 61.790 201.200 ;
        RECT 61.070 199.860 61.330 200.180 ;
        RECT 60.610 198.160 60.870 198.480 ;
        RECT 61.130 197.880 61.270 199.860 ;
        RECT 60.670 197.740 61.270 197.880 ;
        RECT 60.670 196.440 60.810 197.740 ;
        RECT 61.070 197.140 61.330 197.460 ;
        RECT 61.130 196.440 61.270 197.140 ;
        RECT 60.610 196.120 60.870 196.440 ;
        RECT 61.070 196.120 61.330 196.440 ;
        RECT 60.150 195.780 60.410 196.100 ;
        RECT 59.230 195.440 59.490 195.760 ;
        RECT 59.690 195.440 59.950 195.760 ;
        RECT 61.530 195.440 61.790 195.760 ;
        RECT 57.850 194.760 58.110 195.080 ;
        RECT 57.390 192.720 57.650 193.040 ;
        RECT 56.470 192.380 56.730 192.700 ;
        RECT 56.930 192.380 57.190 192.700 ;
        RECT 54.630 192.040 54.890 192.360 ;
        RECT 54.170 191.700 54.430 192.020 ;
        RECT 52.790 190.000 53.050 190.320 ;
        RECT 52.850 187.600 52.990 190.000 ;
        RECT 54.230 187.940 54.370 191.700 ;
        RECT 57.450 190.320 57.590 192.720 ;
        RECT 55.550 190.000 55.810 190.320 ;
        RECT 57.390 190.000 57.650 190.320 ;
        RECT 54.170 187.620 54.430 187.940 ;
        RECT 52.790 187.280 53.050 187.600 ;
        RECT 52.850 181.820 52.990 187.280 ;
        RECT 53.250 186.600 53.510 186.920 ;
        RECT 52.790 181.500 53.050 181.820 ;
        RECT 53.310 178.420 53.450 186.600 ;
        RECT 53.250 178.100 53.510 178.420 ;
        RECT 55.610 176.720 55.750 190.000 ;
        RECT 57.910 187.940 58.050 194.760 ;
        RECT 59.290 192.020 59.430 195.440 ;
        RECT 61.070 195.100 61.330 195.420 ;
        RECT 61.130 193.020 61.270 195.100 ;
        RECT 61.590 193.720 61.730 195.440 ;
        RECT 61.530 193.400 61.790 193.720 ;
        RECT 61.130 192.880 61.730 193.020 ;
        RECT 60.150 192.380 60.410 192.700 ;
        RECT 59.230 191.700 59.490 192.020 ;
        RECT 60.210 190.660 60.350 192.380 ;
        RECT 61.590 192.020 61.730 192.880 ;
        RECT 61.990 192.380 62.250 192.700 ;
        RECT 61.530 191.700 61.790 192.020 ;
        RECT 60.150 190.340 60.410 190.660 ;
        RECT 59.690 189.660 59.950 189.980 ;
        RECT 58.310 188.980 58.570 189.300 ;
        RECT 57.850 187.620 58.110 187.940 ;
        RECT 58.370 186.920 58.510 188.980 ;
        RECT 59.750 187.260 59.890 189.660 ;
        RECT 60.210 189.300 60.350 190.340 ;
        RECT 60.610 190.000 60.870 190.320 ;
        RECT 60.150 188.980 60.410 189.300 ;
        RECT 60.670 187.260 60.810 190.000 ;
        RECT 61.590 187.260 61.730 191.700 ;
        RECT 62.050 190.320 62.190 192.380 ;
        RECT 61.990 190.000 62.250 190.320 ;
        RECT 62.510 189.720 62.650 203.260 ;
        RECT 66.190 200.860 66.330 208.020 ;
        RECT 67.110 205.960 67.250 208.360 ;
        RECT 68.430 208.020 68.690 208.340 ;
        RECT 68.490 206.980 68.630 208.020 ;
        RECT 68.430 206.660 68.690 206.980 ;
        RECT 68.890 205.980 69.150 206.300 ;
        RECT 67.050 205.640 67.310 205.960 ;
        RECT 67.510 205.300 67.770 205.620 ;
        RECT 67.570 204.600 67.710 205.300 ;
        RECT 67.510 204.280 67.770 204.600 ;
        RECT 68.950 201.200 69.090 205.980 ;
        RECT 66.590 200.880 66.850 201.200 ;
        RECT 68.890 200.880 69.150 201.200 ;
        RECT 62.910 200.540 63.170 200.860 ;
        RECT 66.130 200.540 66.390 200.860 ;
        RECT 62.970 193.040 63.110 200.540 ;
        RECT 65.210 200.200 65.470 200.520 ;
        RECT 63.830 199.860 64.090 200.180 ;
        RECT 63.890 198.820 64.030 199.860 ;
        RECT 63.830 198.500 64.090 198.820 ;
        RECT 65.270 198.140 65.410 200.200 ;
        RECT 65.660 199.665 65.940 200.035 ;
        RECT 65.730 198.140 65.870 199.665 ;
        RECT 66.190 199.160 66.330 200.540 ;
        RECT 66.650 199.160 66.790 200.880 ;
        RECT 67.050 200.540 67.310 200.860 ;
        RECT 66.130 198.840 66.390 199.160 ;
        RECT 66.590 198.840 66.850 199.160 ;
        RECT 67.110 198.480 67.250 200.540 ;
        RECT 67.050 198.160 67.310 198.480 ;
        RECT 65.210 197.820 65.470 198.140 ;
        RECT 65.670 197.820 65.930 198.140 ;
        RECT 67.110 195.080 67.250 198.160 ;
        RECT 68.950 198.140 69.090 200.880 ;
        RECT 69.410 198.820 69.550 209.720 ;
        RECT 70.790 209.700 70.930 217.200 ;
        RECT 82.690 216.860 82.950 217.180 ;
        RECT 71.650 216.180 71.910 216.500 ;
        RECT 71.710 212.080 71.850 216.180 ;
        RECT 82.750 213.780 82.890 216.860 ;
        RECT 80.390 213.460 80.650 213.780 ;
        RECT 82.690 213.460 82.950 213.780 ;
        RECT 80.450 212.080 80.590 213.460 ;
        RECT 71.190 211.760 71.450 212.080 ;
        RECT 71.650 211.760 71.910 212.080 ;
        RECT 80.390 211.760 80.650 212.080 ;
        RECT 81.770 211.760 82.030 212.080 ;
        RECT 71.250 211.480 71.390 211.760 ;
        RECT 71.250 211.340 71.850 211.480 ;
        RECT 70.730 209.380 70.990 209.700 ;
        RECT 70.790 206.640 70.930 209.380 ;
        RECT 71.710 209.020 71.850 211.340 ;
        RECT 71.650 208.700 71.910 209.020 ;
        RECT 70.730 206.320 70.990 206.640 ;
        RECT 69.810 199.860 70.070 200.180 ;
        RECT 69.350 198.500 69.610 198.820 ;
        RECT 69.870 198.140 70.010 199.860 ;
        RECT 68.890 197.820 69.150 198.140 ;
        RECT 69.810 197.820 70.070 198.140 ;
        RECT 71.190 197.480 71.450 197.800 ;
        RECT 69.350 197.140 69.610 197.460 ;
        RECT 69.410 195.760 69.550 197.140 ;
        RECT 71.250 196.440 71.390 197.480 ;
        RECT 71.190 196.120 71.450 196.440 ;
        RECT 69.350 195.440 69.610 195.760 ;
        RECT 67.050 194.760 67.310 195.080 ;
        RECT 63.830 194.420 64.090 194.740 ;
        RECT 69.810 194.420 70.070 194.740 ;
        RECT 62.910 192.720 63.170 193.040 ;
        RECT 63.890 190.660 64.030 194.420 ;
        RECT 69.870 193.380 70.010 194.420 ;
        RECT 69.810 193.060 70.070 193.380 ;
        RECT 69.870 192.700 70.010 193.060 ;
        RECT 69.810 192.380 70.070 192.700 ;
        RECT 71.190 192.380 71.450 192.700 ;
        RECT 66.130 191.700 66.390 192.020 ;
        RECT 65.210 190.680 65.470 191.000 ;
        RECT 63.830 190.340 64.090 190.660 ;
        RECT 65.270 190.320 65.410 190.680 ;
        RECT 65.670 190.340 65.930 190.660 ;
        RECT 63.370 190.000 63.630 190.320 ;
        RECT 65.210 190.000 65.470 190.320 ;
        RECT 62.510 189.580 63.110 189.720 ;
        RECT 62.450 188.980 62.710 189.300 ;
        RECT 62.510 187.260 62.650 188.980 ;
        RECT 62.970 187.940 63.110 189.580 ;
        RECT 63.430 187.940 63.570 190.000 ;
        RECT 62.910 187.620 63.170 187.940 ;
        RECT 63.370 187.620 63.630 187.940 ;
        RECT 59.690 186.940 59.950 187.260 ;
        RECT 60.150 186.940 60.410 187.260 ;
        RECT 60.610 186.940 60.870 187.260 ;
        RECT 61.530 186.940 61.790 187.260 ;
        RECT 62.450 186.940 62.710 187.260 ;
        RECT 58.310 186.600 58.570 186.920 ;
        RECT 60.210 185.560 60.350 186.940 ;
        RECT 60.150 185.240 60.410 185.560 ;
        RECT 60.670 185.220 60.810 186.940 ;
        RECT 61.990 185.240 62.250 185.560 ;
        RECT 60.610 184.900 60.870 185.220 ;
        RECT 62.050 184.880 62.190 185.240 ;
        RECT 62.970 184.960 63.110 187.620 ;
        RECT 63.830 186.940 64.090 187.260 ;
        RECT 63.890 185.560 64.030 186.940 ;
        RECT 63.830 185.240 64.090 185.560 ;
        RECT 62.970 184.880 63.570 184.960 ;
        RECT 61.990 184.560 62.250 184.880 ;
        RECT 62.970 184.820 63.630 184.880 ;
        RECT 63.370 184.560 63.630 184.820 ;
        RECT 65.270 183.600 65.410 190.000 ;
        RECT 64.810 183.460 65.410 183.600 ;
        RECT 58.310 182.180 58.570 182.500 ;
        RECT 56.930 179.800 57.190 180.120 ;
        RECT 56.990 179.100 57.130 179.800 ;
        RECT 58.370 179.440 58.510 182.180 ;
        RECT 61.070 181.160 61.330 181.480 ;
        RECT 58.310 179.120 58.570 179.440 ;
        RECT 61.130 179.100 61.270 181.160 ;
        RECT 63.370 180.820 63.630 181.140 ;
        RECT 63.430 179.100 63.570 180.820 ;
        RECT 56.930 178.780 57.190 179.100 ;
        RECT 61.070 178.780 61.330 179.100 ;
        RECT 63.370 178.780 63.630 179.100 ;
        RECT 52.330 176.400 52.590 176.720 ;
        RECT 55.550 176.400 55.810 176.720 ;
        RECT 52.390 157.680 52.530 176.400 ;
        RECT 54.170 173.680 54.430 174.000 ;
        RECT 54.230 171.960 54.370 173.680 ;
        RECT 55.610 173.660 55.750 176.400 ;
        RECT 56.990 176.380 57.130 178.780 ;
        RECT 58.310 178.100 58.570 178.420 ;
        RECT 58.770 178.100 59.030 178.420 ;
        RECT 56.930 176.060 57.190 176.380 ;
        RECT 58.370 174.340 58.510 178.100 ;
        RECT 58.830 176.380 58.970 178.100 ;
        RECT 58.770 176.060 59.030 176.380 ;
        RECT 58.310 174.020 58.570 174.340 ;
        RECT 55.550 173.340 55.810 173.660 ;
        RECT 54.170 171.640 54.430 171.960 ;
        RECT 55.610 168.900 55.750 173.340 ;
        RECT 55.550 168.580 55.810 168.900 ;
        RECT 62.450 167.220 62.710 167.540 ;
        RECT 56.010 165.860 56.270 166.180 ;
        RECT 56.070 163.120 56.210 165.860 ;
        RECT 57.390 165.180 57.650 165.500 ;
        RECT 57.450 163.800 57.590 165.180 ;
        RECT 61.530 164.840 61.790 165.160 ;
        RECT 57.390 163.480 57.650 163.800 ;
        RECT 57.910 163.120 59.430 163.200 ;
        RECT 56.010 163.030 56.270 163.120 ;
        RECT 57.910 163.060 59.490 163.120 ;
        RECT 56.010 162.890 56.670 163.030 ;
        RECT 56.010 162.800 56.270 162.890 ;
        RECT 56.530 160.740 56.670 162.890 ;
        RECT 57.910 162.440 58.050 163.060 ;
        RECT 59.230 162.800 59.490 163.060 ;
        RECT 58.770 162.460 59.030 162.780 ;
        RECT 57.850 162.120 58.110 162.440 ;
        RECT 56.470 160.420 56.730 160.740 ;
        RECT 58.830 160.480 58.970 162.460 ;
        RECT 60.610 161.780 60.870 162.100 ;
        RECT 60.670 161.080 60.810 161.780 ;
        RECT 60.610 160.760 60.870 161.080 ;
        RECT 55.090 159.740 55.350 160.060 ;
        RECT 56.010 159.740 56.270 160.060 ;
        RECT 56.530 159.800 56.670 160.420 ;
        RECT 58.830 160.400 60.350 160.480 ;
        RECT 58.770 160.340 60.350 160.400 ;
        RECT 58.770 160.080 59.030 160.340 ;
        RECT 54.630 159.060 54.890 159.380 ;
        RECT 54.690 158.020 54.830 159.060 ;
        RECT 52.850 157.680 54.370 157.760 ;
        RECT 54.630 157.700 54.890 158.020 ;
        RECT 51.410 157.360 51.670 157.680 ;
        RECT 52.330 157.360 52.590 157.680 ;
        RECT 52.850 157.620 54.430 157.680 ;
        RECT 50.950 157.020 51.210 157.340 ;
        RECT 50.030 156.340 50.290 156.660 ;
        RECT 51.470 155.640 51.610 157.360 ;
        RECT 52.850 157.340 52.990 157.620 ;
        RECT 54.170 157.360 54.430 157.620 ;
        RECT 52.790 157.020 53.050 157.340 ;
        RECT 51.410 155.320 51.670 155.640 ;
        RECT 47.730 154.980 47.990 155.300 ;
        RECT 38.530 154.300 38.790 154.620 ;
        RECT 38.990 154.300 39.250 154.620 ;
        RECT 39.910 154.300 40.170 154.620 ;
        RECT 40.830 154.300 41.090 154.620 ;
        RECT 42.210 154.300 42.470 154.620 ;
        RECT 42.670 154.300 42.930 154.620 ;
        RECT 46.810 154.300 47.070 154.620 ;
        RECT 38.070 152.600 38.330 152.920 ;
        RECT 38.590 152.240 38.730 154.300 ;
        RECT 39.050 152.920 39.190 154.300 ;
        RECT 38.990 152.600 39.250 152.920 ;
        RECT 38.530 151.920 38.790 152.240 ;
        RECT 39.050 151.900 39.190 152.600 ;
        RECT 39.970 152.580 40.110 154.300 ;
        RECT 40.890 152.920 41.030 154.300 ;
        RECT 42.270 153.940 42.410 154.300 ;
        RECT 42.210 153.620 42.470 153.940 ;
        RECT 45.890 153.620 46.150 153.940 ;
        RECT 40.830 152.600 41.090 152.920 ;
        RECT 39.910 152.260 40.170 152.580 ;
        RECT 38.990 151.580 39.250 151.900 ;
        RECT 38.530 150.900 38.790 151.220 ;
        RECT 35.770 149.880 36.030 150.200 ;
        RECT 35.770 149.200 36.030 149.520 ;
        RECT 35.310 147.160 35.570 147.480 ;
        RECT 35.830 146.800 35.970 149.200 ;
        RECT 38.590 149.180 38.730 150.900 ;
        RECT 40.890 150.200 41.030 152.600 ;
        RECT 40.830 149.880 41.090 150.200 ;
        RECT 38.530 148.860 38.790 149.180 ;
        RECT 36.120 147.645 37.660 148.015 ;
        RECT 35.770 146.480 36.030 146.800 ;
        RECT 35.830 144.080 35.970 146.480 ;
        RECT 38.590 146.460 38.730 148.860 ;
        RECT 44.970 148.520 45.230 148.840 ;
        RECT 39.450 147.160 39.710 147.480 ;
        RECT 42.210 147.160 42.470 147.480 ;
        RECT 39.510 146.800 39.650 147.160 ;
        RECT 42.270 146.800 42.410 147.160 ;
        RECT 45.030 147.140 45.170 148.520 ;
        RECT 44.970 146.820 45.230 147.140 ;
        RECT 39.450 146.480 39.710 146.800 ;
        RECT 42.210 146.480 42.470 146.800 ;
        RECT 42.670 146.480 42.930 146.800 ;
        RECT 38.530 146.140 38.790 146.460 ;
        RECT 41.750 145.800 42.010 146.120 ;
        RECT 36.690 145.460 36.950 145.780 ;
        RECT 39.450 145.460 39.710 145.780 ;
        RECT 36.750 144.720 36.890 145.460 ;
        RECT 39.510 144.760 39.650 145.460 ;
        RECT 36.290 144.580 36.890 144.720 ;
        RECT 35.770 143.760 36.030 144.080 ;
        RECT 34.850 143.080 35.110 143.400 ;
        RECT 22.890 141.380 23.150 141.700 ;
        RECT 20.590 140.020 20.850 140.340 ;
        RECT 20.650 138.300 20.790 140.020 ;
        RECT 22.950 139.320 23.090 141.380 ;
        RECT 35.830 141.360 35.970 143.760 ;
        RECT 36.290 143.400 36.430 144.580 ;
        RECT 39.450 144.440 39.710 144.760 ;
        RECT 36.230 143.080 36.490 143.400 ;
        RECT 38.070 142.740 38.330 143.060 ;
        RECT 36.120 142.205 37.660 142.575 ;
        RECT 38.130 141.700 38.270 142.740 ;
        RECT 38.070 141.380 38.330 141.700 ;
        RECT 27.950 141.040 28.210 141.360 ;
        RECT 35.770 141.040 36.030 141.360 ;
        RECT 28.010 139.320 28.150 141.040 ;
        RECT 41.810 141.020 41.950 145.800 ;
        RECT 42.270 145.780 42.410 146.480 ;
        RECT 42.730 146.120 42.870 146.480 ;
        RECT 42.670 145.800 42.930 146.120 ;
        RECT 45.950 145.780 46.090 153.620 ;
        RECT 46.870 146.460 47.010 154.300 ;
        RECT 52.850 149.520 52.990 157.020 ;
        RECT 55.150 157.000 55.290 159.740 ;
        RECT 56.070 158.020 56.210 159.740 ;
        RECT 56.530 159.720 57.590 159.800 ;
        RECT 56.470 159.660 57.590 159.720 ;
        RECT 56.470 159.400 56.730 159.660 ;
        RECT 56.930 159.060 57.190 159.380 ;
        RECT 56.010 157.700 56.270 158.020 ;
        RECT 56.990 157.680 57.130 159.060 ;
        RECT 56.470 157.360 56.730 157.680 ;
        RECT 56.930 157.360 57.190 157.680 ;
        RECT 55.090 156.680 55.350 157.000 ;
        RECT 54.630 156.340 54.890 156.660 ;
        RECT 54.170 152.260 54.430 152.580 ;
        RECT 53.710 151.920 53.970 152.240 ;
        RECT 53.770 149.860 53.910 151.920 ;
        RECT 53.710 149.540 53.970 149.860 ;
        RECT 52.790 149.200 53.050 149.520 ;
        RECT 50.030 148.860 50.290 149.180 ;
        RECT 50.090 146.800 50.230 148.860 ;
        RECT 50.030 146.480 50.290 146.800 ;
        RECT 46.810 146.140 47.070 146.460 ;
        RECT 42.210 145.460 42.470 145.780 ;
        RECT 45.890 145.460 46.150 145.780 ;
        RECT 42.270 142.040 42.410 145.460 ;
        RECT 46.870 144.760 47.010 146.140 ;
        RECT 49.110 145.460 49.370 145.780 ;
        RECT 49.170 144.760 49.310 145.460 ;
        RECT 44.050 144.440 44.310 144.760 ;
        RECT 46.810 144.440 47.070 144.760 ;
        RECT 49.110 144.440 49.370 144.760 ;
        RECT 44.110 142.040 44.250 144.440 ;
        RECT 50.090 144.420 50.230 146.480 ;
        RECT 52.850 146.460 52.990 149.200 ;
        RECT 54.230 148.920 54.370 152.260 ;
        RECT 54.690 152.240 54.830 156.340 ;
        RECT 54.630 151.920 54.890 152.240 ;
        RECT 55.550 151.920 55.810 152.240 ;
        RECT 54.630 150.900 54.890 151.220 ;
        RECT 53.770 148.780 54.370 148.920 ;
        RECT 52.790 146.140 53.050 146.460 ;
        RECT 48.190 144.160 48.450 144.420 ;
        RECT 47.330 144.100 48.450 144.160 ;
        RECT 50.030 144.100 50.290 144.420 ;
        RECT 47.330 144.020 48.390 144.100 ;
        RECT 47.330 143.740 47.470 144.020 ;
        RECT 52.850 143.740 52.990 146.140 ;
        RECT 53.250 145.460 53.510 145.780 ;
        RECT 53.310 144.760 53.450 145.460 ;
        RECT 53.250 144.440 53.510 144.760 ;
        RECT 47.270 143.420 47.530 143.740 ;
        RECT 52.790 143.420 53.050 143.740 ;
        RECT 44.510 142.740 44.770 143.060 ;
        RECT 42.210 141.720 42.470 142.040 ;
        RECT 44.050 141.720 44.310 142.040 ;
        RECT 44.570 141.360 44.710 142.740 ;
        RECT 52.850 142.040 52.990 143.420 ;
        RECT 53.770 143.400 53.910 148.780 ;
        RECT 54.170 145.460 54.430 145.780 ;
        RECT 53.710 143.080 53.970 143.400 ;
        RECT 52.790 141.720 53.050 142.040 ;
        RECT 54.230 141.700 54.370 145.460 ;
        RECT 54.690 144.760 54.830 150.900 ;
        RECT 55.090 149.200 55.350 149.520 ;
        RECT 55.150 147.480 55.290 149.200 ;
        RECT 55.610 148.500 55.750 151.920 ;
        RECT 56.530 149.860 56.670 157.360 ;
        RECT 57.450 153.940 57.590 159.660 ;
        RECT 58.310 157.360 58.570 157.680 ;
        RECT 58.370 155.300 58.510 157.360 ;
        RECT 58.770 156.340 59.030 156.660 ;
        RECT 58.310 154.980 58.570 155.300 ;
        RECT 57.390 153.620 57.650 153.940 ;
        RECT 56.470 149.540 56.730 149.860 ;
        RECT 55.550 148.180 55.810 148.500 ;
        RECT 55.090 147.160 55.350 147.480 ;
        RECT 55.610 146.800 55.750 148.180 ;
        RECT 57.450 147.140 57.590 153.620 ;
        RECT 58.830 152.580 58.970 156.340 ;
        RECT 58.770 152.260 59.030 152.580 ;
        RECT 60.210 152.240 60.350 160.340 ;
        RECT 60.670 159.380 60.810 160.760 ;
        RECT 61.070 159.400 61.330 159.720 ;
        RECT 60.610 159.060 60.870 159.380 ;
        RECT 61.130 157.680 61.270 159.400 ;
        RECT 61.590 158.020 61.730 164.840 ;
        RECT 61.990 164.500 62.250 164.820 ;
        RECT 62.050 163.460 62.190 164.500 ;
        RECT 62.510 163.800 62.650 167.220 ;
        RECT 62.910 165.520 63.170 165.840 ;
        RECT 62.450 163.480 62.710 163.800 ;
        RECT 61.990 163.140 62.250 163.460 ;
        RECT 61.530 157.700 61.790 158.020 ;
        RECT 62.970 157.680 63.110 165.520 ;
        RECT 64.810 165.500 64.950 183.460 ;
        RECT 65.210 182.520 65.470 182.840 ;
        RECT 65.270 178.420 65.410 182.520 ;
        RECT 65.730 179.100 65.870 190.340 ;
        RECT 66.190 189.980 66.330 191.700 ;
        RECT 71.250 190.400 71.390 192.380 ;
        RECT 71.710 191.000 71.850 208.700 ;
        RECT 72.570 205.640 72.830 205.960 ;
        RECT 72.630 196.100 72.770 205.640 ;
        RECT 80.450 204.260 80.590 211.760 ;
        RECT 81.830 210.040 81.970 211.760 ;
        RECT 81.770 209.720 82.030 210.040 ;
        RECT 82.750 209.020 82.890 213.460 ;
        RECT 82.690 208.700 82.950 209.020 ;
        RECT 80.850 205.300 81.110 205.620 ;
        RECT 80.390 203.940 80.650 204.260 ;
        RECT 79.930 203.260 80.190 203.580 ;
        RECT 79.990 201.880 80.130 203.260 ;
        RECT 79.930 201.560 80.190 201.880 ;
        RECT 80.450 201.540 80.590 203.940 ;
        RECT 80.910 203.580 81.050 205.300 ;
        RECT 81.310 204.280 81.570 204.600 ;
        RECT 81.370 203.920 81.510 204.280 ;
        RECT 81.310 203.600 81.570 203.920 ;
        RECT 80.850 203.260 81.110 203.580 ;
        RECT 82.230 202.920 82.490 203.240 ;
        RECT 78.550 201.220 78.810 201.540 ;
        RECT 80.390 201.220 80.650 201.540 ;
        RECT 75.330 200.540 75.590 200.860 ;
        RECT 73.490 199.860 73.750 200.180 ;
        RECT 72.570 195.780 72.830 196.100 ;
        RECT 71.650 190.680 71.910 191.000 ;
        RECT 72.110 190.680 72.370 191.000 ;
        RECT 70.330 190.320 71.390 190.400 ;
        RECT 66.590 190.000 66.850 190.320 ;
        RECT 70.270 190.260 71.390 190.320 ;
        RECT 70.270 190.000 70.530 190.260 ;
        RECT 66.130 189.660 66.390 189.980 ;
        RECT 66.650 187.600 66.790 190.000 ;
        RECT 71.250 189.300 71.390 190.260 ;
        RECT 72.170 189.980 72.310 190.680 ;
        RECT 72.110 189.660 72.370 189.980 ;
        RECT 72.630 189.720 72.770 195.780 ;
        RECT 73.550 195.760 73.690 199.860 ;
        RECT 75.390 199.160 75.530 200.540 ;
        RECT 75.330 198.840 75.590 199.160 ;
        RECT 78.610 198.140 78.750 201.220 ;
        RECT 82.290 201.200 82.430 202.920 ;
        RECT 82.690 202.580 82.950 202.900 ;
        RECT 82.750 201.200 82.890 202.580 ;
        RECT 80.850 200.880 81.110 201.200 ;
        RECT 82.230 200.880 82.490 201.200 ;
        RECT 82.690 200.880 82.950 201.200 ;
        RECT 78.550 197.820 78.810 198.140 ;
        RECT 78.610 196.440 78.750 197.820 ;
        RECT 78.550 196.120 78.810 196.440 ;
        RECT 73.490 195.440 73.750 195.760 ;
        RECT 73.550 193.380 73.690 195.440 ;
        RECT 73.490 193.060 73.750 193.380 ;
        RECT 73.550 191.000 73.690 193.060 ;
        RECT 80.910 192.360 81.050 200.880 ;
        RECT 84.070 197.140 84.330 197.460 ;
        RECT 84.130 196.100 84.270 197.140 ;
        RECT 84.070 195.780 84.330 196.100 ;
        RECT 82.230 194.420 82.490 194.740 ;
        RECT 81.770 193.060 82.030 193.380 ;
        RECT 81.310 192.720 81.570 193.040 ;
        RECT 80.850 192.040 81.110 192.360 ;
        RECT 73.490 190.680 73.750 191.000 ;
        RECT 72.630 189.640 73.690 189.720 ;
        RECT 73.950 189.660 74.210 189.980 ;
        RECT 72.630 189.580 73.750 189.640 ;
        RECT 73.490 189.320 73.750 189.580 ;
        RECT 70.730 188.980 70.990 189.300 ;
        RECT 71.190 188.980 71.450 189.300 ;
        RECT 72.570 188.980 72.830 189.300 ;
        RECT 66.590 187.280 66.850 187.600 ;
        RECT 70.790 187.260 70.930 188.980 ;
        RECT 72.630 187.600 72.770 188.980 ;
        RECT 72.570 187.280 72.830 187.600 ;
        RECT 70.730 186.940 70.990 187.260 ;
        RECT 66.590 186.600 66.850 186.920 ;
        RECT 66.130 184.900 66.390 185.220 ;
        RECT 66.190 181.480 66.330 184.900 ;
        RECT 66.650 184.880 66.790 186.600 ;
        RECT 72.630 184.880 72.770 187.280 ;
        RECT 73.550 186.920 73.690 189.320 ;
        RECT 73.490 186.600 73.750 186.920 ;
        RECT 66.590 184.560 66.850 184.880 ;
        RECT 72.570 184.560 72.830 184.880 ;
        RECT 66.650 182.840 66.790 184.560 ;
        RECT 66.590 182.520 66.850 182.840 ;
        RECT 72.630 181.820 72.770 184.560 ;
        RECT 73.030 184.220 73.290 184.540 ;
        RECT 73.090 182.840 73.230 184.220 ;
        RECT 73.030 182.520 73.290 182.840 ;
        RECT 66.590 181.500 66.850 181.820 ;
        RECT 68.430 181.500 68.690 181.820 ;
        RECT 72.570 181.500 72.830 181.820 ;
        RECT 66.130 181.160 66.390 181.480 ;
        RECT 66.190 179.780 66.330 181.160 ;
        RECT 66.130 179.460 66.390 179.780 ;
        RECT 65.670 178.780 65.930 179.100 ;
        RECT 65.210 178.100 65.470 178.420 ;
        RECT 65.270 174.680 65.410 178.100 ;
        RECT 65.730 177.400 65.870 178.780 ;
        RECT 65.670 177.080 65.930 177.400 ;
        RECT 66.190 177.060 66.330 179.460 ;
        RECT 66.650 179.440 66.790 181.500 ;
        RECT 67.970 181.160 68.230 181.480 ;
        RECT 67.510 180.820 67.770 181.140 ;
        RECT 67.570 180.120 67.710 180.820 ;
        RECT 68.030 180.120 68.170 181.160 ;
        RECT 67.510 179.800 67.770 180.120 ;
        RECT 67.970 179.800 68.230 180.120 ;
        RECT 66.590 179.120 66.850 179.440 ;
        RECT 68.490 178.760 68.630 181.500 ;
        RECT 68.890 180.820 69.150 181.140 ;
        RECT 68.430 178.440 68.690 178.760 ;
        RECT 66.130 176.740 66.390 177.060 ;
        RECT 68.950 176.380 69.090 180.820 ;
        RECT 73.550 179.780 73.690 186.600 ;
        RECT 74.010 186.580 74.150 189.660 ;
        RECT 80.910 188.280 81.050 192.040 ;
        RECT 81.370 189.980 81.510 192.720 ;
        RECT 81.830 191.000 81.970 193.060 ;
        RECT 81.770 190.680 82.030 191.000 ;
        RECT 82.290 190.660 82.430 194.420 ;
        RECT 84.590 193.020 84.730 219.240 ;
        RECT 85.450 218.900 85.710 219.220 ;
        RECT 85.510 214.120 85.650 218.900 ;
        RECT 85.910 216.860 86.170 217.180 ;
        RECT 85.450 213.800 85.710 214.120 ;
        RECT 85.970 212.760 86.110 216.860 ;
        RECT 87.350 212.760 87.490 219.580 ;
        RECT 85.910 212.440 86.170 212.760 ;
        RECT 87.290 212.440 87.550 212.760 ;
        RECT 86.370 212.100 86.630 212.420 ;
        RECT 86.430 210.040 86.570 212.100 ;
        RECT 86.370 209.720 86.630 210.040 ;
        RECT 86.430 209.020 86.570 209.720 ;
        RECT 86.370 208.700 86.630 209.020 ;
        RECT 85.910 208.020 86.170 208.340 ;
        RECT 84.990 205.300 85.250 205.620 ;
        RECT 85.050 198.140 85.190 205.300 ;
        RECT 85.970 204.600 86.110 208.020 ;
        RECT 85.910 204.280 86.170 204.600 ;
        RECT 85.910 202.920 86.170 203.240 ;
        RECT 85.970 201.880 86.110 202.920 ;
        RECT 85.910 201.560 86.170 201.880 ;
        RECT 84.990 197.820 85.250 198.140 ;
        RECT 85.910 197.140 86.170 197.460 ;
        RECT 85.970 196.440 86.110 197.140 ;
        RECT 85.910 196.120 86.170 196.440 ;
        RECT 84.590 192.880 85.190 193.020 ;
        RECT 82.230 190.340 82.490 190.660 ;
        RECT 81.310 189.660 81.570 189.980 ;
        RECT 80.850 187.960 81.110 188.280 ;
        RECT 81.370 187.260 81.510 189.660 ;
        RECT 81.310 186.940 81.570 187.260 ;
        RECT 73.950 186.260 74.210 186.580 ;
        RECT 78.090 183.540 78.350 183.860 ;
        RECT 74.410 181.160 74.670 181.480 ;
        RECT 73.490 179.460 73.750 179.780 ;
        RECT 74.470 178.760 74.610 181.160 ;
        RECT 78.150 180.120 78.290 183.540 ;
        RECT 83.610 181.500 83.870 181.820 ;
        RECT 78.090 179.800 78.350 180.120 ;
        RECT 83.670 179.780 83.810 181.500 ;
        RECT 83.610 179.460 83.870 179.780 ;
        RECT 78.090 179.120 78.350 179.440 ;
        RECT 74.410 178.440 74.670 178.760 ;
        RECT 68.890 176.060 69.150 176.380 ;
        RECT 78.150 175.700 78.290 179.120 ;
        RECT 83.670 176.720 83.810 179.460 ;
        RECT 84.530 178.100 84.790 178.420 ;
        RECT 83.610 176.400 83.870 176.720 ;
        RECT 78.090 175.380 78.350 175.700 ;
        RECT 65.210 174.360 65.470 174.680 ;
        RECT 83.150 173.910 83.410 174.000 ;
        RECT 82.750 173.770 83.410 173.910 ;
        RECT 82.750 170.940 82.890 173.770 ;
        RECT 83.150 173.680 83.410 173.770 ;
        RECT 83.670 173.660 83.810 176.400 ;
        RECT 83.610 173.340 83.870 173.660 ;
        RECT 83.670 171.280 83.810 173.340 ;
        RECT 84.590 171.960 84.730 178.100 ;
        RECT 85.050 176.720 85.190 192.880 ;
        RECT 86.830 192.040 87.090 192.360 ;
        RECT 85.910 188.980 86.170 189.300 ;
        RECT 85.970 186.920 86.110 188.980 ;
        RECT 85.910 186.600 86.170 186.920 ;
        RECT 86.370 186.600 86.630 186.920 ;
        RECT 86.430 184.540 86.570 186.600 ;
        RECT 86.370 184.220 86.630 184.540 ;
        RECT 86.430 181.820 86.570 184.220 ;
        RECT 86.370 181.500 86.630 181.820 ;
        RECT 84.990 176.400 85.250 176.720 ;
        RECT 85.050 172.980 85.190 176.400 ;
        RECT 85.910 173.340 86.170 173.660 ;
        RECT 84.990 172.660 85.250 172.980 ;
        RECT 84.530 171.640 84.790 171.960 ;
        RECT 85.970 171.620 86.110 173.340 ;
        RECT 85.910 171.300 86.170 171.620 ;
        RECT 83.610 170.960 83.870 171.280 ;
        RECT 82.690 170.620 82.950 170.940 ;
        RECT 84.070 170.620 84.330 170.940 ;
        RECT 82.750 168.900 82.890 170.620 ;
        RECT 82.690 168.580 82.950 168.900 ;
        RECT 84.130 168.560 84.270 170.620 ;
        RECT 86.890 170.600 87.030 192.040 ;
        RECT 87.290 175.380 87.550 175.700 ;
        RECT 87.350 174.340 87.490 175.380 ;
        RECT 87.810 174.340 87.950 220.260 ;
        RECT 89.130 219.580 89.390 219.900 ;
        RECT 103.390 219.580 103.650 219.900 ;
        RECT 88.210 218.900 88.470 219.220 ;
        RECT 87.290 174.020 87.550 174.340 ;
        RECT 87.750 174.020 88.010 174.340 ;
        RECT 87.810 171.620 87.950 174.020 ;
        RECT 88.270 174.000 88.410 218.900 ;
        RECT 89.190 218.200 89.330 219.580 ;
        RECT 89.590 219.240 89.850 219.560 ;
        RECT 89.650 218.200 89.790 219.240 ;
        RECT 90.970 218.900 91.230 219.220 ;
        RECT 89.130 217.880 89.390 218.200 ;
        RECT 89.590 217.880 89.850 218.200 ;
        RECT 90.510 217.540 90.770 217.860 ;
        RECT 89.590 215.160 89.850 215.480 ;
        RECT 89.650 212.080 89.790 215.160 ;
        RECT 90.570 212.080 90.710 217.540 ;
        RECT 91.030 212.080 91.170 218.900 ;
        RECT 93.270 217.880 93.530 218.200 ;
        RECT 93.330 217.520 93.470 217.880 ;
        RECT 103.450 217.860 103.590 219.580 ;
        RECT 95.570 217.540 95.830 217.860 ;
        RECT 97.410 217.540 97.670 217.860 ;
        RECT 103.390 217.540 103.650 217.860 ;
        RECT 93.270 217.200 93.530 217.520 ;
        RECT 93.330 216.500 93.470 217.200 ;
        RECT 93.270 216.180 93.530 216.500 ;
        RECT 91.890 213.800 92.150 214.120 ;
        RECT 91.950 212.760 92.090 213.800 ;
        RECT 91.890 212.440 92.150 212.760 ;
        RECT 89.590 211.760 89.850 212.080 ;
        RECT 90.510 211.760 90.770 212.080 ;
        RECT 90.970 211.760 91.230 212.080 ;
        RECT 92.350 211.760 92.610 212.080 ;
        RECT 89.130 210.740 89.390 211.060 ;
        RECT 89.190 209.020 89.330 210.740 ;
        RECT 89.130 208.700 89.390 209.020 ;
        RECT 89.190 206.640 89.330 208.700 ;
        RECT 89.650 206.980 89.790 211.760 ;
        RECT 90.570 211.060 90.710 211.760 ;
        RECT 90.510 210.740 90.770 211.060 ;
        RECT 90.570 209.020 90.710 210.740 ;
        RECT 91.030 210.040 91.170 211.760 ;
        RECT 90.970 209.720 91.230 210.040 ;
        RECT 92.410 209.700 92.550 211.760 ;
        RECT 95.630 211.740 95.770 217.540 ;
        RECT 96.490 217.200 96.750 217.520 ;
        RECT 96.550 216.840 96.690 217.200 ;
        RECT 96.490 216.750 96.750 216.840 ;
        RECT 96.490 216.610 97.150 216.750 ;
        RECT 96.490 216.520 96.750 216.610 ;
        RECT 96.490 214.140 96.750 214.460 ;
        RECT 96.550 212.420 96.690 214.140 ;
        RECT 97.010 213.780 97.150 216.610 ;
        RECT 97.470 215.480 97.610 217.540 ;
        RECT 98.790 216.860 99.050 217.180 ;
        RECT 97.410 215.160 97.670 215.480 ;
        RECT 96.950 213.460 97.210 213.780 ;
        RECT 96.490 212.100 96.750 212.420 ;
        RECT 95.570 211.420 95.830 211.740 ;
        RECT 93.270 211.310 93.530 211.400 ;
        RECT 92.870 211.170 93.530 211.310 ;
        RECT 92.350 209.380 92.610 209.700 ;
        RECT 92.870 209.020 93.010 211.170 ;
        RECT 93.270 211.080 93.530 211.170 ;
        RECT 90.510 208.700 90.770 209.020 ;
        RECT 92.810 208.700 93.070 209.020 ;
        RECT 95.570 208.020 95.830 208.340 ;
        RECT 89.590 206.660 89.850 206.980 ;
        RECT 89.130 206.320 89.390 206.640 ;
        RECT 89.650 201.540 89.790 206.660 ;
        RECT 94.190 206.320 94.450 206.640 ;
        RECT 91.430 205.300 91.690 205.620 ;
        RECT 91.490 203.580 91.630 205.300 ;
        RECT 91.430 203.260 91.690 203.580 ;
        RECT 89.590 201.220 89.850 201.540 ;
        RECT 89.130 198.050 89.390 198.140 ;
        RECT 89.650 198.050 89.790 201.220 ;
        RECT 91.490 199.160 91.630 203.260 ;
        RECT 94.250 202.900 94.390 206.320 ;
        RECT 94.650 205.300 94.910 205.620 ;
        RECT 94.190 202.580 94.450 202.900 ;
        RECT 94.250 201.880 94.390 202.580 ;
        RECT 94.190 201.560 94.450 201.880 ;
        RECT 94.710 201.200 94.850 205.300 ;
        RECT 95.630 204.600 95.770 208.020 ;
        RECT 96.030 206.320 96.290 206.640 ;
        RECT 96.090 204.600 96.230 206.320 ;
        RECT 95.570 204.280 95.830 204.600 ;
        RECT 96.030 204.280 96.290 204.600 ;
        RECT 95.630 201.880 95.770 204.280 ;
        RECT 96.550 203.920 96.690 212.100 ;
        RECT 97.010 211.060 97.150 213.460 ;
        RECT 98.850 212.080 98.990 216.860 ;
        RECT 103.450 215.480 103.590 217.540 ;
        RECT 106.610 216.520 106.870 216.840 ;
        RECT 104.310 216.180 104.570 216.500 ;
        RECT 103.390 215.160 103.650 215.480 ;
        RECT 100.630 213.800 100.890 214.120 ;
        RECT 103.390 213.800 103.650 214.120 ;
        RECT 97.410 211.760 97.670 212.080 ;
        RECT 98.790 211.760 99.050 212.080 ;
        RECT 96.950 210.740 97.210 211.060 ;
        RECT 96.490 203.600 96.750 203.920 ;
        RECT 95.570 201.560 95.830 201.880 ;
        RECT 95.630 201.280 95.770 201.560 ;
        RECT 92.350 200.880 92.610 201.200 ;
        RECT 94.650 200.880 94.910 201.200 ;
        RECT 95.630 201.140 96.230 201.280 ;
        RECT 92.410 199.160 92.550 200.880 ;
        RECT 94.710 200.600 94.850 200.880 ;
        RECT 94.250 200.460 94.850 200.600 ;
        RECT 91.430 198.840 91.690 199.160 ;
        RECT 92.350 198.840 92.610 199.160 ;
        RECT 90.500 198.305 90.780 198.675 ;
        RECT 90.570 198.140 90.710 198.305 ;
        RECT 94.250 198.140 94.390 200.460 ;
        RECT 94.650 199.860 94.910 200.180 ;
        RECT 94.710 198.820 94.850 199.860 ;
        RECT 94.650 198.500 94.910 198.820 ;
        RECT 96.090 198.480 96.230 201.140 ;
        RECT 96.030 198.160 96.290 198.480 ;
        RECT 89.130 197.910 89.790 198.050 ;
        RECT 89.130 197.820 89.390 197.910 ;
        RECT 90.510 197.820 90.770 198.140 ;
        RECT 94.190 197.820 94.450 198.140 ;
        RECT 95.570 197.820 95.830 198.140 ;
        RECT 90.570 196.440 90.710 197.820 ;
        RECT 94.250 197.460 94.390 197.820 ;
        RECT 94.190 197.140 94.450 197.460 ;
        RECT 94.650 197.140 94.910 197.460 ;
        RECT 90.510 196.120 90.770 196.440 ;
        RECT 94.190 192.380 94.450 192.700 ;
        RECT 90.970 191.700 91.230 192.020 ;
        RECT 91.030 191.000 91.170 191.700 ;
        RECT 90.970 190.680 91.230 191.000 ;
        RECT 94.250 190.400 94.390 192.380 ;
        RECT 94.710 191.000 94.850 197.140 ;
        RECT 95.630 192.700 95.770 197.820 ;
        RECT 96.020 197.625 96.300 197.995 ;
        RECT 96.090 197.460 96.230 197.625 ;
        RECT 96.030 197.140 96.290 197.460 ;
        RECT 96.550 193.720 96.690 203.600 ;
        RECT 96.950 201.395 97.210 201.540 ;
        RECT 96.940 201.025 97.220 201.395 ;
        RECT 96.490 193.400 96.750 193.720 ;
        RECT 95.570 192.380 95.830 192.700 ;
        RECT 94.650 190.680 94.910 191.000 ;
        RECT 94.250 190.260 94.850 190.400 ;
        RECT 94.710 187.940 94.850 190.260 ;
        RECT 96.490 190.000 96.750 190.320 ;
        RECT 96.950 190.000 97.210 190.320 ;
        RECT 94.650 187.620 94.910 187.940 ;
        RECT 94.650 184.560 94.910 184.880 ;
        RECT 94.710 180.120 94.850 184.560 ;
        RECT 95.110 184.220 95.370 184.540 ;
        RECT 94.650 179.800 94.910 180.120 ;
        RECT 95.170 177.400 95.310 184.220 ;
        RECT 96.030 183.540 96.290 183.860 ;
        RECT 96.090 182.160 96.230 183.540 ;
        RECT 96.030 181.840 96.290 182.160 ;
        RECT 95.570 180.820 95.830 181.140 ;
        RECT 96.030 180.820 96.290 181.140 ;
        RECT 95.110 177.080 95.370 177.400 ;
        RECT 90.970 174.020 91.230 174.340 ;
        RECT 88.210 173.680 88.470 174.000 ;
        RECT 87.750 171.360 88.010 171.620 ;
        RECT 87.350 171.300 88.010 171.360 ;
        RECT 87.350 171.220 87.950 171.300 ;
        RECT 87.350 170.940 87.490 171.220 ;
        RECT 88.270 170.940 88.410 173.680 ;
        RECT 88.670 173.000 88.930 173.320 ;
        RECT 88.730 171.960 88.870 173.000 ;
        RECT 88.670 171.640 88.930 171.960 ;
        RECT 89.590 171.300 89.850 171.620 ;
        RECT 89.650 170.940 89.790 171.300 ;
        RECT 87.290 170.620 87.550 170.940 ;
        RECT 88.210 170.850 88.470 170.940 ;
        RECT 87.810 170.710 88.470 170.850 ;
        RECT 86.830 170.280 87.090 170.600 ;
        RECT 84.070 168.240 84.330 168.560 ;
        RECT 67.050 167.900 67.310 168.220 ;
        RECT 79.470 167.900 79.730 168.220 ;
        RECT 63.370 165.180 63.630 165.500 ;
        RECT 64.750 165.180 65.010 165.500 ;
        RECT 63.430 161.080 63.570 165.180 ;
        RECT 64.810 164.820 64.950 165.180 ;
        RECT 67.110 165.160 67.250 167.900 ;
        RECT 79.530 166.520 79.670 167.900 ;
        RECT 82.690 167.220 82.950 167.540 ;
        RECT 82.750 166.520 82.890 167.220 ;
        RECT 79.470 166.200 79.730 166.520 ;
        RECT 82.690 166.430 82.950 166.520 ;
        RECT 82.290 166.290 82.950 166.430 ;
        RECT 71.650 165.520 71.910 165.840 ;
        RECT 67.510 165.180 67.770 165.500 ;
        RECT 67.050 164.840 67.310 165.160 ;
        RECT 64.750 164.500 65.010 164.820 ;
        RECT 63.370 160.760 63.630 161.080 ;
        RECT 64.810 160.060 64.950 164.500 ;
        RECT 67.110 162.100 67.250 164.840 ;
        RECT 67.570 162.440 67.710 165.180 ;
        RECT 69.350 164.840 69.610 165.160 ;
        RECT 68.890 162.460 69.150 162.780 ;
        RECT 67.510 162.120 67.770 162.440 ;
        RECT 67.050 161.780 67.310 162.100 ;
        RECT 65.210 160.760 65.470 161.080 ;
        RECT 64.290 159.740 64.550 160.060 ;
        RECT 64.750 159.740 65.010 160.060 ;
        RECT 64.350 158.020 64.490 159.740 ;
        RECT 64.290 157.700 64.550 158.020 ;
        RECT 60.610 157.360 60.870 157.680 ;
        RECT 61.070 157.360 61.330 157.680 ;
        RECT 62.910 157.360 63.170 157.680 ;
        RECT 60.670 157.000 60.810 157.360 ;
        RECT 64.810 157.340 64.950 159.740 ;
        RECT 65.270 158.020 65.410 160.760 ;
        RECT 66.590 159.400 66.850 159.720 ;
        RECT 66.650 158.020 66.790 159.400 ;
        RECT 65.210 157.700 65.470 158.020 ;
        RECT 66.590 157.700 66.850 158.020 ;
        RECT 64.750 157.020 65.010 157.340 ;
        RECT 60.610 156.680 60.870 157.000 ;
        RECT 66.650 155.300 66.790 157.700 ;
        RECT 67.570 157.000 67.710 162.120 ;
        RECT 67.970 161.780 68.230 162.100 ;
        RECT 68.030 160.060 68.170 161.780 ;
        RECT 67.970 159.740 68.230 160.060 ;
        RECT 68.430 159.740 68.690 160.060 ;
        RECT 67.510 156.680 67.770 157.000 ;
        RECT 66.590 154.980 66.850 155.300 ;
        RECT 60.610 154.640 60.870 154.960 ;
        RECT 60.670 152.580 60.810 154.640 ;
        RECT 64.750 153.960 65.010 154.280 ;
        RECT 62.450 153.620 62.710 153.940 ;
        RECT 61.070 152.600 61.330 152.920 ;
        RECT 60.610 152.260 60.870 152.580 ;
        RECT 60.150 151.920 60.410 152.240 ;
        RECT 58.310 150.900 58.570 151.220 ;
        RECT 58.370 150.200 58.510 150.900 ;
        RECT 58.310 149.880 58.570 150.200 ;
        RECT 60.210 149.520 60.350 151.920 ;
        RECT 60.150 149.200 60.410 149.520 ;
        RECT 61.130 147.140 61.270 152.600 ;
        RECT 62.510 152.580 62.650 153.620 ;
        RECT 62.450 152.260 62.710 152.580 ;
        RECT 64.810 150.200 64.950 153.960 ;
        RECT 68.490 153.940 68.630 159.740 ;
        RECT 68.430 153.620 68.690 153.940 ;
        RECT 68.490 152.920 68.630 153.620 ;
        RECT 68.430 152.600 68.690 152.920 ;
        RECT 64.750 149.880 65.010 150.200 ;
        RECT 66.130 149.540 66.390 149.860 ;
        RECT 62.450 149.200 62.710 149.520 ;
        RECT 57.390 146.820 57.650 147.140 ;
        RECT 61.070 146.820 61.330 147.140 ;
        RECT 62.510 146.800 62.650 149.200 ;
        RECT 62.910 148.860 63.170 149.180 ;
        RECT 62.970 147.140 63.110 148.860 ;
        RECT 64.750 148.180 65.010 148.500 ;
        RECT 64.810 147.140 64.950 148.180 ;
        RECT 66.190 147.480 66.330 149.540 ;
        RECT 68.950 149.520 69.090 162.460 ;
        RECT 69.410 156.660 69.550 164.840 ;
        RECT 70.730 162.800 70.990 163.120 ;
        RECT 70.790 161.080 70.930 162.800 ;
        RECT 71.710 162.780 71.850 165.520 ;
        RECT 73.030 164.840 73.290 165.160 ;
        RECT 73.950 164.840 74.210 165.160 ;
        RECT 74.870 164.840 75.130 165.160 ;
        RECT 80.390 164.840 80.650 165.160 ;
        RECT 73.090 163.800 73.230 164.840 ;
        RECT 73.030 163.480 73.290 163.800 ;
        RECT 71.650 162.460 71.910 162.780 ;
        RECT 73.490 162.460 73.750 162.780 ;
        RECT 71.650 161.780 71.910 162.100 ;
        RECT 70.730 160.760 70.990 161.080 ;
        RECT 70.270 160.080 70.530 160.400 ;
        RECT 70.330 157.680 70.470 160.080 ;
        RECT 71.710 158.020 71.850 161.780 ;
        RECT 73.550 160.400 73.690 162.460 ;
        RECT 73.490 160.080 73.750 160.400 ;
        RECT 74.010 160.060 74.150 164.840 ;
        RECT 74.930 162.440 75.070 164.840 ;
        RECT 79.010 164.500 79.270 164.820 ;
        RECT 79.070 163.460 79.210 164.500 ;
        RECT 79.010 163.140 79.270 163.460 ;
        RECT 74.870 162.120 75.130 162.440 ;
        RECT 73.950 159.740 74.210 160.060 ;
        RECT 74.010 158.440 74.150 159.740 ;
        RECT 74.010 158.360 74.610 158.440 ;
        RECT 74.010 158.300 74.670 158.360 ;
        RECT 74.410 158.040 74.670 158.300 ;
        RECT 71.650 157.700 71.910 158.020 ;
        RECT 70.270 157.360 70.530 157.680 ;
        RECT 69.350 156.340 69.610 156.660 ;
        RECT 68.890 149.200 69.150 149.520 ;
        RECT 66.590 148.520 66.850 148.840 ;
        RECT 66.130 147.160 66.390 147.480 ;
        RECT 62.910 146.880 63.170 147.140 ;
        RECT 62.910 146.820 63.570 146.880 ;
        RECT 64.750 146.820 65.010 147.140 ;
        RECT 55.550 146.480 55.810 146.800 ;
        RECT 62.450 146.480 62.710 146.800 ;
        RECT 62.970 146.740 63.570 146.820 ;
        RECT 54.630 144.440 54.890 144.760 ;
        RECT 62.510 143.740 62.650 146.480 ;
        RECT 62.910 145.460 63.170 145.780 ;
        RECT 62.970 144.760 63.110 145.460 ;
        RECT 63.430 144.760 63.570 146.740 ;
        RECT 62.910 144.440 63.170 144.760 ;
        RECT 63.370 144.440 63.630 144.760 ;
        RECT 62.450 143.420 62.710 143.740 ;
        RECT 54.170 141.380 54.430 141.700 ;
        RECT 66.650 141.360 66.790 148.520 ;
        RECT 68.950 146.800 69.090 149.200 ;
        RECT 70.330 149.180 70.470 157.360 ;
        RECT 73.950 154.300 74.210 154.620 ;
        RECT 74.010 152.240 74.150 154.300 ;
        RECT 74.930 153.940 75.070 162.120 ;
        RECT 75.790 161.780 76.050 162.100 ;
        RECT 75.850 160.060 75.990 161.780 ;
        RECT 75.790 159.740 76.050 160.060 ;
        RECT 79.070 159.720 79.210 163.140 ;
        RECT 80.450 162.690 80.590 164.840 ;
        RECT 80.850 162.690 81.110 162.780 ;
        RECT 80.450 162.550 81.110 162.690 ;
        RECT 80.850 162.460 81.110 162.550 ;
        RECT 82.290 160.060 82.430 166.290 ;
        RECT 82.690 166.200 82.950 166.290 ;
        RECT 82.690 164.840 82.950 165.160 ;
        RECT 82.750 163.800 82.890 164.840 ;
        RECT 82.690 163.480 82.950 163.800 ;
        RECT 85.450 162.800 85.710 163.120 ;
        RECT 83.150 161.780 83.410 162.100 ;
        RECT 83.210 160.060 83.350 161.780 ;
        RECT 85.510 161.080 85.650 162.800 ;
        RECT 86.370 162.460 86.630 162.780 ;
        RECT 85.450 160.760 85.710 161.080 ;
        RECT 86.430 160.060 86.570 162.460 ;
        RECT 82.230 159.740 82.490 160.060 ;
        RECT 83.150 159.740 83.410 160.060 ;
        RECT 86.370 159.740 86.630 160.060 ;
        RECT 79.010 159.400 79.270 159.720 ;
        RECT 78.550 159.060 78.810 159.380 ;
        RECT 74.870 153.620 75.130 153.940 ;
        RECT 76.250 153.620 76.510 153.940 ;
        RECT 73.950 151.920 74.210 152.240 ;
        RECT 75.330 151.580 75.590 151.900 ;
        RECT 73.490 150.900 73.750 151.220 ;
        RECT 70.270 148.860 70.530 149.180 ;
        RECT 68.890 146.480 69.150 146.800 ;
        RECT 44.510 141.040 44.770 141.360 ;
        RECT 66.590 141.040 66.850 141.360 ;
        RECT 41.750 140.700 42.010 141.020 ;
        RECT 31.170 140.020 31.430 140.340 ;
        RECT 22.890 139.000 23.150 139.320 ;
        RECT 27.950 139.000 28.210 139.320 ;
        RECT 31.230 138.640 31.370 140.020 ;
        RECT 32.820 139.485 34.360 139.855 ;
        RECT 31.630 139.000 31.890 139.320 ;
        RECT 31.690 138.720 31.830 139.000 ;
        RECT 31.170 138.320 31.430 138.640 ;
        RECT 31.690 138.580 32.290 138.720 ;
        RECT 32.550 138.660 32.810 138.980 ;
        RECT 20.590 137.980 20.850 138.300 ;
        RECT 24.730 137.980 24.990 138.300 ;
        RECT 30.250 137.980 30.510 138.300 ;
        RECT 24.270 137.640 24.530 137.960 ;
        RECT 21.050 135.260 21.310 135.580 ;
        RECT 19.270 133.140 19.870 133.280 ;
        RECT 19.730 132.860 19.870 133.140 ;
        RECT 19.670 132.600 19.930 132.860 ;
        RECT 21.110 132.600 21.250 135.260 ;
        RECT 19.670 132.540 21.250 132.600 ;
        RECT 19.730 132.460 21.250 132.540 ;
        RECT 15.350 131.945 17.000 132.210 ;
        RECT 14.575 131.100 15.140 131.415 ;
        RECT 13.735 130.295 14.315 130.565 ;
        RECT 13.090 129.210 13.550 129.350 ;
        RECT 13.410 120.510 13.550 129.210 ;
        RECT 14.045 121.515 14.315 130.295 ;
        RECT 14.825 122.725 15.140 131.100 ;
        RECT 15.980 129.625 16.260 129.995 ;
        RECT 15.990 129.480 16.250 129.625 ;
        RECT 15.990 127.955 16.250 128.100 ;
        RECT 15.980 127.585 16.260 127.955 ;
        RECT 15.480 123.380 16.180 123.980 ;
        RECT 14.825 122.410 15.460 122.725 ;
        RECT 14.045 121.245 14.795 121.515 ;
        RECT 13.410 120.370 13.890 120.510 ;
        RECT 12.295 117.210 12.585 119.425 ;
        RECT 12.100 116.560 12.780 117.210 ;
        RECT 11.850 94.120 12.110 94.440 ;
        RECT 11.910 86.550 12.050 94.120 ;
        RECT 13.750 92.980 13.890 120.370 ;
        RECT 14.525 110.490 14.795 121.245 ;
        RECT 15.145 112.065 15.460 122.410 ;
        RECT 15.980 119.425 16.260 119.795 ;
        RECT 15.990 119.280 16.250 119.425 ;
        RECT 15.990 112.995 16.250 113.140 ;
        RECT 15.980 112.625 16.260 112.995 ;
        RECT 15.145 111.750 16.450 112.065 ;
        RECT 14.525 110.390 15.750 110.490 ;
        RECT 14.360 109.790 15.750 110.390 ;
        RECT 14.700 109.720 15.750 109.790 ;
        RECT 16.095 107.045 16.450 111.750 ;
        RECT 15.225 107.010 16.465 107.045 ;
        RECT 15.015 106.990 16.465 107.010 ;
        RECT 14.990 106.695 16.465 106.990 ;
        RECT 14.990 106.515 16.445 106.695 ;
        RECT 14.990 106.390 15.990 106.515 ;
        RECT 15.015 106.370 15.565 106.390 ;
        RECT 16.735 103.690 17.000 131.945 ;
        RECT 20.190 125.040 20.330 132.460 ;
        RECT 21.970 132.200 22.230 132.520 ;
        RECT 22.030 131.160 22.170 132.200 ;
        RECT 21.970 130.840 22.230 131.160 ;
        RECT 24.330 130.480 24.470 137.640 ;
        RECT 24.790 135.580 24.930 137.980 ;
        RECT 30.310 136.600 30.450 137.980 ;
        RECT 31.170 137.640 31.430 137.960 ;
        RECT 30.250 136.280 30.510 136.600 ;
        RECT 26.110 135.600 26.370 135.920 ;
        RECT 24.730 135.260 24.990 135.580 ;
        RECT 26.170 133.880 26.310 135.600 ;
        RECT 26.110 133.560 26.370 133.880 ;
        RECT 30.310 132.180 30.450 136.280 ;
        RECT 31.230 133.540 31.370 137.640 ;
        RECT 32.150 135.920 32.290 138.580 ;
        RECT 32.610 136.600 32.750 138.660 ;
        RECT 66.650 137.960 66.790 141.040 ;
        RECT 66.590 137.640 66.850 137.960 ;
        RECT 36.120 136.765 37.660 137.135 ;
        RECT 32.550 136.280 32.810 136.600 ;
        RECT 32.090 135.600 32.350 135.920 ;
        RECT 65.210 135.600 65.470 135.920 ;
        RECT 31.630 134.580 31.890 134.900 ;
        RECT 31.170 133.220 31.430 133.540 ;
        RECT 26.110 131.860 26.370 132.180 ;
        RECT 30.250 131.860 30.510 132.180 ;
        RECT 26.170 130.820 26.310 131.860 ;
        RECT 26.110 130.500 26.370 130.820 ;
        RECT 24.270 130.160 24.530 130.480 ;
        RECT 21.970 127.100 22.230 127.420 ;
        RECT 21.050 126.420 21.310 126.740 ;
        RECT 20.130 124.720 20.390 125.040 ;
        RECT 19.210 123.700 19.470 124.020 ;
        RECT 19.270 122.320 19.410 123.700 ;
        RECT 19.210 122.000 19.470 122.320 ;
        RECT 20.190 120.280 20.330 124.720 ;
        RECT 21.110 123.875 21.250 126.420 ;
        RECT 21.040 123.505 21.320 123.875 ;
        RECT 21.510 121.320 21.770 121.640 ;
        RECT 21.570 120.280 21.710 121.320 ;
        RECT 22.030 121.300 22.170 127.100 ;
        RECT 21.970 120.980 22.230 121.300 ;
        RECT 22.030 120.280 22.170 120.980 ;
        RECT 24.330 120.280 24.470 130.160 ;
        RECT 25.650 127.100 25.910 127.420 ;
        RECT 25.710 125.720 25.850 127.100 ;
        RECT 26.570 126.760 26.830 127.080 ;
        RECT 25.650 125.400 25.910 125.720 ;
        RECT 26.110 124.720 26.370 125.040 ;
        RECT 26.170 124.020 26.310 124.720 ;
        RECT 26.110 123.700 26.370 124.020 ;
        RECT 26.170 121.980 26.310 123.700 ;
        RECT 26.110 121.660 26.370 121.980 ;
        RECT 20.130 119.960 20.390 120.280 ;
        RECT 21.510 119.960 21.770 120.280 ;
        RECT 21.970 119.960 22.230 120.280 ;
        RECT 24.270 119.960 24.530 120.280 ;
        RECT 20.130 119.280 20.390 119.600 ;
        RECT 20.190 117.075 20.330 119.280 ;
        RECT 24.330 117.120 24.470 119.960 ;
        RECT 26.170 119.260 26.310 121.660 ;
        RECT 26.630 119.600 26.770 126.760 ;
        RECT 31.230 124.700 31.370 133.220 ;
        RECT 31.690 132.860 31.830 134.580 ;
        RECT 31.630 132.540 31.890 132.860 ;
        RECT 31.630 126.420 31.890 126.740 ;
        RECT 31.690 125.040 31.830 126.420 ;
        RECT 31.630 124.720 31.890 125.040 ;
        RECT 31.170 124.380 31.430 124.700 ;
        RECT 29.790 123.700 30.050 124.020 ;
        RECT 28.870 122.680 29.130 123.000 ;
        RECT 27.490 120.980 27.750 121.300 ;
        RECT 26.570 119.280 26.830 119.600 ;
        RECT 26.110 118.940 26.370 119.260 ;
        RECT 20.120 116.705 20.400 117.075 ;
        RECT 24.330 116.980 24.930 117.120 ;
        RECT 24.270 113.840 24.530 114.160 ;
        RECT 23.810 113.500 24.070 113.820 ;
        RECT 20.130 111.800 20.390 112.120 ;
        RECT 18.280 109.905 18.560 110.275 ;
        RECT 18.350 109.400 18.490 109.905 ;
        RECT 18.290 109.080 18.550 109.400 ;
        RECT 20.190 108.720 20.330 111.800 ;
        RECT 20.130 108.400 20.390 108.720 ;
        RECT 21.970 108.400 22.230 108.720 ;
        RECT 18.280 106.505 18.560 106.875 ;
        RECT 16.610 103.475 17.120 103.690 ;
        RECT 16.610 103.105 17.180 103.475 ;
        RECT 16.610 102.600 17.120 103.105 ;
        RECT 16.610 102.340 17.170 102.600 ;
        RECT 16.620 102.310 17.170 102.340 ;
        RECT 16.910 102.280 17.170 102.310 ;
        RECT 18.350 102.260 18.490 106.505 ;
        RECT 19.210 104.660 19.470 104.980 ;
        RECT 19.270 103.280 19.410 104.660 ;
        RECT 22.030 103.280 22.170 108.400 ;
        RECT 23.870 103.280 24.010 113.500 ;
        RECT 24.330 112.120 24.470 113.840 ;
        RECT 24.270 111.800 24.530 112.120 ;
        RECT 24.790 106.680 24.930 116.980 ;
        RECT 26.170 113.730 26.310 118.940 ;
        RECT 27.550 114.500 27.690 120.980 ;
        RECT 27.950 118.260 28.210 118.580 ;
        RECT 27.490 114.180 27.750 114.500 ;
        RECT 27.030 113.730 27.290 113.820 ;
        RECT 26.170 113.590 27.290 113.730 ;
        RECT 27.030 113.500 27.290 113.590 ;
        RECT 25.650 112.820 25.910 113.140 ;
        RECT 25.710 111.100 25.850 112.820 ;
        RECT 27.090 111.100 27.230 113.500 ;
        RECT 27.550 111.440 27.690 114.180 ;
        RECT 27.490 111.120 27.750 111.440 ;
        RECT 25.650 110.780 25.910 111.100 ;
        RECT 27.030 110.780 27.290 111.100 ;
        RECT 27.090 107.700 27.230 110.780 ;
        RECT 27.030 107.380 27.290 107.700 ;
        RECT 24.730 106.360 24.990 106.680 ;
        RECT 27.090 105.660 27.230 107.380 ;
        RECT 28.010 105.660 28.150 118.260 ;
        RECT 28.930 116.540 29.070 122.680 ;
        RECT 29.850 121.640 29.990 123.700 ;
        RECT 29.790 121.320 30.050 121.640 ;
        RECT 29.330 119.280 29.590 119.600 ;
        RECT 28.870 116.220 29.130 116.540 ;
        RECT 28.870 115.770 29.130 115.860 ;
        RECT 29.390 115.770 29.530 119.280 ;
        RECT 29.850 118.580 29.990 121.320 ;
        RECT 30.250 119.280 30.510 119.600 ;
        RECT 29.790 118.260 30.050 118.580 ;
        RECT 29.850 116.540 29.990 118.260 ;
        RECT 29.790 116.220 30.050 116.540 ;
        RECT 28.870 115.630 29.530 115.770 ;
        RECT 28.870 115.540 29.130 115.630 ;
        RECT 28.930 108.380 29.070 115.540 ;
        RECT 30.310 114.920 30.450 119.280 ;
        RECT 29.390 114.780 30.450 114.920 ;
        RECT 28.870 108.120 29.130 108.380 ;
        RECT 28.470 108.060 29.130 108.120 ;
        RECT 28.470 107.980 29.070 108.060 ;
        RECT 27.030 105.340 27.290 105.660 ;
        RECT 27.950 105.340 28.210 105.660 ;
        RECT 25.650 105.000 25.910 105.320 ;
        RECT 25.710 103.960 25.850 105.000 ;
        RECT 25.650 103.640 25.910 103.960 ;
        RECT 19.210 102.960 19.470 103.280 ;
        RECT 21.970 102.960 22.230 103.280 ;
        RECT 23.810 102.960 24.070 103.280 ;
        RECT 25.650 102.960 25.910 103.280 ;
        RECT 18.290 101.940 18.550 102.260 ;
        RECT 25.710 98.520 25.850 102.960 ;
        RECT 26.110 101.940 26.370 102.260 ;
        RECT 25.650 98.200 25.910 98.520 ;
        RECT 15.070 94.800 15.330 95.120 ;
        RECT 13.690 92.660 13.950 92.980 ;
        RECT 12.910 91.970 13.330 92.390 ;
        RECT 15.130 87.220 15.270 94.800 ;
        RECT 18.290 94.460 18.550 94.780 ;
        RECT 24.730 94.460 24.990 94.780 ;
        RECT 15.005 86.920 15.395 87.220 ;
        RECT 15.130 86.550 15.270 86.920 ;
        RECT 18.350 86.550 18.490 94.460 ;
        RECT 21.510 93.780 21.770 94.100 ;
        RECT 21.570 92.350 21.710 93.780 ;
        RECT 21.470 92.020 21.810 92.350 ;
        RECT 21.570 86.550 21.710 92.020 ;
        RECT 24.790 88.985 24.930 94.460 ;
        RECT 25.710 94.440 25.850 98.200 ;
        RECT 26.170 98.180 26.310 101.940 ;
        RECT 27.090 100.220 27.230 105.340 ;
        RECT 28.470 102.600 28.610 107.980 ;
        RECT 28.870 103.300 29.130 103.620 ;
        RECT 28.410 102.280 28.670 102.600 ;
        RECT 27.490 101.940 27.750 102.260 ;
        RECT 27.550 100.220 27.690 101.940 ;
        RECT 27.030 99.900 27.290 100.220 ;
        RECT 27.490 99.900 27.750 100.220 ;
        RECT 26.570 99.560 26.830 99.880 ;
        RECT 26.630 98.520 26.770 99.560 ;
        RECT 26.570 98.200 26.830 98.520 ;
        RECT 26.110 97.860 26.370 98.180 ;
        RECT 27.090 97.500 27.230 99.900 ;
        RECT 27.550 98.180 27.690 99.900 ;
        RECT 28.410 99.220 28.670 99.540 ;
        RECT 28.470 98.520 28.610 99.220 ;
        RECT 28.410 98.200 28.670 98.520 ;
        RECT 27.490 97.860 27.750 98.180 ;
        RECT 27.030 97.180 27.290 97.500 ;
        RECT 27.550 94.440 27.690 97.860 ;
        RECT 28.470 94.780 28.610 98.200 ;
        RECT 28.930 95.800 29.070 103.300 ;
        RECT 29.390 102.940 29.530 114.780 ;
        RECT 30.710 113.840 30.970 114.160 ;
        RECT 30.770 112.120 30.910 113.840 ;
        RECT 30.710 111.800 30.970 112.120 ;
        RECT 30.710 110.100 30.970 110.420 ;
        RECT 30.770 109.400 30.910 110.100 ;
        RECT 30.710 109.080 30.970 109.400 ;
        RECT 29.790 105.340 30.050 105.660 ;
        RECT 29.330 102.620 29.590 102.940 ;
        RECT 29.390 97.500 29.530 102.620 ;
        RECT 29.330 97.180 29.590 97.500 ;
        RECT 29.850 95.800 29.990 105.340 ;
        RECT 30.770 98.520 30.910 109.080 ;
        RECT 31.230 106.680 31.370 124.380 ;
        RECT 32.150 121.640 32.290 135.600 ;
        RECT 32.820 134.045 34.360 134.415 ;
        RECT 65.270 133.880 65.410 135.600 ;
        RECT 66.130 134.580 66.390 134.900 ;
        RECT 65.210 133.560 65.470 133.880 ;
        RECT 61.990 132.540 62.250 132.860 ;
        RECT 32.550 132.200 32.810 132.520 ;
        RECT 35.770 132.200 36.030 132.520 ;
        RECT 32.610 130.140 32.750 132.200 ;
        RECT 34.850 131.860 35.110 132.180 ;
        RECT 32.550 129.820 32.810 130.140 ;
        RECT 32.820 128.605 34.360 128.975 ;
        RECT 34.910 124.700 35.050 131.860 ;
        RECT 35.310 124.720 35.570 125.040 ;
        RECT 34.850 124.380 35.110 124.700 ;
        RECT 32.820 123.165 34.360 123.535 ;
        RECT 34.910 121.720 35.050 124.380 ;
        RECT 35.370 123.000 35.510 124.720 ;
        RECT 35.310 122.680 35.570 123.000 ;
        RECT 32.090 121.320 32.350 121.640 ;
        RECT 34.450 121.580 35.050 121.720 ;
        RECT 34.450 119.260 34.590 121.580 ;
        RECT 34.850 120.980 35.110 121.300 ;
        RECT 34.390 118.940 34.650 119.260 ;
        RECT 34.910 118.920 35.050 120.980 ;
        RECT 35.370 119.940 35.510 122.680 ;
        RECT 35.830 120.280 35.970 132.200 ;
        RECT 36.120 131.325 37.660 131.695 ;
        RECT 62.050 130.480 62.190 132.540 ;
        RECT 64.750 132.200 65.010 132.520 ;
        RECT 61.990 130.160 62.250 130.480 ;
        RECT 64.810 128.440 64.950 132.200 ;
        RECT 64.750 128.120 65.010 128.440 ;
        RECT 66.190 127.760 66.330 134.580 ;
        RECT 66.650 130.820 66.790 137.640 ;
        RECT 67.050 135.600 67.310 135.920 ;
        RECT 68.430 135.600 68.690 135.920 ;
        RECT 67.110 134.900 67.250 135.600 ;
        RECT 67.050 134.580 67.310 134.900 ;
        RECT 67.110 132.860 67.250 134.580 ;
        RECT 68.490 133.880 68.630 135.600 ;
        RECT 68.430 133.560 68.690 133.880 ;
        RECT 67.050 132.540 67.310 132.860 ;
        RECT 68.430 131.860 68.690 132.180 ;
        RECT 66.590 130.500 66.850 130.820 ;
        RECT 66.590 129.820 66.850 130.140 ;
        RECT 66.130 127.440 66.390 127.760 ;
        RECT 36.120 125.885 37.660 126.255 ;
        RECT 36.120 120.445 37.660 120.815 ;
        RECT 35.770 119.960 36.030 120.280 ;
        RECT 35.310 119.620 35.570 119.940 ;
        RECT 35.310 118.940 35.570 119.260 ;
        RECT 34.850 118.600 35.110 118.920 ;
        RECT 32.820 117.725 34.360 118.095 ;
        RECT 32.090 114.520 32.350 114.840 ;
        RECT 32.150 111.100 32.290 114.520 ;
        RECT 32.820 112.285 34.360 112.655 ;
        RECT 32.090 110.780 32.350 111.100 ;
        RECT 32.820 106.845 34.360 107.215 ;
        RECT 31.170 106.360 31.430 106.680 ;
        RECT 35.370 106.340 35.510 118.940 ;
        RECT 36.120 115.005 37.660 115.375 ;
        RECT 66.650 114.160 66.790 129.820 ;
        RECT 68.490 126.740 68.630 131.860 ;
        RECT 68.950 127.420 69.090 146.480 ;
        RECT 70.330 146.460 70.470 148.860 ;
        RECT 73.550 147.140 73.690 150.900 ;
        RECT 73.490 146.820 73.750 147.140 ;
        RECT 70.270 146.140 70.530 146.460 ;
        RECT 70.330 144.720 70.470 146.140 ;
        RECT 75.390 144.760 75.530 151.580 ;
        RECT 76.310 148.500 76.450 153.620 ;
        RECT 78.610 152.920 78.750 159.060 ;
        RECT 86.890 156.660 87.030 170.280 ;
        RECT 87.810 170.260 87.950 170.710 ;
        RECT 88.210 170.620 88.470 170.710 ;
        RECT 89.590 170.620 89.850 170.940 ;
        RECT 87.750 169.940 88.010 170.260 ;
        RECT 88.210 169.940 88.470 170.260 ;
        RECT 87.810 167.540 87.950 169.940 ;
        RECT 88.270 168.755 88.410 169.940 ;
        RECT 88.670 168.920 88.930 169.240 ;
        RECT 88.200 168.385 88.480 168.755 ;
        RECT 88.210 167.900 88.470 168.220 ;
        RECT 87.750 167.220 88.010 167.540 ;
        RECT 88.270 162.100 88.410 167.900 ;
        RECT 88.730 163.120 88.870 168.920 ;
        RECT 89.130 168.580 89.390 168.900 ;
        RECT 88.670 162.800 88.930 163.120 ;
        RECT 88.210 161.780 88.470 162.100 ;
        RECT 88.270 161.080 88.410 161.780 ;
        RECT 88.210 160.760 88.470 161.080 ;
        RECT 89.190 160.060 89.330 168.580 ;
        RECT 89.650 168.560 89.790 170.620 ;
        RECT 89.590 168.240 89.850 168.560 ;
        RECT 91.030 160.060 91.170 174.020 ;
        RECT 92.350 171.640 92.610 171.960 ;
        RECT 92.410 168.560 92.550 171.640 ;
        RECT 92.350 168.240 92.610 168.560 ;
        RECT 93.270 162.460 93.530 162.780 ;
        RECT 89.130 159.740 89.390 160.060 ;
        RECT 90.970 159.740 91.230 160.060 ;
        RECT 92.810 159.400 93.070 159.720 ;
        RECT 88.210 159.060 88.470 159.380 ;
        RECT 87.290 157.020 87.550 157.340 ;
        RECT 86.830 156.340 87.090 156.660 ;
        RECT 79.010 154.300 79.270 154.620 ;
        RECT 79.930 154.300 80.190 154.620 ;
        RECT 78.550 152.600 78.810 152.920 ;
        RECT 78.090 151.580 78.350 151.900 ;
        RECT 76.710 150.900 76.970 151.220 ;
        RECT 76.770 150.200 76.910 150.900 ;
        RECT 76.710 149.880 76.970 150.200 ;
        RECT 78.150 149.860 78.290 151.580 ;
        RECT 78.090 149.540 78.350 149.860 ;
        RECT 77.170 149.200 77.430 149.520 ;
        RECT 76.250 148.180 76.510 148.500 ;
        RECT 69.870 144.580 70.470 144.720 ;
        RECT 69.870 141.020 70.010 144.580 ;
        RECT 75.330 144.440 75.590 144.760 ;
        RECT 72.110 143.420 72.370 143.740 ;
        RECT 69.810 140.700 70.070 141.020 ;
        RECT 69.870 135.920 70.010 140.700 ;
        RECT 70.270 138.320 70.530 138.640 ;
        RECT 70.330 137.620 70.470 138.320 ;
        RECT 70.270 137.300 70.530 137.620 ;
        RECT 69.810 135.600 70.070 135.920 ;
        RECT 72.170 133.200 72.310 143.420 ;
        RECT 77.230 141.700 77.370 149.200 ;
        RECT 78.150 142.040 78.290 149.540 ;
        RECT 79.070 148.840 79.210 154.300 ;
        RECT 79.470 153.620 79.730 153.940 ;
        RECT 79.530 151.900 79.670 153.620 ;
        RECT 79.470 151.580 79.730 151.900 ;
        RECT 79.530 149.180 79.670 151.580 ;
        RECT 79.470 148.860 79.730 149.180 ;
        RECT 78.550 148.520 78.810 148.840 ;
        RECT 79.010 148.520 79.270 148.840 ;
        RECT 78.610 147.140 78.750 148.520 ;
        RECT 79.070 147.480 79.210 148.520 ;
        RECT 79.470 148.240 79.730 148.500 ;
        RECT 79.990 148.240 80.130 154.300 ;
        RECT 83.610 153.620 83.870 153.940 ;
        RECT 80.390 152.600 80.650 152.920 ;
        RECT 80.450 149.180 80.590 152.600 ;
        RECT 83.670 151.220 83.810 153.620 ;
        RECT 86.370 152.260 86.630 152.580 ;
        RECT 85.910 151.920 86.170 152.240 ;
        RECT 83.610 150.900 83.870 151.220 ;
        RECT 83.670 149.520 83.810 150.900 ;
        RECT 85.970 150.200 86.110 151.920 ;
        RECT 86.430 150.200 86.570 152.260 ;
        RECT 85.910 149.880 86.170 150.200 ;
        RECT 86.370 149.880 86.630 150.200 ;
        RECT 83.610 149.200 83.870 149.520 ;
        RECT 80.390 148.860 80.650 149.180 ;
        RECT 81.770 148.520 82.030 148.840 ;
        RECT 79.470 148.180 80.130 148.240 ;
        RECT 79.530 148.100 80.130 148.180 ;
        RECT 79.010 147.160 79.270 147.480 ;
        RECT 78.550 146.820 78.810 147.140 ;
        RECT 78.610 144.420 78.750 146.820 ;
        RECT 79.070 146.460 79.210 147.160 ;
        RECT 79.010 146.140 79.270 146.460 ;
        RECT 79.530 146.120 79.670 148.100 ;
        RECT 79.930 146.480 80.190 146.800 ;
        RECT 79.470 145.800 79.730 146.120 ;
        RECT 78.550 144.100 78.810 144.420 ;
        RECT 79.530 143.740 79.670 145.800 ;
        RECT 79.990 144.760 80.130 146.480 ;
        RECT 81.830 146.460 81.970 148.520 ;
        RECT 81.770 146.140 82.030 146.460 ;
        RECT 82.230 146.140 82.490 146.460 ;
        RECT 79.930 144.440 80.190 144.760 ;
        RECT 79.470 143.420 79.730 143.740 ;
        RECT 78.090 141.720 78.350 142.040 ;
        RECT 77.170 141.610 77.430 141.700 ;
        RECT 77.170 141.470 77.830 141.610 ;
        RECT 77.170 141.380 77.430 141.470 ;
        RECT 76.250 140.700 76.510 141.020 ;
        RECT 76.310 139.320 76.450 140.700 ;
        RECT 72.570 139.000 72.830 139.320 ;
        RECT 76.250 139.000 76.510 139.320 ;
        RECT 72.110 132.880 72.370 133.200 ;
        RECT 72.170 131.160 72.310 132.880 ;
        RECT 72.110 130.840 72.370 131.160 ;
        RECT 70.730 130.160 70.990 130.480 ;
        RECT 70.790 128.440 70.930 130.160 ;
        RECT 70.730 128.120 70.990 128.440 ;
        RECT 72.630 127.760 72.770 139.000 ;
        RECT 73.490 138.660 73.750 138.980 ;
        RECT 73.550 136.600 73.690 138.660 ;
        RECT 73.950 138.320 74.210 138.640 ;
        RECT 73.490 136.280 73.750 136.600 ;
        RECT 74.010 132.860 74.150 138.320 ;
        RECT 76.310 134.900 76.450 139.000 ;
        RECT 77.170 137.980 77.430 138.300 ;
        RECT 77.230 135.920 77.370 137.980 ;
        RECT 77.690 137.620 77.830 141.470 ;
        RECT 81.830 141.020 81.970 146.140 ;
        RECT 82.290 144.760 82.430 146.140 ;
        RECT 82.230 144.440 82.490 144.760 ;
        RECT 83.670 144.720 83.810 149.200 ;
        RECT 86.370 148.180 86.630 148.500 ;
        RECT 86.430 145.780 86.570 148.180 ;
        RECT 85.450 145.460 85.710 145.780 ;
        RECT 86.370 145.460 86.630 145.780 ;
        RECT 83.210 144.580 83.810 144.720 ;
        RECT 82.690 141.040 82.950 141.360 ;
        RECT 81.770 140.700 82.030 141.020 ;
        RECT 82.750 138.300 82.890 141.040 ;
        RECT 82.690 137.980 82.950 138.300 ;
        RECT 77.630 137.300 77.890 137.620 ;
        RECT 77.690 135.920 77.830 137.300 ;
        RECT 82.750 136.000 82.890 137.980 ;
        RECT 82.290 135.920 82.890 136.000 ;
        RECT 77.170 135.600 77.430 135.920 ;
        RECT 77.630 135.600 77.890 135.920 ;
        RECT 82.230 135.860 82.890 135.920 ;
        RECT 82.230 135.600 82.490 135.860 ;
        RECT 76.250 134.580 76.510 134.900 ;
        RECT 76.310 133.880 76.450 134.580 ;
        RECT 77.230 133.880 77.370 135.600 ;
        RECT 80.390 135.320 80.650 135.580 ;
        RECT 80.390 135.260 81.970 135.320 ;
        RECT 80.450 135.240 81.970 135.260 ;
        RECT 80.450 135.180 82.030 135.240 ;
        RECT 81.770 134.920 82.030 135.180 ;
        RECT 79.930 134.580 80.190 134.900 ;
        RECT 82.230 134.580 82.490 134.900 ;
        RECT 79.990 133.880 80.130 134.580 ;
        RECT 76.250 133.560 76.510 133.880 ;
        RECT 77.170 133.560 77.430 133.880 ;
        RECT 79.930 133.560 80.190 133.880 ;
        RECT 73.950 132.540 74.210 132.860 ;
        RECT 73.030 129.140 73.290 129.460 ;
        RECT 77.170 129.140 77.430 129.460 ;
        RECT 72.570 127.440 72.830 127.760 ;
        RECT 68.890 127.100 69.150 127.420 ;
        RECT 73.090 127.080 73.230 129.140 ;
        RECT 77.230 127.080 77.370 129.140 ;
        RECT 82.290 127.760 82.430 134.580 ;
        RECT 82.690 130.160 82.950 130.480 ;
        RECT 82.750 128.440 82.890 130.160 ;
        RECT 82.690 128.120 82.950 128.440 ;
        RECT 82.230 127.440 82.490 127.760 ;
        RECT 73.030 126.760 73.290 127.080 ;
        RECT 77.170 126.760 77.430 127.080 ;
        RECT 68.430 126.420 68.690 126.740 ;
        RECT 71.650 126.420 71.910 126.740 ;
        RECT 66.590 113.840 66.850 114.160 ;
        RECT 66.650 111.100 66.790 113.840 ;
        RECT 68.430 111.460 68.690 111.780 ;
        RECT 61.530 110.780 61.790 111.100 ;
        RECT 66.590 110.780 66.850 111.100 ;
        RECT 36.120 109.565 37.660 109.935 ;
        RECT 35.310 106.080 35.570 106.340 ;
        RECT 34.450 106.020 35.570 106.080 ;
        RECT 34.450 105.940 35.510 106.020 ;
        RECT 34.450 105.660 34.590 105.940 ;
        RECT 61.070 105.680 61.330 106.000 ;
        RECT 32.550 105.340 32.810 105.660 ;
        RECT 34.390 105.340 34.650 105.660 ;
        RECT 35.310 105.340 35.570 105.660 ;
        RECT 31.170 105.000 31.430 105.320 ;
        RECT 31.230 103.280 31.370 105.000 ;
        RECT 31.170 102.960 31.430 103.280 ;
        RECT 32.090 103.190 32.350 103.280 ;
        RECT 31.690 103.050 32.350 103.190 ;
        RECT 31.690 100.640 31.830 103.050 ;
        RECT 32.090 102.960 32.350 103.050 ;
        RECT 32.610 102.170 32.750 105.340 ;
        RECT 33.930 104.660 34.190 104.980 ;
        RECT 33.470 102.960 33.730 103.280 ;
        RECT 33.530 102.260 33.670 102.960 ;
        RECT 33.990 102.260 34.130 104.660 ;
        RECT 35.370 103.620 35.510 105.340 ;
        RECT 35.770 104.660 36.030 104.980 ;
        RECT 35.310 103.300 35.570 103.620 ;
        RECT 35.310 102.620 35.570 102.940 ;
        RECT 32.150 102.030 32.750 102.170 ;
        RECT 32.150 101.240 32.290 102.030 ;
        RECT 33.470 101.940 33.730 102.260 ;
        RECT 33.930 101.940 34.190 102.260 ;
        RECT 34.850 101.940 35.110 102.260 ;
        RECT 32.820 101.405 34.360 101.775 ;
        RECT 32.090 100.920 32.350 101.240 ;
        RECT 31.690 100.500 32.750 100.640 ;
        RECT 32.610 100.220 32.750 100.500 ;
        RECT 32.090 99.900 32.350 100.220 ;
        RECT 32.550 99.900 32.810 100.220 ;
        RECT 33.930 99.900 34.190 100.220 ;
        RECT 31.170 99.220 31.430 99.540 ;
        RECT 30.710 98.200 30.970 98.520 ;
        RECT 31.230 97.840 31.370 99.220 ;
        RECT 31.170 97.520 31.430 97.840 ;
        RECT 28.870 95.480 29.130 95.800 ;
        RECT 29.790 95.480 30.050 95.800 ;
        RECT 32.150 95.710 32.290 99.900 ;
        RECT 32.610 96.820 32.750 99.900 ;
        RECT 33.470 99.560 33.730 99.880 ;
        RECT 33.530 97.840 33.670 99.560 ;
        RECT 33.990 98.520 34.130 99.900 ;
        RECT 33.930 98.200 34.190 98.520 ;
        RECT 33.470 97.520 33.730 97.840 ;
        RECT 32.550 96.500 32.810 96.820 ;
        RECT 32.820 95.965 34.360 96.335 ;
        RECT 32.150 95.570 33.670 95.710 ;
        RECT 33.530 94.780 33.670 95.570 ;
        RECT 34.910 95.460 35.050 101.940 ;
        RECT 35.370 100.560 35.510 102.620 ;
        RECT 35.310 100.240 35.570 100.560 ;
        RECT 35.310 99.220 35.570 99.540 ;
        RECT 35.370 98.180 35.510 99.220 ;
        RECT 35.310 97.860 35.570 98.180 ;
        RECT 35.310 97.410 35.570 97.500 ;
        RECT 35.830 97.410 35.970 104.660 ;
        RECT 36.120 104.125 37.660 104.495 ;
        RECT 61.130 103.620 61.270 105.680 ;
        RECT 36.690 103.300 36.950 103.620 ;
        RECT 61.070 103.300 61.330 103.620 ;
        RECT 36.750 99.880 36.890 103.300 ;
        RECT 61.590 103.280 61.730 110.780 ;
        RECT 64.750 110.440 65.010 110.760 ;
        RECT 64.810 109.400 64.950 110.440 ;
        RECT 64.750 109.080 65.010 109.400 ;
        RECT 68.490 109.060 68.630 111.460 ;
        RECT 71.190 111.120 71.450 111.440 ;
        RECT 70.270 110.100 70.530 110.420 ;
        RECT 70.730 110.100 70.990 110.420 ;
        RECT 67.050 108.740 67.310 109.060 ;
        RECT 68.430 108.740 68.690 109.060 ;
        RECT 67.110 106.000 67.250 108.740 ;
        RECT 69.350 106.020 69.610 106.340 ;
        RECT 67.050 105.680 67.310 106.000 ;
        RECT 68.430 105.340 68.690 105.660 ;
        RECT 64.290 104.660 64.550 104.980 ;
        RECT 67.050 104.660 67.310 104.980 ;
        RECT 64.350 103.620 64.490 104.660 ;
        RECT 64.290 103.300 64.550 103.620 ;
        RECT 38.530 102.960 38.790 103.280 ;
        RECT 39.910 102.960 40.170 103.280 ;
        RECT 41.290 102.960 41.550 103.280 ;
        RECT 41.750 102.960 42.010 103.280 ;
        RECT 61.530 102.960 61.790 103.280 ;
        RECT 64.750 102.960 65.010 103.280 ;
        RECT 38.070 101.940 38.330 102.260 ;
        RECT 36.690 99.560 36.950 99.880 ;
        RECT 36.120 98.685 37.660 99.055 ;
        RECT 37.610 97.520 37.870 97.840 ;
        RECT 35.310 97.270 35.970 97.410 ;
        RECT 35.310 97.180 35.570 97.270 ;
        RECT 36.230 97.180 36.490 97.500 ;
        RECT 36.290 95.800 36.430 97.180 ;
        RECT 36.690 96.500 36.950 96.820 ;
        RECT 36.750 95.800 36.890 96.500 ;
        RECT 36.230 95.480 36.490 95.800 ;
        RECT 36.690 95.480 36.950 95.800 ;
        RECT 37.670 95.460 37.810 97.520 ;
        RECT 38.130 95.460 38.270 101.940 ;
        RECT 38.590 97.840 38.730 102.960 ;
        RECT 39.450 100.240 39.710 100.560 ;
        RECT 39.510 99.960 39.650 100.240 ;
        RECT 39.050 99.820 39.650 99.960 ;
        RECT 38.530 97.520 38.790 97.840 ;
        RECT 39.050 96.820 39.190 99.820 ;
        RECT 39.970 99.540 40.110 102.960 ;
        RECT 40.830 102.620 41.090 102.940 ;
        RECT 40.370 99.900 40.630 100.220 ;
        RECT 39.910 99.280 40.170 99.540 ;
        RECT 39.510 99.220 40.170 99.280 ;
        RECT 39.510 99.140 40.110 99.220 ;
        RECT 39.510 97.840 39.650 99.140 ;
        RECT 39.450 97.520 39.710 97.840 ;
        RECT 38.990 96.500 39.250 96.820 ;
        RECT 34.850 95.140 35.110 95.460 ;
        RECT 37.610 95.140 37.870 95.460 ;
        RECT 38.070 95.140 38.330 95.460 ;
        RECT 28.410 94.460 28.670 94.780 ;
        RECT 31.170 94.460 31.430 94.780 ;
        RECT 33.470 94.460 33.730 94.780 ;
        RECT 34.850 94.690 35.110 94.780 ;
        RECT 34.450 94.550 35.110 94.690 ;
        RECT 25.650 94.120 25.910 94.440 ;
        RECT 27.490 94.120 27.750 94.440 ;
        RECT 27.950 93.780 28.210 94.100 ;
        RECT 28.010 92.950 28.150 93.780 ;
        RECT 27.920 92.690 28.240 92.950 ;
        RECT 24.710 88.595 25.010 88.985 ;
        RECT 24.790 86.550 24.930 88.595 ;
        RECT 28.010 86.550 28.150 92.690 ;
        RECT 31.230 86.550 31.370 94.460 ;
        RECT 33.530 93.080 33.670 94.460 ;
        RECT 33.470 92.760 33.730 93.080 ;
        RECT 34.450 91.090 34.590 94.550 ;
        RECT 34.850 94.460 35.110 94.550 ;
        RECT 38.070 94.460 38.330 94.780 ;
        RECT 36.120 93.245 37.660 93.615 ;
        RECT 34.825 91.090 35.215 91.170 ;
        RECT 34.450 90.950 35.215 91.090 ;
        RECT 34.450 86.550 34.590 90.950 ;
        RECT 34.825 90.870 35.215 90.950 ;
        RECT 38.130 89.080 38.270 94.460 ;
        RECT 39.050 94.100 39.190 96.500 ;
        RECT 39.510 95.800 39.650 97.520 ;
        RECT 40.430 97.500 40.570 99.900 ;
        RECT 40.890 99.880 41.030 102.620 ;
        RECT 41.350 100.900 41.490 102.960 ;
        RECT 41.290 100.580 41.550 100.900 ;
        RECT 40.830 99.560 41.090 99.880 ;
        RECT 40.890 97.840 41.030 99.560 ;
        RECT 41.810 98.520 41.950 102.960 ;
        RECT 43.590 102.280 43.850 102.600 ;
        RECT 42.210 100.920 42.470 101.240 ;
        RECT 41.750 98.200 42.010 98.520 ;
        RECT 42.270 97.840 42.410 100.920 ;
        RECT 43.650 98.520 43.790 102.280 ;
        RECT 44.510 101.940 44.770 102.260 ;
        RECT 58.770 101.940 59.030 102.260 ;
        RECT 43.590 98.200 43.850 98.520 ;
        RECT 44.570 97.840 44.710 101.940 ;
        RECT 48.190 100.580 48.450 100.900 ;
        RECT 46.810 99.900 47.070 100.220 ;
        RECT 45.890 99.220 46.150 99.540 ;
        RECT 45.950 97.840 46.090 99.220 ;
        RECT 40.830 97.520 41.090 97.840 ;
        RECT 42.210 97.520 42.470 97.840 ;
        RECT 44.510 97.520 44.770 97.840 ;
        RECT 45.890 97.520 46.150 97.840 ;
        RECT 40.370 97.180 40.630 97.500 ;
        RECT 40.890 95.800 41.030 97.520 ;
        RECT 39.450 95.480 39.710 95.800 ;
        RECT 40.830 95.480 41.090 95.800 ;
        RECT 42.270 95.460 42.410 97.520 ;
        RECT 42.210 95.140 42.470 95.460 ;
        RECT 40.830 94.460 41.090 94.780 ;
        RECT 44.050 94.460 44.310 94.780 ;
        RECT 38.990 93.780 39.250 94.100 ;
        RECT 40.890 89.770 41.030 94.460 ;
        RECT 44.110 90.620 44.250 94.460 ;
        RECT 45.950 94.440 46.090 97.520 ;
        RECT 46.870 96.820 47.010 99.900 ;
        RECT 48.250 98.520 48.390 100.580 ;
        RECT 58.830 99.880 58.970 101.940 ;
        RECT 61.590 101.240 61.730 102.960 ;
        RECT 61.530 100.920 61.790 101.240 ;
        RECT 61.590 100.220 61.730 100.920 ;
        RECT 61.530 99.900 61.790 100.220 ;
        RECT 58.770 99.560 59.030 99.880 ;
        RECT 48.190 98.200 48.450 98.520 ;
        RECT 61.590 98.180 61.730 99.900 ;
        RECT 61.530 97.860 61.790 98.180 ;
        RECT 56.930 97.520 57.190 97.840 ;
        RECT 61.990 97.520 62.250 97.840 ;
        RECT 46.810 96.500 47.070 96.820 ;
        RECT 48.650 96.500 48.910 96.820 ;
        RECT 48.710 95.800 48.850 96.500 ;
        RECT 48.650 95.480 48.910 95.800 ;
        RECT 47.270 94.460 47.530 94.780 ;
        RECT 50.490 94.460 50.750 94.780 ;
        RECT 53.710 94.460 53.970 94.780 ;
        RECT 45.890 94.120 46.150 94.440 ;
        RECT 47.330 92.175 47.470 94.460 ;
        RECT 47.730 93.780 47.990 94.100 ;
        RECT 47.790 93.080 47.930 93.780 ;
        RECT 47.730 92.760 47.990 93.080 ;
        RECT 47.250 91.785 47.550 92.175 ;
        RECT 43.920 89.980 45.010 90.620 ;
        RECT 40.730 89.320 41.420 89.770 ;
        RECT 37.670 88.940 38.270 89.080 ;
        RECT 37.670 86.550 37.810 88.940 ;
        RECT 40.890 86.550 41.030 89.320 ;
        RECT 44.110 86.550 44.250 89.980 ;
        RECT 11.840 81.280 12.120 86.550 ;
        RECT 15.060 82.550 15.340 86.550 ;
        RECT 18.280 85.910 18.560 86.550 ;
        RECT 18.180 85.490 18.640 85.910 ;
        RECT 18.280 82.550 18.560 85.490 ;
        RECT 21.500 82.550 21.780 86.550 ;
        RECT 24.720 82.550 25.000 86.550 ;
        RECT 27.940 82.550 28.220 86.550 ;
        RECT 31.160 81.990 31.440 86.550 ;
        RECT 34.380 82.550 34.660 86.550 ;
        RECT 37.600 82.550 37.880 86.550 ;
        RECT 40.820 82.550 41.100 86.550 ;
        RECT 44.040 82.550 44.320 86.550 ;
        RECT 47.260 82.550 47.540 91.785 ;
        RECT 50.550 88.180 50.690 94.460 ;
        RECT 50.360 87.680 51.620 88.180 ;
        RECT 50.550 86.550 50.690 87.680 ;
        RECT 53.770 86.550 53.910 94.460 ;
        RECT 56.990 86.550 57.130 97.520 ;
        RECT 62.050 95.800 62.190 97.520 ;
        RECT 61.990 95.480 62.250 95.800 ;
        RECT 60.150 95.140 60.410 95.460 ;
        RECT 57.850 94.460 58.110 94.780 ;
        RECT 57.910 93.080 58.050 94.460 ;
        RECT 57.850 92.760 58.110 93.080 ;
        RECT 60.210 86.550 60.350 95.140 ;
        RECT 64.810 94.440 64.950 102.960 ;
        RECT 66.130 101.940 66.390 102.260 ;
        RECT 66.190 94.440 66.330 101.940 ;
        RECT 67.110 95.460 67.250 104.660 ;
        RECT 68.490 101.240 68.630 105.340 ;
        RECT 68.890 104.660 69.150 104.980 ;
        RECT 68.430 100.920 68.690 101.240 ;
        RECT 68.430 99.900 68.690 100.220 ;
        RECT 67.970 99.560 68.230 99.880 ;
        RECT 67.510 98.200 67.770 98.520 ;
        RECT 67.050 95.140 67.310 95.460 ;
        RECT 67.570 94.780 67.710 98.200 ;
        RECT 68.030 95.800 68.170 99.560 ;
        RECT 68.490 96.420 68.630 99.900 ;
        RECT 68.950 98.520 69.090 104.660 ;
        RECT 69.410 103.960 69.550 106.020 ;
        RECT 69.350 103.640 69.610 103.960 ;
        RECT 70.330 100.220 70.470 110.100 ;
        RECT 70.790 108.040 70.930 110.100 ;
        RECT 70.730 107.720 70.990 108.040 ;
        RECT 71.250 106.000 71.390 111.120 ;
        RECT 71.710 108.380 71.850 126.420 ;
        RECT 73.090 117.640 73.230 126.760 ;
        RECT 80.390 119.960 80.650 120.280 ;
        RECT 79.010 119.280 79.270 119.600 ;
        RECT 73.950 118.940 74.210 119.260 ;
        RECT 72.630 117.500 73.230 117.640 ;
        RECT 72.630 111.100 72.770 117.500 ;
        RECT 73.030 116.560 73.290 116.880 ;
        RECT 73.090 114.840 73.230 116.560 ;
        RECT 74.010 115.860 74.150 118.940 ;
        RECT 76.250 118.260 76.510 118.580 ;
        RECT 76.310 116.200 76.450 118.260 ;
        RECT 76.250 115.880 76.510 116.200 ;
        RECT 73.490 115.540 73.750 115.860 ;
        RECT 73.950 115.540 74.210 115.860 ;
        RECT 73.030 114.520 73.290 114.840 ;
        RECT 73.550 114.500 73.690 115.540 ;
        RECT 73.490 114.180 73.750 114.500 ;
        RECT 74.010 111.780 74.150 115.540 ;
        RECT 79.070 113.140 79.210 119.280 ;
        RECT 79.930 118.600 80.190 118.920 ;
        RECT 79.990 115.860 80.130 118.600 ;
        RECT 79.930 115.540 80.190 115.860 ;
        RECT 79.990 114.840 80.130 115.540 ;
        RECT 79.930 114.520 80.190 114.840 ;
        RECT 77.630 112.820 77.890 113.140 ;
        RECT 79.010 112.820 79.270 113.140 ;
        RECT 73.950 111.460 74.210 111.780 ;
        RECT 72.570 110.780 72.830 111.100 ;
        RECT 74.010 110.840 74.150 111.460 ;
        RECT 73.550 110.700 74.150 110.840 ;
        RECT 71.650 108.060 71.910 108.380 ;
        RECT 71.190 105.680 71.450 106.000 ;
        RECT 70.730 103.640 70.990 103.960 ;
        RECT 70.790 103.475 70.930 103.640 ;
        RECT 70.720 103.105 71.000 103.475 ;
        RECT 71.250 102.680 71.390 105.680 ;
        RECT 71.710 103.475 71.850 108.060 ;
        RECT 72.110 105.000 72.370 105.320 ;
        RECT 73.030 105.000 73.290 105.320 ;
        RECT 72.170 103.620 72.310 105.000 ;
        RECT 73.090 103.960 73.230 105.000 ;
        RECT 73.030 103.640 73.290 103.960 ;
        RECT 71.640 103.105 71.920 103.475 ;
        RECT 72.110 103.300 72.370 103.620 ;
        RECT 71.650 102.680 71.910 102.940 ;
        RECT 71.250 102.620 71.910 102.680 ;
        RECT 71.250 102.540 71.850 102.620 ;
        RECT 71.190 100.920 71.450 101.240 ;
        RECT 70.270 99.900 70.530 100.220 ;
        RECT 69.810 99.560 70.070 99.880 ;
        RECT 68.890 98.200 69.150 98.520 ;
        RECT 68.950 97.160 69.090 98.200 ;
        RECT 68.890 96.840 69.150 97.160 ;
        RECT 69.350 96.500 69.610 96.820 ;
        RECT 68.490 96.280 69.090 96.420 ;
        RECT 67.970 95.480 68.230 95.800 ;
        RECT 67.510 94.460 67.770 94.780 ;
        RECT 63.370 94.120 63.630 94.440 ;
        RECT 64.750 94.120 65.010 94.440 ;
        RECT 66.130 94.120 66.390 94.440 ;
        RECT 63.430 86.550 63.570 94.120 ;
        RECT 66.590 93.780 66.850 94.100 ;
        RECT 66.650 86.550 66.790 93.780 ;
        RECT 68.950 93.080 69.090 96.280 ;
        RECT 69.410 95.460 69.550 96.500 ;
        RECT 69.350 95.140 69.610 95.460 ;
        RECT 68.890 92.760 69.150 93.080 ;
        RECT 69.870 86.550 70.010 99.560 ;
        RECT 71.250 96.420 71.390 100.920 ;
        RECT 72.170 99.960 72.310 103.300 ;
        RECT 73.090 100.220 73.230 103.640 ;
        RECT 73.550 103.280 73.690 110.700 ;
        RECT 74.410 105.680 74.670 106.000 ;
        RECT 73.950 103.640 74.210 103.960 ;
        RECT 73.490 102.960 73.750 103.280 ;
        RECT 71.710 99.820 72.310 99.960 ;
        RECT 73.030 99.900 73.290 100.220 ;
        RECT 71.710 97.840 71.850 99.820 ;
        RECT 72.110 99.220 72.370 99.540 ;
        RECT 72.170 98.520 72.310 99.220 ;
        RECT 72.110 98.200 72.370 98.520 ;
        RECT 71.650 97.520 71.910 97.840 ;
        RECT 73.490 97.520 73.750 97.840 ;
        RECT 72.570 97.180 72.830 97.500 ;
        RECT 71.250 96.280 71.850 96.420 ;
        RECT 71.180 94.945 71.460 95.315 ;
        RECT 71.710 95.120 71.850 96.280 ;
        RECT 72.630 95.120 72.770 97.180 ;
        RECT 71.250 94.780 71.390 94.945 ;
        RECT 71.650 94.800 71.910 95.120 ;
        RECT 72.570 94.800 72.830 95.120 ;
        RECT 73.550 94.780 73.690 97.520 ;
        RECT 74.010 97.500 74.150 103.640 ;
        RECT 74.470 98.180 74.610 105.680 ;
        RECT 75.330 105.000 75.590 105.320 ;
        RECT 74.410 97.860 74.670 98.180 ;
        RECT 75.390 97.840 75.530 105.000 ;
        RECT 75.790 101.940 76.050 102.260 ;
        RECT 75.850 99.880 75.990 101.940 ;
        RECT 75.790 99.560 76.050 99.880 ;
        RECT 75.330 97.520 75.590 97.840 ;
        RECT 73.950 97.180 74.210 97.500 ;
        RECT 77.690 94.780 77.830 112.820 ;
        RECT 79.070 111.440 79.210 112.820 ;
        RECT 79.010 111.120 79.270 111.440 ;
        RECT 78.090 110.780 78.350 111.100 ;
        RECT 78.150 108.040 78.290 110.780 ;
        RECT 78.090 107.720 78.350 108.040 ;
        RECT 78.150 103.280 78.290 107.720 ;
        RECT 79.470 107.380 79.730 107.700 ;
        RECT 79.530 103.620 79.670 107.380 ;
        RECT 79.470 103.300 79.730 103.620 ;
        RECT 78.090 102.960 78.350 103.280 ;
        RECT 78.090 102.280 78.350 102.600 ;
        RECT 78.150 99.540 78.290 102.280 ;
        RECT 78.090 99.220 78.350 99.540 ;
        RECT 78.150 94.780 78.290 99.220 ;
        RECT 79.990 94.780 80.130 114.520 ;
        RECT 80.450 114.500 80.590 119.960 ;
        RECT 80.850 116.220 81.110 116.540 ;
        RECT 80.390 114.180 80.650 114.500 ;
        RECT 80.910 103.280 81.050 116.220 ;
        RECT 83.210 107.700 83.350 144.580 ;
        RECT 85.510 143.740 85.650 145.460 ;
        RECT 85.450 143.420 85.710 143.740 ;
        RECT 85.910 141.380 86.170 141.700 ;
        RECT 85.450 141.040 85.710 141.360 ;
        RECT 85.510 139.320 85.650 141.040 ;
        RECT 85.450 139.000 85.710 139.320 ;
        RECT 85.970 138.300 86.110 141.380 ;
        RECT 86.370 140.700 86.630 141.020 ;
        RECT 85.910 137.980 86.170 138.300 ;
        RECT 85.970 135.920 86.110 137.980 ;
        RECT 85.910 135.600 86.170 135.920 ;
        RECT 84.530 134.580 84.790 134.900 ;
        RECT 84.590 133.200 84.730 134.580 ;
        RECT 84.530 132.880 84.790 133.200 ;
        RECT 86.430 132.860 86.570 140.700 ;
        RECT 86.890 137.960 87.030 156.340 ;
        RECT 87.350 155.640 87.490 157.020 ;
        RECT 87.290 155.320 87.550 155.640 ;
        RECT 87.750 148.860 88.010 149.180 ;
        RECT 87.810 147.480 87.950 148.860 ;
        RECT 88.270 148.840 88.410 159.060 ;
        RECT 92.870 158.360 93.010 159.400 ;
        RECT 92.810 158.040 93.070 158.360 ;
        RECT 90.510 152.260 90.770 152.580 ;
        RECT 90.570 149.520 90.710 152.260 ;
        RECT 90.510 149.200 90.770 149.520 ;
        RECT 88.210 148.520 88.470 148.840 ;
        RECT 87.750 147.160 88.010 147.480 ;
        RECT 87.750 146.140 88.010 146.460 ;
        RECT 87.290 145.460 87.550 145.780 ;
        RECT 87.350 143.740 87.490 145.460 ;
        RECT 87.810 144.080 87.950 146.140 ;
        RECT 87.750 143.760 88.010 144.080 ;
        RECT 87.290 143.420 87.550 143.740 ;
        RECT 87.350 141.360 87.490 143.420 ;
        RECT 87.290 141.040 87.550 141.360 ;
        RECT 87.290 140.020 87.550 140.340 ;
        RECT 87.350 138.640 87.490 140.020 ;
        RECT 87.290 138.320 87.550 138.640 ;
        RECT 86.830 137.640 87.090 137.960 ;
        RECT 87.810 136.000 87.950 143.760 ;
        RECT 89.590 143.080 89.850 143.400 ;
        RECT 89.650 142.040 89.790 143.080 ;
        RECT 89.590 141.720 89.850 142.040 ;
        RECT 90.050 140.700 90.310 141.020 ;
        RECT 90.110 138.300 90.250 140.700 ;
        RECT 93.330 138.300 93.470 162.460 ;
        RECT 94.190 160.760 94.450 161.080 ;
        RECT 94.250 154.960 94.390 160.760 ;
        RECT 95.630 158.360 95.770 180.820 ;
        RECT 96.090 176.380 96.230 180.820 ;
        RECT 96.030 176.060 96.290 176.380 ;
        RECT 96.030 159.060 96.290 159.380 ;
        RECT 95.570 158.040 95.830 158.360 ;
        RECT 94.190 154.640 94.450 154.960 ;
        RECT 93.730 153.960 93.990 154.280 ;
        RECT 93.790 152.920 93.930 153.960 ;
        RECT 93.730 152.600 93.990 152.920 ;
        RECT 93.790 151.900 93.930 152.600 ;
        RECT 94.250 152.580 94.390 154.640 ;
        RECT 94.650 153.960 94.910 154.280 ;
        RECT 94.190 152.260 94.450 152.580 ;
        RECT 93.730 151.580 93.990 151.900 ;
        RECT 94.710 151.560 94.850 153.960 ;
        RECT 94.650 151.240 94.910 151.560 ;
        RECT 94.190 150.900 94.450 151.220 ;
        RECT 94.250 149.180 94.390 150.900 ;
        RECT 94.190 148.860 94.450 149.180 ;
        RECT 95.110 142.740 95.370 143.060 ;
        RECT 95.170 142.040 95.310 142.740 ;
        RECT 95.110 141.720 95.370 142.040 ;
        RECT 90.050 137.980 90.310 138.300 ;
        RECT 93.270 137.980 93.530 138.300 ;
        RECT 89.590 137.640 89.850 137.960 ;
        RECT 88.210 137.300 88.470 137.620 ;
        RECT 88.270 136.260 88.410 137.300 ;
        RECT 87.350 135.920 87.950 136.000 ;
        RECT 88.210 135.940 88.470 136.260 ;
        RECT 87.290 135.860 87.950 135.920 ;
        RECT 87.290 135.600 87.550 135.860 ;
        RECT 87.810 133.200 87.950 135.860 ;
        RECT 87.750 132.880 88.010 133.200 ;
        RECT 86.370 132.540 86.630 132.860 ;
        RECT 86.430 127.420 86.570 132.540 ;
        RECT 86.830 131.860 87.090 132.180 ;
        RECT 86.890 130.480 87.030 131.860 ;
        RECT 87.810 130.820 87.950 132.880 ;
        RECT 87.750 130.500 88.010 130.820 ;
        RECT 86.830 130.160 87.090 130.480 ;
        RECT 86.370 127.100 86.630 127.420 ;
        RECT 86.370 126.420 86.630 126.740 ;
        RECT 85.910 121.320 86.170 121.640 ;
        RECT 83.610 119.620 83.870 119.940 ;
        RECT 83.670 114.500 83.810 119.620 ;
        RECT 85.450 118.940 85.710 119.260 ;
        RECT 84.070 118.260 84.330 118.580 ;
        RECT 83.610 114.180 83.870 114.500 ;
        RECT 83.150 107.380 83.410 107.700 ;
        RECT 83.670 106.000 83.810 114.180 ;
        RECT 84.130 111.780 84.270 118.260 ;
        RECT 84.530 115.880 84.790 116.200 ;
        RECT 84.590 112.120 84.730 115.880 ;
        RECT 84.990 115.540 85.250 115.860 ;
        RECT 85.050 114.160 85.190 115.540 ;
        RECT 84.990 113.840 85.250 114.160 ;
        RECT 84.530 111.800 84.790 112.120 ;
        RECT 84.070 111.460 84.330 111.780 ;
        RECT 83.610 105.680 83.870 106.000 ;
        RECT 85.050 105.320 85.190 113.840 ;
        RECT 84.990 105.000 85.250 105.320 ;
        RECT 81.770 104.660 82.030 104.980 ;
        RECT 81.830 103.280 81.970 104.660 ;
        RECT 80.850 102.960 81.110 103.280 ;
        RECT 81.770 102.960 82.030 103.280 ;
        RECT 80.910 100.220 81.050 102.960 ;
        RECT 85.050 100.560 85.190 105.000 ;
        RECT 85.510 102.260 85.650 118.940 ;
        RECT 85.970 105.660 86.110 121.320 ;
        RECT 86.430 120.280 86.570 126.420 ;
        RECT 86.830 124.720 87.090 125.040 ;
        RECT 86.370 119.960 86.630 120.280 ;
        RECT 86.370 116.450 86.630 116.540 ;
        RECT 86.890 116.450 87.030 124.720 ;
        RECT 87.810 124.700 87.950 130.500 ;
        RECT 89.650 127.420 89.790 137.640 ;
        RECT 90.510 137.300 90.770 137.620 ;
        RECT 90.970 137.300 91.230 137.620 ;
        RECT 90.570 134.900 90.710 137.300 ;
        RECT 90.510 134.580 90.770 134.900 ;
        RECT 91.030 132.860 91.170 137.300 ;
        RECT 90.970 132.540 91.230 132.860 ;
        RECT 89.590 127.100 89.850 127.420 ;
        RECT 88.670 126.760 88.930 127.080 ;
        RECT 88.730 125.040 88.870 126.760 ;
        RECT 89.650 125.040 89.790 127.100 ;
        RECT 93.330 125.800 93.470 137.980 ;
        RECT 94.650 137.300 94.910 137.620 ;
        RECT 93.730 134.580 93.990 134.900 ;
        RECT 93.790 133.200 93.930 134.580 ;
        RECT 93.730 132.880 93.990 133.200 ;
        RECT 94.710 132.180 94.850 137.300 ;
        RECT 94.650 131.860 94.910 132.180 ;
        RECT 93.330 125.660 93.930 125.800 ;
        RECT 88.670 124.720 88.930 125.040 ;
        RECT 89.590 124.720 89.850 125.040 ;
        RECT 87.750 124.380 88.010 124.700 ;
        RECT 93.270 124.380 93.530 124.700 ;
        RECT 91.890 122.680 92.150 123.000 ;
        RECT 88.670 122.340 88.930 122.660 ;
        RECT 88.210 120.980 88.470 121.300 ;
        RECT 87.750 118.600 88.010 118.920 ;
        RECT 86.370 116.310 87.030 116.450 ;
        RECT 86.370 116.220 86.630 116.310 ;
        RECT 86.890 114.160 87.030 116.310 ;
        RECT 86.830 113.840 87.090 114.160 ;
        RECT 86.370 113.500 86.630 113.820 ;
        RECT 87.810 113.560 87.950 118.600 ;
        RECT 88.270 114.160 88.410 120.980 ;
        RECT 88.730 117.560 88.870 122.340 ;
        RECT 90.050 119.960 90.310 120.280 ;
        RECT 89.130 119.280 89.390 119.600 ;
        RECT 88.670 117.240 88.930 117.560 ;
        RECT 89.190 115.860 89.330 119.280 ;
        RECT 89.590 116.220 89.850 116.540 ;
        RECT 89.130 115.540 89.390 115.860 ;
        RECT 88.210 113.840 88.470 114.160 ;
        RECT 86.430 112.120 86.570 113.500 ;
        RECT 86.890 113.480 87.950 113.560 ;
        RECT 86.830 113.420 87.950 113.480 ;
        RECT 86.830 113.160 87.090 113.420 ;
        RECT 86.370 111.800 86.630 112.120 ;
        RECT 86.370 107.720 86.630 108.040 ;
        RECT 86.430 105.660 86.570 107.720 ;
        RECT 87.810 106.000 87.950 113.420 ;
        RECT 89.190 110.760 89.330 115.540 ;
        RECT 89.650 111.100 89.790 116.220 ;
        RECT 90.110 115.860 90.250 119.960 ;
        RECT 91.950 119.600 92.090 122.680 ;
        RECT 93.330 122.320 93.470 124.380 ;
        RECT 93.270 122.000 93.530 122.320 ;
        RECT 93.790 119.600 93.930 125.660 ;
        RECT 91.890 119.510 92.150 119.600 ;
        RECT 91.890 119.370 93.010 119.510 ;
        RECT 91.890 119.280 92.150 119.370 ;
        RECT 90.050 115.540 90.310 115.860 ;
        RECT 89.590 110.780 89.850 111.100 ;
        RECT 89.130 110.440 89.390 110.760 ;
        RECT 89.650 108.120 89.790 110.780 ;
        RECT 90.510 110.440 90.770 110.760 ;
        RECT 89.190 107.980 89.790 108.120 ;
        RECT 87.750 105.680 88.010 106.000 ;
        RECT 85.910 105.340 86.170 105.660 ;
        RECT 86.370 105.340 86.630 105.660 ;
        RECT 85.970 103.620 86.110 105.340 ;
        RECT 87.290 104.660 87.550 104.980 ;
        RECT 85.910 103.300 86.170 103.620 ;
        RECT 85.450 101.940 85.710 102.260 ;
        RECT 84.990 100.240 85.250 100.560 ;
        RECT 80.850 99.900 81.110 100.220 ;
        RECT 85.970 99.960 86.110 103.300 ;
        RECT 87.350 102.260 87.490 104.660 ;
        RECT 87.810 103.960 87.950 105.680 ;
        RECT 87.750 103.640 88.010 103.960 ;
        RECT 87.290 101.940 87.550 102.260 ;
        RECT 87.750 101.940 88.010 102.260 ;
        RECT 82.690 99.560 82.950 99.880 ;
        RECT 85.970 99.820 87.030 99.960 ;
        RECT 82.750 97.840 82.890 99.560 ;
        RECT 85.910 97.860 86.170 98.180 ;
        RECT 82.690 97.520 82.950 97.840 ;
        RECT 85.970 95.800 86.110 97.860 ;
        RECT 85.910 95.480 86.170 95.800 ;
        RECT 86.890 95.120 87.030 99.820 ;
        RECT 87.350 95.120 87.490 101.940 ;
        RECT 87.810 95.460 87.950 101.940 ;
        RECT 89.190 99.540 89.330 107.980 ;
        RECT 89.590 107.380 89.850 107.700 ;
        RECT 89.650 103.960 89.790 107.380 ;
        RECT 90.570 106.080 90.710 110.440 ;
        RECT 91.890 110.100 92.150 110.420 ;
        RECT 90.110 105.940 91.630 106.080 ;
        RECT 90.110 105.320 90.250 105.940 ;
        RECT 90.510 105.340 90.770 105.660 ;
        RECT 90.050 105.000 90.310 105.320 ;
        RECT 89.590 103.640 89.850 103.960 ;
        RECT 90.050 103.640 90.310 103.960 ;
        RECT 89.590 99.560 89.850 99.880 ;
        RECT 89.130 99.220 89.390 99.540 ;
        RECT 89.650 95.800 89.790 99.560 ;
        RECT 90.110 98.035 90.250 103.640 ;
        RECT 90.570 101.240 90.710 105.340 ;
        RECT 90.510 100.920 90.770 101.240 ;
        RECT 91.490 98.520 91.630 105.940 ;
        RECT 91.430 98.200 91.690 98.520 ;
        RECT 90.040 97.665 90.320 98.035 ;
        RECT 90.110 97.160 90.250 97.665 ;
        RECT 90.050 96.840 90.310 97.160 ;
        RECT 89.590 95.480 89.850 95.800 ;
        RECT 87.750 95.140 88.010 95.460 ;
        RECT 86.830 94.800 87.090 95.120 ;
        RECT 87.290 94.800 87.550 95.120 ;
        RECT 91.950 94.780 92.090 110.100 ;
        RECT 92.870 105.660 93.010 119.370 ;
        RECT 93.730 119.280 93.990 119.600 ;
        RECT 93.790 117.220 93.930 119.280 ;
        RECT 95.110 118.940 95.370 119.260 ;
        RECT 95.170 117.560 95.310 118.940 ;
        RECT 95.110 117.240 95.370 117.560 ;
        RECT 93.730 116.900 93.990 117.220 ;
        RECT 95.570 116.900 95.830 117.220 ;
        RECT 95.110 116.560 95.370 116.880 ;
        RECT 93.730 115.540 93.990 115.860 ;
        RECT 93.790 113.140 93.930 115.540 ;
        RECT 94.650 114.180 94.910 114.500 ;
        RECT 93.730 112.820 93.990 113.140 ;
        RECT 93.790 111.100 93.930 112.820 ;
        RECT 93.730 110.780 93.990 111.100 ;
        RECT 93.790 109.400 93.930 110.780 ;
        RECT 94.710 109.480 94.850 114.180 ;
        RECT 95.170 113.140 95.310 116.560 ;
        RECT 95.630 114.160 95.770 116.900 ;
        RECT 95.570 113.840 95.830 114.160 ;
        RECT 95.110 112.820 95.370 113.140 ;
        RECT 93.730 109.080 93.990 109.400 ;
        RECT 94.710 109.340 95.310 109.480 ;
        RECT 94.650 107.380 94.910 107.700 ;
        RECT 94.190 106.360 94.450 106.680 ;
        RECT 92.810 105.340 93.070 105.660 ;
        RECT 92.810 103.640 93.070 103.960 ;
        RECT 92.870 102.940 93.010 103.640 ;
        RECT 93.730 102.960 93.990 103.280 ;
        RECT 92.810 102.620 93.070 102.940 ;
        RECT 92.350 100.920 92.610 101.240 ;
        RECT 92.410 97.500 92.550 100.920 ;
        RECT 93.790 100.900 93.930 102.960 ;
        RECT 93.730 100.580 93.990 100.900 ;
        RECT 93.270 99.560 93.530 99.880 ;
        RECT 92.800 97.665 93.080 98.035 ;
        RECT 93.330 97.840 93.470 99.560 ;
        RECT 94.250 99.540 94.390 106.360 ;
        RECT 94.190 99.220 94.450 99.540 ;
        RECT 92.810 97.520 93.070 97.665 ;
        RECT 93.270 97.520 93.530 97.840 ;
        RECT 94.180 97.665 94.460 98.035 ;
        RECT 94.710 97.840 94.850 107.380 ;
        RECT 95.170 102.940 95.310 109.340 ;
        RECT 96.090 105.660 96.230 159.060 ;
        RECT 96.550 157.000 96.690 190.000 ;
        RECT 97.010 184.200 97.150 190.000 ;
        RECT 97.470 184.280 97.610 211.760 ;
        RECT 98.330 210.740 98.590 211.060 ;
        RECT 98.390 209.020 98.530 210.740 ;
        RECT 98.850 209.700 98.990 211.760 ;
        RECT 99.710 211.080 99.970 211.400 ;
        RECT 98.790 209.380 99.050 209.700 ;
        RECT 99.770 209.020 99.910 211.080 ;
        RECT 100.690 210.040 100.830 213.800 ;
        RECT 102.930 211.420 103.190 211.740 ;
        RECT 100.630 209.720 100.890 210.040 ;
        RECT 98.330 208.700 98.590 209.020 ;
        RECT 99.710 208.700 99.970 209.020 ;
        RECT 97.870 204.280 98.130 204.600 ;
        RECT 97.930 197.800 98.070 204.280 ;
        RECT 99.250 202.920 99.510 203.240 ;
        RECT 99.310 201.880 99.450 202.920 ;
        RECT 101.550 202.580 101.810 202.900 ;
        RECT 99.250 201.560 99.510 201.880 ;
        RECT 99.250 200.880 99.510 201.200 ;
        RECT 98.330 199.860 98.590 200.180 ;
        RECT 98.390 198.140 98.530 199.860 ;
        RECT 98.330 197.820 98.590 198.140 ;
        RECT 98.790 197.820 99.050 198.140 ;
        RECT 99.310 197.880 99.450 200.880 ;
        RECT 99.710 200.540 99.970 200.860 ;
        RECT 99.770 198.820 99.910 200.540 ;
        RECT 99.710 198.500 99.970 198.820 ;
        RECT 100.170 198.160 100.430 198.480 ;
        RECT 101.080 198.305 101.360 198.675 ;
        RECT 100.230 197.880 100.370 198.160 ;
        RECT 101.150 198.140 101.290 198.305 ;
        RECT 97.870 197.480 98.130 197.800 ;
        RECT 98.850 196.440 98.990 197.820 ;
        RECT 99.310 197.740 100.370 197.880 ;
        RECT 101.090 197.820 101.350 198.140 ;
        RECT 101.610 197.800 101.750 202.580 ;
        RECT 102.990 201.880 103.130 211.420 ;
        RECT 103.450 208.680 103.590 213.800 ;
        RECT 104.370 212.080 104.510 216.180 ;
        RECT 106.670 212.080 106.810 216.520 ;
        RECT 107.070 213.800 107.330 214.120 ;
        RECT 107.130 212.760 107.270 213.800 ;
        RECT 107.070 212.440 107.330 212.760 ;
        RECT 104.310 211.760 104.570 212.080 ;
        RECT 106.610 211.760 106.870 212.080 ;
        RECT 103.390 208.360 103.650 208.680 ;
        RECT 102.930 201.560 103.190 201.880 ;
        RECT 102.460 201.025 102.740 201.395 ;
        RECT 102.470 200.880 102.730 201.025 ;
        RECT 102.930 197.820 103.190 198.140 ;
        RECT 98.790 196.120 99.050 196.440 ;
        RECT 98.330 195.440 98.590 195.760 ;
        RECT 98.790 195.670 99.050 195.760 ;
        RECT 99.310 195.670 99.450 197.740 ;
        RECT 100.630 197.480 100.890 197.800 ;
        RECT 101.550 197.480 101.810 197.800 ;
        RECT 100.170 197.140 100.430 197.460 ;
        RECT 98.790 195.530 99.450 195.670 ;
        RECT 98.790 195.440 99.050 195.530 ;
        RECT 97.870 189.660 98.130 189.980 ;
        RECT 97.930 188.280 98.070 189.660 ;
        RECT 97.870 187.960 98.130 188.280 ;
        RECT 98.390 184.880 98.530 195.440 ;
        RECT 99.710 193.400 99.970 193.720 ;
        RECT 99.770 187.600 99.910 193.400 ;
        RECT 100.230 189.980 100.370 197.140 ;
        RECT 100.690 196.350 100.830 197.480 ;
        RECT 102.010 197.140 102.270 197.460 ;
        RECT 102.470 197.140 102.730 197.460 ;
        RECT 101.090 196.350 101.350 196.440 ;
        RECT 100.690 196.210 101.350 196.350 ;
        RECT 100.690 195.420 100.830 196.210 ;
        RECT 101.090 196.120 101.350 196.210 ;
        RECT 102.070 195.760 102.210 197.140 ;
        RECT 102.530 196.100 102.670 197.140 ;
        RECT 102.470 195.780 102.730 196.100 ;
        RECT 101.550 195.440 101.810 195.760 ;
        RECT 102.010 195.440 102.270 195.760 ;
        RECT 100.630 195.100 100.890 195.420 ;
        RECT 101.610 193.720 101.750 195.440 ;
        RECT 102.990 193.720 103.130 197.820 ;
        RECT 101.550 193.400 101.810 193.720 ;
        RECT 102.930 193.400 103.190 193.720 ;
        RECT 101.610 193.020 101.750 193.400 ;
        RECT 103.450 193.040 103.590 208.360 ;
        RECT 106.150 202.920 106.410 203.240 ;
        RECT 103.850 202.580 104.110 202.900 ;
        RECT 103.910 201.540 104.050 202.580 ;
        RECT 103.850 201.220 104.110 201.540 ;
        RECT 106.210 201.200 106.350 202.920 ;
        RECT 106.150 200.880 106.410 201.200 ;
        RECT 107.130 200.860 107.270 212.440 ;
        RECT 107.990 209.040 108.250 209.360 ;
        RECT 108.050 206.640 108.190 209.040 ;
        RECT 107.990 206.320 108.250 206.640 ;
        RECT 108.050 204.000 108.190 206.320 ;
        RECT 108.450 205.980 108.710 206.300 ;
        RECT 107.590 203.860 108.190 204.000 ;
        RECT 107.590 201.880 107.730 203.860 ;
        RECT 107.990 203.260 108.250 203.580 ;
        RECT 107.530 201.560 107.790 201.880 ;
        RECT 103.850 200.540 104.110 200.860 ;
        RECT 104.770 200.540 105.030 200.860 ;
        RECT 105.230 200.540 105.490 200.860 ;
        RECT 107.070 200.540 107.330 200.860 ;
        RECT 103.910 196.440 104.050 200.540 ;
        RECT 104.830 199.160 104.970 200.540 ;
        RECT 104.770 198.840 105.030 199.160 ;
        RECT 105.290 197.995 105.430 200.540 ;
        RECT 106.610 199.860 106.870 200.180 ;
        RECT 105.680 198.305 105.960 198.675 ;
        RECT 105.750 198.140 105.890 198.305 ;
        RECT 106.670 198.140 106.810 199.860 ;
        RECT 107.530 198.160 107.790 198.480 ;
        RECT 105.220 197.625 105.500 197.995 ;
        RECT 105.690 197.820 105.950 198.140 ;
        RECT 106.610 197.820 106.870 198.140 ;
        RECT 105.230 197.140 105.490 197.460 ;
        RECT 105.290 196.440 105.430 197.140 ;
        RECT 103.850 196.120 104.110 196.440 ;
        RECT 105.230 196.120 105.490 196.440 ;
        RECT 106.670 195.420 106.810 197.820 ;
        RECT 106.610 195.100 106.870 195.420 ;
        RECT 107.590 193.040 107.730 198.160 ;
        RECT 108.050 195.760 108.190 203.260 ;
        RECT 108.510 202.900 108.650 205.980 ;
        RECT 114.890 202.920 115.150 203.240 ;
        RECT 108.450 202.580 108.710 202.900 ;
        RECT 108.510 198.820 108.650 202.580 ;
        RECT 114.950 201.880 115.090 202.920 ;
        RECT 114.890 201.560 115.150 201.880 ;
        RECT 120.870 200.880 121.130 201.200 ;
        RECT 108.450 198.500 108.710 198.820 ;
        RECT 117.190 197.820 117.450 198.140 ;
        RECT 110.290 197.140 110.550 197.460 ;
        RECT 110.350 196.100 110.490 197.140 ;
        RECT 110.290 195.780 110.550 196.100 ;
        RECT 107.990 195.440 108.250 195.760 ;
        RECT 108.050 193.040 108.190 195.440 ;
        RECT 117.250 194.740 117.390 197.820 ;
        RECT 118.110 197.480 118.370 197.800 ;
        RECT 117.190 194.420 117.450 194.740 ;
        RECT 118.170 193.720 118.310 197.480 ;
        RECT 120.930 196.440 121.070 200.880 ;
        RECT 124.550 197.820 124.810 198.140 ;
        RECT 125.010 197.820 125.270 198.140 ;
        RECT 122.250 197.140 122.510 197.460 ;
        RECT 120.870 196.120 121.130 196.440 ;
        RECT 120.870 195.100 121.130 195.420 ;
        RECT 114.890 193.400 115.150 193.720 ;
        RECT 118.110 193.400 118.370 193.720 ;
        RECT 101.610 192.880 102.210 193.020 ;
        RECT 102.070 190.320 102.210 192.880 ;
        RECT 103.390 192.720 103.650 193.040 ;
        RECT 107.530 192.720 107.790 193.040 ;
        RECT 107.990 192.720 108.250 193.040 ;
        RECT 102.010 190.000 102.270 190.320 ;
        RECT 100.170 189.660 100.430 189.980 ;
        RECT 103.450 189.640 103.590 192.720 ;
        RECT 106.610 191.700 106.870 192.020 ;
        RECT 106.670 191.000 106.810 191.700 ;
        RECT 106.610 190.680 106.870 191.000 ;
        RECT 107.590 189.980 107.730 192.720 ;
        RECT 108.050 190.660 108.190 192.720 ;
        RECT 108.450 192.040 108.710 192.360 ;
        RECT 108.510 191.000 108.650 192.040 ;
        RECT 108.450 190.680 108.710 191.000 ;
        RECT 111.670 190.680 111.930 191.000 ;
        RECT 107.990 190.340 108.250 190.660 ;
        RECT 107.530 189.660 107.790 189.980 ;
        RECT 103.390 189.320 103.650 189.640 ;
        RECT 102.470 188.980 102.730 189.300 ;
        RECT 102.530 187.600 102.670 188.980 ;
        RECT 103.450 187.600 103.590 189.320 ;
        RECT 99.710 187.280 99.970 187.600 ;
        RECT 102.470 187.280 102.730 187.600 ;
        RECT 103.390 187.280 103.650 187.600 ;
        RECT 99.770 184.880 99.910 187.280 ;
        RECT 101.090 186.940 101.350 187.260 ;
        RECT 110.290 186.940 110.550 187.260 ;
        RECT 110.750 186.940 111.010 187.260 ;
        RECT 98.330 184.560 98.590 184.880 ;
        RECT 99.710 184.560 99.970 184.880 ;
        RECT 96.950 183.880 97.210 184.200 ;
        RECT 97.470 184.140 98.070 184.280 ;
        RECT 97.410 183.540 97.670 183.860 ;
        RECT 97.470 180.120 97.610 183.540 ;
        RECT 97.410 179.800 97.670 180.120 ;
        RECT 96.950 179.120 97.210 179.440 ;
        RECT 97.010 177.400 97.150 179.120 ;
        RECT 96.950 177.080 97.210 177.400 ;
        RECT 96.950 169.940 97.210 170.260 ;
        RECT 97.010 168.900 97.150 169.940 ;
        RECT 96.950 168.580 97.210 168.900 ;
        RECT 97.010 165.840 97.150 168.580 ;
        RECT 97.930 166.520 98.070 184.140 ;
        RECT 98.390 182.840 98.530 184.560 ;
        RECT 98.330 182.520 98.590 182.840 ;
        RECT 101.150 182.160 101.290 186.940 ;
        RECT 107.530 186.260 107.790 186.580 ;
        RECT 108.450 186.260 108.710 186.580 ;
        RECT 105.230 184.220 105.490 184.540 ;
        RECT 102.930 183.540 103.190 183.860 ;
        RECT 102.990 182.160 103.130 183.540 ;
        RECT 98.330 181.840 98.590 182.160 ;
        RECT 101.090 181.840 101.350 182.160 ;
        RECT 102.930 181.840 103.190 182.160 ;
        RECT 98.390 179.100 98.530 181.840 ;
        RECT 100.630 179.120 100.890 179.440 ;
        RECT 105.290 179.220 105.430 184.220 ;
        RECT 105.690 183.540 105.950 183.860 ;
        RECT 105.750 181.820 105.890 183.540 ;
        RECT 105.690 181.500 105.950 181.820 ;
        RECT 106.610 181.500 106.870 181.820 ;
        RECT 98.330 178.780 98.590 179.100 ;
        RECT 99.710 176.060 99.970 176.380 ;
        RECT 99.770 174.000 99.910 176.060 ;
        RECT 100.170 174.360 100.430 174.680 ;
        RECT 98.790 173.680 99.050 174.000 ;
        RECT 99.710 173.680 99.970 174.000 ;
        RECT 98.850 171.960 98.990 173.680 ;
        RECT 98.790 171.640 99.050 171.960 ;
        RECT 98.850 168.560 98.990 171.640 ;
        RECT 99.770 168.755 99.910 173.680 ;
        RECT 98.790 168.240 99.050 168.560 ;
        RECT 99.250 168.240 99.510 168.560 ;
        RECT 99.700 168.385 99.980 168.755 ;
        RECT 100.230 168.560 100.370 174.360 ;
        RECT 100.690 170.940 100.830 179.120 ;
        RECT 104.370 179.080 105.430 179.220 ;
        RECT 103.850 176.400 104.110 176.720 ;
        RECT 103.390 175.720 103.650 176.040 ;
        RECT 101.090 170.960 101.350 171.280 ;
        RECT 100.630 170.620 100.890 170.940 ;
        RECT 100.630 168.920 100.890 169.240 ;
        RECT 99.710 168.240 99.970 168.385 ;
        RECT 100.170 168.240 100.430 168.560 ;
        RECT 99.310 167.540 99.450 168.240 ;
        RECT 100.690 167.880 100.830 168.920 ;
        RECT 100.630 167.560 100.890 167.880 ;
        RECT 99.250 167.220 99.510 167.540 ;
        RECT 97.870 166.200 98.130 166.520 ;
        RECT 96.950 165.520 97.210 165.840 ;
        RECT 97.410 165.180 97.670 165.500 ;
        RECT 97.470 160.740 97.610 165.180 ;
        RECT 101.150 163.120 101.290 170.960 ;
        RECT 102.930 170.620 103.190 170.940 ;
        RECT 102.990 169.240 103.130 170.620 ;
        RECT 102.930 168.920 103.190 169.240 ;
        RECT 101.090 162.800 101.350 163.120 ;
        RECT 101.150 161.080 101.290 162.800 ;
        RECT 101.090 160.760 101.350 161.080 ;
        RECT 97.410 160.420 97.670 160.740 ;
        RECT 97.870 159.740 98.130 160.060 ;
        RECT 97.410 159.060 97.670 159.380 ;
        RECT 97.470 157.340 97.610 159.060 ;
        RECT 97.930 157.340 98.070 159.740 ;
        RECT 98.330 157.360 98.590 157.680 ;
        RECT 101.090 157.360 101.350 157.680 ;
        RECT 102.930 157.360 103.190 157.680 ;
        RECT 97.410 157.020 97.670 157.340 ;
        RECT 97.870 157.020 98.130 157.340 ;
        RECT 96.490 156.680 96.750 157.000 ;
        RECT 97.470 154.620 97.610 157.020 ;
        RECT 97.410 154.300 97.670 154.620 ;
        RECT 98.390 153.940 98.530 157.360 ;
        RECT 98.330 153.620 98.590 153.940 ;
        RECT 98.390 152.240 98.530 153.620 ;
        RECT 101.150 152.240 101.290 157.360 ;
        RECT 96.950 151.920 97.210 152.240 ;
        RECT 98.330 151.920 98.590 152.240 ;
        RECT 101.090 151.920 101.350 152.240 ;
        RECT 97.010 144.760 97.150 151.920 ;
        RECT 101.150 150.200 101.290 151.920 ;
        RECT 101.090 149.880 101.350 150.200 ;
        RECT 102.470 149.540 102.730 149.860 ;
        RECT 98.790 148.860 99.050 149.180 ;
        RECT 98.850 146.800 98.990 148.860 ;
        RECT 101.550 148.180 101.810 148.500 ;
        RECT 101.610 147.140 101.750 148.180 ;
        RECT 101.550 146.820 101.810 147.140 ;
        RECT 97.410 146.480 97.670 146.800 ;
        RECT 98.790 146.480 99.050 146.800 ;
        RECT 99.710 146.480 99.970 146.800 ;
        RECT 96.950 144.440 97.210 144.760 ;
        RECT 96.490 126.420 96.750 126.740 ;
        RECT 96.550 125.380 96.690 126.420 ;
        RECT 96.490 125.060 96.750 125.380 ;
        RECT 96.490 118.260 96.750 118.580 ;
        RECT 96.550 114.070 96.690 118.260 ;
        RECT 97.470 114.840 97.610 146.480 ;
        RECT 98.850 143.740 98.990 146.480 ;
        RECT 99.770 144.420 99.910 146.480 ;
        RECT 102.530 144.760 102.670 149.540 ;
        RECT 102.990 149.180 103.130 157.360 ;
        RECT 102.930 148.860 103.190 149.180 ;
        RECT 102.470 144.440 102.730 144.760 ;
        RECT 99.710 144.160 99.970 144.420 ;
        RECT 99.710 144.100 100.370 144.160 ;
        RECT 99.770 144.020 100.370 144.100 ;
        RECT 98.790 143.420 99.050 143.740 ;
        RECT 99.710 143.420 99.970 143.740 ;
        RECT 98.850 138.980 98.990 143.420 ;
        RECT 98.790 138.660 99.050 138.980 ;
        RECT 98.790 132.540 99.050 132.860 ;
        RECT 98.330 131.860 98.590 132.180 ;
        RECT 98.390 127.080 98.530 131.860 ;
        RECT 98.850 130.140 98.990 132.540 ;
        RECT 98.790 129.820 99.050 130.140 ;
        RECT 98.330 126.760 98.590 127.080 ;
        RECT 99.250 126.420 99.510 126.740 ;
        RECT 99.310 121.980 99.450 126.420 ;
        RECT 99.250 121.660 99.510 121.980 ;
        RECT 97.410 114.520 97.670 114.840 ;
        RECT 97.410 114.070 97.670 114.160 ;
        RECT 96.550 113.930 97.670 114.070 ;
        RECT 97.410 113.840 97.670 113.930 ;
        RECT 96.490 111.120 96.750 111.440 ;
        RECT 96.030 105.340 96.290 105.660 ;
        RECT 95.110 102.620 95.370 102.940 ;
        RECT 95.170 100.560 95.310 102.620 ;
        RECT 95.110 100.240 95.370 100.560 ;
        RECT 95.570 100.130 95.830 100.220 ;
        RECT 96.090 100.130 96.230 105.340 ;
        RECT 96.550 104.980 96.690 111.120 ;
        RECT 97.470 110.760 97.610 113.840 ;
        RECT 98.330 112.820 98.590 113.140 ;
        RECT 98.390 111.440 98.530 112.820 ;
        RECT 98.330 111.120 98.590 111.440 ;
        RECT 97.410 110.440 97.670 110.760 ;
        RECT 99.770 105.320 99.910 143.420 ;
        RECT 100.230 138.640 100.370 144.020 ;
        RECT 101.550 143.420 101.810 143.740 ;
        RECT 100.170 138.320 100.430 138.640 ;
        RECT 101.610 128.100 101.750 143.420 ;
        RECT 102.470 140.930 102.730 141.020 ;
        RECT 103.450 140.930 103.590 175.720 ;
        RECT 103.910 174.340 104.050 176.400 ;
        RECT 104.370 175.700 104.510 179.080 ;
        RECT 105.230 176.060 105.490 176.380 ;
        RECT 105.750 176.120 105.890 181.500 ;
        RECT 106.670 177.400 106.810 181.500 ;
        RECT 107.070 178.100 107.330 178.420 ;
        RECT 107.590 178.275 107.730 186.260 ;
        RECT 107.990 184.560 108.250 184.880 ;
        RECT 108.050 182.160 108.190 184.560 ;
        RECT 107.990 181.840 108.250 182.160 ;
        RECT 108.050 179.440 108.190 181.840 ;
        RECT 108.510 180.120 108.650 186.260 ;
        RECT 110.350 185.560 110.490 186.940 ;
        RECT 110.290 185.240 110.550 185.560 ;
        RECT 110.290 184.560 110.550 184.880 ;
        RECT 108.450 179.800 108.710 180.120 ;
        RECT 107.990 179.120 108.250 179.440 ;
        RECT 106.610 177.080 106.870 177.400 ;
        RECT 107.130 177.310 107.270 178.100 ;
        RECT 107.520 177.905 107.800 178.275 ;
        RECT 108.050 177.595 108.190 179.120 ;
        RECT 107.530 177.310 107.790 177.400 ;
        RECT 107.130 177.170 107.790 177.310 ;
        RECT 107.980 177.225 108.260 177.595 ;
        RECT 107.530 177.080 107.790 177.170 ;
        RECT 107.990 176.800 108.250 177.060 ;
        RECT 107.590 176.740 108.250 176.800 ;
        RECT 107.590 176.660 108.190 176.740 ;
        RECT 104.310 175.380 104.570 175.700 ;
        RECT 105.290 175.555 105.430 176.060 ;
        RECT 105.750 175.980 105.935 176.120 ;
        RECT 105.795 175.950 105.935 175.980 ;
        RECT 105.795 175.810 106.350 175.950 ;
        RECT 105.220 175.185 105.500 175.555 ;
        RECT 105.230 174.360 105.490 174.680 ;
        RECT 103.850 174.020 104.110 174.340 ;
        RECT 105.290 169.240 105.430 174.360 ;
        RECT 106.210 173.400 106.350 175.810 ;
        RECT 107.590 175.700 107.730 176.660 ;
        RECT 108.450 176.400 108.710 176.720 ;
        RECT 107.980 175.865 108.260 176.235 ;
        RECT 107.530 175.380 107.790 175.700 ;
        RECT 108.050 174.000 108.190 175.865 ;
        RECT 108.510 174.340 108.650 176.400 ;
        RECT 110.350 175.555 110.490 184.560 ;
        RECT 110.810 180.120 110.950 186.940 ;
        RECT 111.210 184.560 111.470 184.880 ;
        RECT 110.750 179.800 111.010 180.120 ;
        RECT 111.270 177.400 111.410 184.560 ;
        RECT 111.210 177.080 111.470 177.400 ;
        RECT 110.750 175.720 111.010 176.040 ;
        RECT 110.280 175.185 110.560 175.555 ;
        RECT 108.450 174.020 108.710 174.340 ;
        RECT 107.990 173.680 108.250 174.000 ;
        RECT 110.350 173.660 110.490 175.185 ;
        RECT 106.210 173.260 106.810 173.400 ;
        RECT 110.290 173.340 110.550 173.660 ;
        RECT 106.150 172.660 106.410 172.980 ;
        RECT 105.230 168.920 105.490 169.240 ;
        RECT 106.210 168.900 106.350 172.660 ;
        RECT 106.670 169.240 106.810 173.260 ;
        RECT 108.450 172.660 108.710 172.980 ;
        RECT 107.070 171.300 107.330 171.620 ;
        RECT 106.610 168.920 106.870 169.240 ;
        RECT 106.150 168.580 106.410 168.900 ;
        RECT 106.670 168.560 106.810 168.920 ;
        RECT 107.130 168.560 107.270 171.300 ;
        RECT 108.510 168.560 108.650 172.660 ;
        RECT 110.350 172.320 110.490 173.340 ;
        RECT 109.890 172.180 110.490 172.320 ;
        RECT 109.890 170.260 110.030 172.180 ;
        RECT 110.290 171.640 110.550 171.960 ;
        RECT 109.830 169.940 110.090 170.260 ;
        RECT 110.350 168.560 110.490 171.640 ;
        RECT 106.610 168.240 106.870 168.560 ;
        RECT 107.070 168.240 107.330 168.560 ;
        RECT 108.450 168.240 108.710 168.560 ;
        RECT 110.290 168.240 110.550 168.560 ;
        RECT 109.830 165.180 110.090 165.500 ;
        RECT 109.890 163.800 110.030 165.180 ;
        RECT 109.830 163.480 110.090 163.800 ;
        RECT 107.980 160.905 108.260 161.275 ;
        RECT 107.990 160.760 108.250 160.905 ;
        RECT 109.890 160.740 110.030 163.480 ;
        RECT 109.830 160.420 110.090 160.740 ;
        RECT 110.810 160.400 110.950 175.720 ;
        RECT 111.270 174.340 111.410 177.080 ;
        RECT 111.210 174.020 111.470 174.340 ;
        RECT 110.750 160.080 111.010 160.400 ;
        RECT 104.310 159.400 104.570 159.720 ;
        RECT 108.450 159.400 108.710 159.720 ;
        RECT 104.370 158.360 104.510 159.400 ;
        RECT 104.310 158.040 104.570 158.360 ;
        RECT 107.990 157.700 108.250 158.020 ;
        RECT 106.150 157.360 106.410 157.680 ;
        RECT 103.850 156.340 104.110 156.660 ;
        RECT 103.910 152.580 104.050 156.340 ;
        RECT 106.210 155.640 106.350 157.360 ;
        RECT 108.050 155.640 108.190 157.700 ;
        RECT 108.510 157.340 108.650 159.400 ;
        RECT 108.450 157.020 108.710 157.340 ;
        RECT 111.730 155.640 111.870 190.680 ;
        RECT 114.950 190.320 115.090 193.400 ;
        RECT 120.930 193.040 121.070 195.100 ;
        RECT 120.870 192.720 121.130 193.040 ;
        RECT 118.570 192.380 118.830 192.700 ;
        RECT 116.270 191.700 116.530 192.020 ;
        RECT 116.330 191.000 116.470 191.700 ;
        RECT 118.630 191.000 118.770 192.380 ;
        RECT 119.950 191.700 120.210 192.020 ;
        RECT 116.270 190.680 116.530 191.000 ;
        RECT 118.570 190.680 118.830 191.000 ;
        RECT 114.890 190.000 115.150 190.320 ;
        RECT 117.190 190.000 117.450 190.320 ;
        RECT 116.270 189.320 116.530 189.640 ;
        RECT 115.810 186.600 116.070 186.920 ;
        RECT 112.130 186.260 112.390 186.580 ;
        RECT 112.190 176.720 112.330 186.260 ;
        RECT 113.970 185.240 114.230 185.560 ;
        RECT 114.030 181.140 114.170 185.240 ;
        RECT 115.350 183.880 115.610 184.200 ;
        RECT 115.410 182.840 115.550 183.880 ;
        RECT 115.350 182.520 115.610 182.840 ;
        RECT 114.430 181.500 114.690 181.820 ;
        RECT 113.970 180.820 114.230 181.140 ;
        RECT 114.030 177.060 114.170 180.820 ;
        RECT 113.970 176.740 114.230 177.060 ;
        RECT 112.130 176.400 112.390 176.720 ;
        RECT 114.490 175.700 114.630 181.500 ;
        RECT 114.890 179.800 115.150 180.120 ;
        RECT 114.950 176.380 115.090 179.800 ;
        RECT 115.410 179.440 115.550 182.520 ;
        RECT 115.350 179.120 115.610 179.440 ;
        RECT 114.890 176.060 115.150 176.380 ;
        RECT 114.430 175.380 114.690 175.700 ;
        RECT 113.050 173.680 113.310 174.000 ;
        RECT 112.590 173.340 112.850 173.660 ;
        RECT 112.650 171.960 112.790 173.340 ;
        RECT 113.110 171.960 113.250 173.680 ;
        RECT 114.950 173.660 115.090 176.060 ;
        RECT 115.350 174.020 115.610 174.340 ;
        RECT 114.890 173.340 115.150 173.660 ;
        RECT 112.590 171.640 112.850 171.960 ;
        RECT 113.050 171.640 113.310 171.960 ;
        RECT 112.650 171.280 112.790 171.640 ;
        RECT 112.590 170.960 112.850 171.280 ;
        RECT 113.110 168.560 113.250 171.640 ;
        RECT 114.950 171.620 115.090 173.340 ;
        RECT 114.890 171.300 115.150 171.620 ;
        RECT 115.410 170.940 115.550 174.020 ;
        RECT 115.350 170.620 115.610 170.940 ;
        RECT 113.050 168.240 113.310 168.560 ;
        RECT 115.410 168.220 115.550 170.620 ;
        RECT 115.870 169.240 116.010 186.600 ;
        RECT 116.330 176.040 116.470 189.320 ;
        RECT 116.270 175.720 116.530 176.040 ;
        RECT 115.810 168.920 116.070 169.240 ;
        RECT 115.350 167.900 115.610 168.220 ;
        RECT 113.510 167.560 113.770 167.880 ;
        RECT 113.570 166.520 113.710 167.560 ;
        RECT 115.810 167.220 116.070 167.540 ;
        RECT 113.510 166.200 113.770 166.520 ;
        RECT 112.580 165.665 112.860 166.035 ;
        RECT 112.650 163.460 112.790 165.665 ;
        RECT 115.870 165.500 116.010 167.220 ;
        RECT 115.810 165.180 116.070 165.500 ;
        RECT 116.270 164.840 116.530 165.160 ;
        RECT 113.970 164.500 114.230 164.820 ;
        RECT 116.330 164.675 116.470 164.840 ;
        RECT 112.590 163.140 112.850 163.460 ;
        RECT 114.030 163.120 114.170 164.500 ;
        RECT 116.260 164.305 116.540 164.675 ;
        RECT 117.250 163.200 117.390 190.000 ;
        RECT 118.630 188.280 118.770 190.680 ;
        RECT 118.570 187.960 118.830 188.280 ;
        RECT 117.650 179.120 117.910 179.440 ;
        RECT 118.560 179.265 118.840 179.635 ;
        RECT 118.570 179.120 118.830 179.265 ;
        RECT 117.710 176.720 117.850 179.120 ;
        RECT 118.110 178.440 118.370 178.760 ;
        RECT 117.650 176.400 117.910 176.720 ;
        RECT 117.710 174.340 117.850 176.400 ;
        RECT 118.170 176.120 118.310 178.440 ;
        RECT 118.630 177.060 118.770 179.120 ;
        RECT 119.480 178.585 119.760 178.955 ;
        RECT 119.550 177.400 119.690 178.585 ;
        RECT 119.490 177.080 119.750 177.400 ;
        RECT 118.570 176.740 118.830 177.060 ;
        RECT 118.570 176.120 118.830 176.380 ;
        RECT 118.170 176.060 118.830 176.120 ;
        RECT 119.030 176.060 119.290 176.380 ;
        RECT 118.170 175.980 118.770 176.060 ;
        RECT 117.650 174.020 117.910 174.340 ;
        RECT 117.650 173.340 117.910 173.660 ;
        RECT 117.710 166.180 117.850 173.340 ;
        RECT 118.110 172.660 118.370 172.980 ;
        RECT 118.170 170.940 118.310 172.660 ;
        RECT 118.630 171.360 118.770 175.980 ;
        RECT 119.090 171.960 119.230 176.060 ;
        RECT 119.030 171.640 119.290 171.960 ;
        RECT 119.490 171.640 119.750 171.960 ;
        RECT 119.550 171.360 119.690 171.640 ;
        RECT 118.630 171.220 119.690 171.360 ;
        RECT 118.110 170.620 118.370 170.940 ;
        RECT 118.170 169.240 118.310 170.620 ;
        RECT 118.630 170.260 118.770 171.220 ;
        RECT 118.570 169.940 118.830 170.260 ;
        RECT 118.110 168.920 118.370 169.240 ;
        RECT 118.630 168.560 118.770 169.940 ;
        RECT 118.570 168.240 118.830 168.560 ;
        RECT 119.030 168.240 119.290 168.560 ;
        RECT 118.110 167.220 118.370 167.540 ;
        RECT 117.650 165.860 117.910 166.180 ;
        RECT 117.650 165.180 117.910 165.500 ;
        RECT 117.710 163.800 117.850 165.180 ;
        RECT 117.650 163.480 117.910 163.800 ;
        RECT 113.970 162.800 114.230 163.120 ;
        RECT 116.270 162.800 116.530 163.120 ;
        RECT 117.250 163.060 117.850 163.200 ;
        RECT 115.810 162.460 116.070 162.780 ;
        RECT 116.330 162.635 116.470 162.800 ;
        RECT 112.130 162.120 112.390 162.440 ;
        RECT 112.190 160.060 112.330 162.120 ;
        RECT 115.350 161.780 115.610 162.100 ;
        RECT 112.590 160.080 112.850 160.400 ;
        RECT 112.130 159.740 112.390 160.060 ;
        RECT 106.150 155.320 106.410 155.640 ;
        RECT 107.990 155.320 108.250 155.640 ;
        RECT 111.670 155.320 111.930 155.640 ;
        RECT 112.130 154.300 112.390 154.620 ;
        RECT 112.190 152.580 112.330 154.300 ;
        RECT 103.850 152.260 104.110 152.580 ;
        RECT 112.130 152.260 112.390 152.580 ;
        RECT 102.470 140.790 103.590 140.930 ;
        RECT 102.470 140.700 102.730 140.790 ;
        RECT 102.530 136.600 102.670 140.700 ;
        RECT 103.910 140.680 104.050 152.260 ;
        RECT 104.770 151.920 105.030 152.240 ;
        RECT 104.830 147.480 104.970 151.920 ;
        RECT 112.190 151.900 112.330 152.260 ;
        RECT 109.370 151.580 109.630 151.900 ;
        RECT 112.130 151.580 112.390 151.900 ;
        RECT 106.150 149.540 106.410 149.860 ;
        RECT 104.770 147.160 105.030 147.480 ;
        RECT 105.690 147.160 105.950 147.480 ;
        RECT 105.750 146.800 105.890 147.160 ;
        RECT 105.690 146.480 105.950 146.800 ;
        RECT 105.750 144.080 105.890 146.480 ;
        RECT 106.210 144.760 106.350 149.540 ;
        RECT 106.610 148.180 106.870 148.500 ;
        RECT 106.670 147.140 106.810 148.180 ;
        RECT 106.610 146.820 106.870 147.140 ;
        RECT 109.430 146.800 109.570 151.580 ;
        RECT 109.370 146.480 109.630 146.800 ;
        RECT 106.150 144.440 106.410 144.760 ;
        RECT 105.690 143.760 105.950 144.080 ;
        RECT 105.230 141.720 105.490 142.040 ;
        RECT 104.310 141.380 104.570 141.700 ;
        RECT 103.850 140.360 104.110 140.680 ;
        RECT 103.910 139.320 104.050 140.360 ;
        RECT 103.850 139.000 104.110 139.320 ;
        RECT 103.390 138.660 103.650 138.980 ;
        RECT 102.470 136.280 102.730 136.600 ;
        RECT 103.450 133.200 103.590 138.660 ;
        RECT 104.370 138.300 104.510 141.380 ;
        RECT 104.310 137.980 104.570 138.300 ;
        RECT 104.370 133.200 104.510 137.980 ;
        RECT 104.770 137.300 105.030 137.620 ;
        RECT 104.830 136.260 104.970 137.300 ;
        RECT 104.770 135.940 105.030 136.260 ;
        RECT 103.390 132.880 103.650 133.200 ;
        RECT 104.310 132.880 104.570 133.200 ;
        RECT 103.450 131.160 103.590 132.880 ;
        RECT 103.390 130.840 103.650 131.160 ;
        RECT 102.470 129.140 102.730 129.460 ;
        RECT 101.550 127.780 101.810 128.100 ;
        RECT 102.530 127.080 102.670 129.140 ;
        RECT 103.450 127.760 103.590 130.840 ;
        RECT 104.370 130.820 104.510 132.880 ;
        RECT 104.310 130.500 104.570 130.820 ;
        RECT 103.390 127.440 103.650 127.760 ;
        RECT 102.010 126.760 102.270 127.080 ;
        RECT 102.470 126.760 102.730 127.080 ;
        RECT 102.070 125.720 102.210 126.760 ;
        RECT 103.850 126.420 104.110 126.740 ;
        RECT 102.010 125.400 102.270 125.720 ;
        RECT 101.550 123.700 101.810 124.020 ;
        RECT 101.610 120.280 101.750 123.700 ;
        RECT 102.070 121.980 102.210 125.400 ;
        RECT 103.910 125.040 104.050 126.420 ;
        RECT 104.370 125.380 104.510 130.500 ;
        RECT 104.310 125.060 104.570 125.380 ;
        RECT 103.850 124.720 104.110 125.040 ;
        RECT 103.910 121.980 104.050 124.720 ;
        RECT 104.370 121.980 104.510 125.060 ;
        RECT 102.010 121.660 102.270 121.980 ;
        RECT 103.850 121.660 104.110 121.980 ;
        RECT 104.310 121.660 104.570 121.980 ;
        RECT 101.550 119.960 101.810 120.280 ;
        RECT 102.070 119.680 102.210 121.660 ;
        RECT 102.070 119.600 102.670 119.680 ;
        RECT 103.910 119.600 104.050 121.660 ;
        RECT 104.370 119.940 104.510 121.660 ;
        RECT 105.290 120.280 105.430 141.720 ;
        RECT 109.370 141.040 109.630 141.360 ;
        RECT 107.070 140.020 107.330 140.340 ;
        RECT 108.450 140.020 108.710 140.340 ;
        RECT 107.130 138.640 107.270 140.020 ;
        RECT 107.070 138.320 107.330 138.640 ;
        RECT 105.690 137.980 105.950 138.300 ;
        RECT 105.750 123.000 105.890 137.980 ;
        RECT 108.510 136.260 108.650 140.020 ;
        RECT 108.450 135.940 108.710 136.260 ;
        RECT 107.070 130.840 107.330 131.160 ;
        RECT 107.130 130.480 107.270 130.840 ;
        RECT 109.430 130.820 109.570 141.040 ;
        RECT 110.290 140.700 110.550 141.020 ;
        RECT 110.350 139.320 110.490 140.700 ;
        RECT 110.290 139.000 110.550 139.320 ;
        RECT 112.650 138.640 112.790 160.080 ;
        RECT 115.410 160.060 115.550 161.780 ;
        RECT 115.870 161.080 116.010 162.460 ;
        RECT 116.260 162.265 116.540 162.635 ;
        RECT 115.810 160.760 116.070 161.080 ;
        RECT 116.730 160.420 116.990 160.740 ;
        RECT 115.350 159.740 115.610 160.060 ;
        RECT 114.890 158.040 115.150 158.360 ;
        RECT 114.950 157.340 115.090 158.040 ;
        RECT 115.410 157.680 115.550 159.740 ;
        RECT 115.350 157.360 115.610 157.680 ;
        RECT 114.890 157.020 115.150 157.340 ;
        RECT 115.410 157.080 115.550 157.360 ;
        RECT 115.410 156.940 116.010 157.080 ;
        RECT 115.870 156.660 116.010 156.940 ;
        RECT 114.890 156.340 115.150 156.660 ;
        RECT 115.350 156.340 115.610 156.660 ;
        RECT 115.810 156.340 116.070 156.660 ;
        RECT 114.950 155.300 115.090 156.340 ;
        RECT 114.890 154.980 115.150 155.300 ;
        RECT 115.410 154.620 115.550 156.340 ;
        RECT 116.790 154.960 116.930 160.420 ;
        RECT 117.190 159.060 117.450 159.380 ;
        RECT 117.250 157.680 117.390 159.060 ;
        RECT 117.190 157.360 117.450 157.680 ;
        RECT 117.190 156.680 117.450 157.000 ;
        RECT 116.730 154.640 116.990 154.960 ;
        RECT 115.350 154.300 115.610 154.620 ;
        RECT 115.810 153.620 116.070 153.940 ;
        RECT 115.870 151.755 116.010 153.620 ;
        RECT 117.250 152.240 117.390 156.680 ;
        RECT 117.190 151.920 117.450 152.240 ;
        RECT 115.800 151.385 116.080 151.755 ;
        RECT 114.890 143.760 115.150 144.080 ;
        RECT 113.970 142.740 114.230 143.060 ;
        RECT 113.510 141.040 113.770 141.360 ;
        RECT 112.590 138.320 112.850 138.640 ;
        RECT 111.670 137.980 111.930 138.300 ;
        RECT 111.730 136.260 111.870 137.980 ;
        RECT 112.650 136.600 112.790 138.320 ;
        RECT 112.590 136.280 112.850 136.600 ;
        RECT 111.670 135.940 111.930 136.260 ;
        RECT 111.730 132.860 111.870 135.940 ;
        RECT 113.570 133.880 113.710 141.040 ;
        RECT 113.510 133.560 113.770 133.880 ;
        RECT 111.670 132.540 111.930 132.860 ;
        RECT 109.370 130.500 109.630 130.820 ;
        RECT 106.610 130.160 106.870 130.480 ;
        RECT 107.070 130.160 107.330 130.480 ;
        RECT 107.990 130.160 108.250 130.480 ;
        RECT 111.200 130.305 111.480 130.675 ;
        RECT 111.730 130.480 111.870 132.540 ;
        RECT 105.690 122.680 105.950 123.000 ;
        RECT 105.230 119.960 105.490 120.280 ;
        RECT 104.310 119.620 104.570 119.940 ;
        RECT 105.290 119.680 105.430 119.960 ;
        RECT 101.550 119.280 101.810 119.600 ;
        RECT 102.070 119.540 102.730 119.600 ;
        RECT 102.470 119.280 102.730 119.540 ;
        RECT 103.850 119.280 104.110 119.600 ;
        RECT 100.630 116.220 100.890 116.540 ;
        RECT 101.090 116.220 101.350 116.540 ;
        RECT 100.690 113.480 100.830 116.220 ;
        RECT 101.150 114.840 101.290 116.220 ;
        RECT 101.610 114.840 101.750 119.280 ;
        RECT 104.370 118.920 104.510 119.620 ;
        RECT 104.830 119.540 105.430 119.680 ;
        RECT 104.310 118.600 104.570 118.920 ;
        RECT 104.830 116.540 104.970 119.540 ;
        RECT 105.230 118.940 105.490 119.260 ;
        RECT 106.150 118.940 106.410 119.260 ;
        RECT 104.770 116.220 105.030 116.540 ;
        RECT 103.390 115.540 103.650 115.860 ;
        RECT 101.090 114.520 101.350 114.840 ;
        RECT 101.550 114.520 101.810 114.840 ;
        RECT 101.610 114.160 101.750 114.520 ;
        RECT 101.550 113.840 101.810 114.160 ;
        RECT 102.930 113.840 103.190 114.160 ;
        RECT 100.630 113.160 100.890 113.480 ;
        RECT 102.990 112.120 103.130 113.840 ;
        RECT 102.930 111.800 103.190 112.120 ;
        RECT 103.450 111.780 103.590 115.540 ;
        RECT 105.290 114.160 105.430 118.940 ;
        RECT 106.210 117.560 106.350 118.940 ;
        RECT 106.150 117.240 106.410 117.560 ;
        RECT 105.230 113.840 105.490 114.160 ;
        RECT 103.390 111.460 103.650 111.780 ;
        RECT 101.090 111.120 101.350 111.440 ;
        RECT 99.710 105.000 99.970 105.320 ;
        RECT 96.490 104.660 96.750 104.980 ;
        RECT 99.250 104.660 99.510 104.980 ;
        RECT 95.570 99.990 96.230 100.130 ;
        RECT 95.570 99.900 95.830 99.990 ;
        RECT 99.310 97.840 99.450 104.660 ;
        RECT 101.150 103.280 101.290 111.120 ;
        RECT 103.850 108.060 104.110 108.380 ;
        RECT 103.390 105.680 103.650 106.000 ;
        RECT 102.010 104.660 102.270 104.980 ;
        RECT 101.090 102.960 101.350 103.280 ;
        RECT 92.350 97.240 92.610 97.500 ;
        RECT 93.730 97.240 93.990 97.500 ;
        RECT 92.350 97.180 93.990 97.240 ;
        RECT 92.410 97.100 93.930 97.180 ;
        RECT 94.250 94.780 94.390 97.665 ;
        RECT 94.650 97.520 94.910 97.840 ;
        RECT 99.250 97.520 99.510 97.840 ;
        RECT 97.410 97.180 97.670 97.500 ;
        RECT 100.630 97.410 100.890 97.500 ;
        RECT 101.150 97.410 101.290 102.960 ;
        RECT 101.550 99.560 101.810 99.880 ;
        RECT 101.610 98.520 101.750 99.560 ;
        RECT 101.550 98.200 101.810 98.520 ;
        RECT 100.630 97.270 101.290 97.410 ;
        RECT 100.630 97.180 100.890 97.270 ;
        RECT 95.110 96.500 95.370 96.820 ;
        RECT 95.170 95.460 95.310 96.500 ;
        RECT 95.110 95.140 95.370 95.460 ;
        RECT 95.570 95.140 95.830 95.460 ;
        RECT 71.190 94.460 71.450 94.780 ;
        RECT 73.490 94.460 73.750 94.780 ;
        RECT 77.630 94.460 77.890 94.780 ;
        RECT 78.090 94.460 78.350 94.780 ;
        RECT 79.930 94.460 80.190 94.780 ;
        RECT 91.890 94.460 92.150 94.780 ;
        RECT 94.190 94.460 94.450 94.780 ;
        RECT 89.130 94.120 89.390 94.440 ;
        RECT 92.350 94.120 92.610 94.440 ;
        RECT 73.030 93.780 73.290 94.100 ;
        RECT 76.250 93.780 76.510 94.100 ;
        RECT 79.470 93.780 79.730 94.100 ;
        RECT 82.690 93.780 82.950 94.100 ;
        RECT 85.910 93.780 86.170 94.100 ;
        RECT 73.090 86.550 73.230 93.780 ;
        RECT 76.310 86.550 76.450 93.780 ;
        RECT 79.530 86.550 79.670 93.780 ;
        RECT 82.750 86.550 82.890 93.780 ;
        RECT 85.970 86.550 86.110 93.780 ;
        RECT 89.190 86.550 89.330 94.120 ;
        RECT 92.410 86.550 92.550 94.120 ;
        RECT 95.630 86.550 95.770 95.140 ;
        RECT 97.470 94.780 97.610 97.180 ;
        RECT 102.070 97.160 102.210 104.660 ;
        RECT 103.450 103.960 103.590 105.680 ;
        RECT 103.910 105.320 104.050 108.060 ;
        RECT 103.850 105.000 104.110 105.320 ;
        RECT 103.910 103.960 104.050 105.000 ;
        RECT 104.310 104.660 104.570 104.980 ;
        RECT 103.390 103.640 103.650 103.960 ;
        RECT 103.850 103.640 104.110 103.960 ;
        RECT 102.930 101.940 103.190 102.260 ;
        RECT 102.990 100.560 103.130 101.940 ;
        RECT 104.370 101.240 104.510 104.660 ;
        RECT 104.310 100.920 104.570 101.240 ;
        RECT 102.930 100.240 103.190 100.560 ;
        RECT 102.010 96.840 102.270 97.160 ;
        RECT 102.990 94.780 103.130 100.240 ;
        RECT 104.370 100.220 104.510 100.920 ;
        RECT 105.290 100.900 105.430 113.840 ;
        RECT 105.690 105.680 105.950 106.000 ;
        RECT 105.750 103.280 105.890 105.680 ;
        RECT 105.690 102.960 105.950 103.280 ;
        RECT 106.670 101.240 106.810 130.160 ;
        RECT 107.130 124.440 107.270 130.160 ;
        RECT 108.050 129.460 108.190 130.160 ;
        RECT 111.270 130.140 111.410 130.305 ;
        RECT 111.670 130.160 111.930 130.480 ;
        RECT 112.130 130.160 112.390 130.480 ;
        RECT 111.210 129.820 111.470 130.140 ;
        RECT 107.990 129.140 108.250 129.460 ;
        RECT 108.050 127.760 108.190 129.140 ;
        RECT 112.190 128.440 112.330 130.160 ;
        RECT 112.130 128.120 112.390 128.440 ;
        RECT 107.990 127.440 108.250 127.760 ;
        RECT 108.910 126.760 109.170 127.080 ;
        RECT 113.500 126.905 113.780 127.275 ;
        RECT 113.510 126.760 113.770 126.905 ;
        RECT 108.440 124.440 108.720 124.555 ;
        RECT 107.130 124.300 108.720 124.440 ;
        RECT 108.440 124.185 108.720 124.300 ;
        RECT 108.510 122.320 108.650 124.185 ;
        RECT 108.450 122.000 108.710 122.320 ;
        RECT 108.970 119.940 109.110 126.760 ;
        RECT 113.570 122.400 113.710 126.760 ;
        RECT 114.030 124.440 114.170 142.740 ;
        RECT 114.430 137.870 114.690 137.960 ;
        RECT 114.950 137.870 115.090 143.760 ;
        RECT 114.430 137.730 115.090 137.870 ;
        RECT 114.430 137.640 114.690 137.730 ;
        RECT 114.950 127.760 115.090 137.730 ;
        RECT 115.350 134.920 115.610 135.240 ;
        RECT 115.410 133.880 115.550 134.920 ;
        RECT 115.350 133.560 115.610 133.880 ;
        RECT 115.410 127.760 115.550 133.560 ;
        RECT 114.890 127.440 115.150 127.760 ;
        RECT 115.350 127.440 115.610 127.760 ;
        RECT 114.950 125.040 115.090 127.440 ;
        RECT 115.870 125.720 116.010 151.385 ;
        RECT 117.710 146.800 117.850 163.060 ;
        RECT 118.170 157.680 118.310 167.220 ;
        RECT 118.630 166.180 118.770 168.240 ;
        RECT 118.570 165.860 118.830 166.180 ;
        RECT 119.090 166.035 119.230 168.240 ;
        RECT 119.020 165.665 119.300 166.035 ;
        RECT 118.570 165.180 118.830 165.500 ;
        RECT 118.630 163.120 118.770 165.180 ;
        RECT 119.030 164.500 119.290 164.820 ;
        RECT 118.570 162.800 118.830 163.120 ;
        RECT 118.630 161.080 118.770 162.800 ;
        RECT 118.570 160.760 118.830 161.080 ;
        RECT 119.090 160.595 119.230 164.500 ;
        RECT 119.490 163.140 119.750 163.460 ;
        RECT 119.020 160.225 119.300 160.595 ;
        RECT 119.550 160.060 119.690 163.140 ;
        RECT 119.490 159.740 119.750 160.060 ;
        RECT 118.110 157.360 118.370 157.680 ;
        RECT 118.570 157.360 118.830 157.680 ;
        RECT 118.170 156.660 118.310 157.360 ;
        RECT 118.110 156.340 118.370 156.660 ;
        RECT 118.170 154.280 118.310 156.340 ;
        RECT 118.110 153.960 118.370 154.280 ;
        RECT 118.630 149.860 118.770 157.360 ;
        RECT 119.490 157.020 119.750 157.340 ;
        RECT 119.550 155.640 119.690 157.020 ;
        RECT 119.490 155.320 119.750 155.640 ;
        RECT 119.030 154.300 119.290 154.620 ;
        RECT 119.090 152.920 119.230 154.300 ;
        RECT 119.030 152.600 119.290 152.920 ;
        RECT 118.570 149.540 118.830 149.860 ;
        RECT 119.490 148.860 119.750 149.180 ;
        RECT 117.650 146.480 117.910 146.800 ;
        RECT 116.270 145.460 116.530 145.780 ;
        RECT 117.650 145.460 117.910 145.780 ;
        RECT 116.330 143.400 116.470 145.460 ;
        RECT 116.270 143.080 116.530 143.400 ;
        RECT 117.710 141.360 117.850 145.460 ;
        RECT 117.650 141.040 117.910 141.360 ;
        RECT 118.570 140.360 118.830 140.680 ;
        RECT 116.730 137.640 116.990 137.960 ;
        RECT 116.790 136.600 116.930 137.640 ;
        RECT 116.730 136.280 116.990 136.600 ;
        RECT 118.630 135.920 118.770 140.360 ;
        RECT 117.650 135.600 117.910 135.920 ;
        RECT 118.570 135.600 118.830 135.920 ;
        RECT 117.710 128.440 117.850 135.600 ;
        RECT 118.630 133.200 118.770 135.600 ;
        RECT 119.550 134.900 119.690 148.860 ;
        RECT 120.010 139.320 120.150 191.700 ;
        RECT 120.930 189.640 121.070 192.720 ;
        RECT 120.870 189.320 121.130 189.640 ;
        RECT 122.310 187.260 122.450 197.140 ;
        RECT 123.630 195.780 123.890 196.100 ;
        RECT 123.690 190.660 123.830 195.780 ;
        RECT 123.630 190.340 123.890 190.660 ;
        RECT 123.690 187.600 123.830 190.340 ;
        RECT 124.090 190.000 124.350 190.320 ;
        RECT 124.150 188.280 124.290 190.000 ;
        RECT 124.090 187.960 124.350 188.280 ;
        RECT 123.630 187.280 123.890 187.600 ;
        RECT 122.250 186.940 122.510 187.260 ;
        RECT 123.630 184.220 123.890 184.540 ;
        RECT 123.690 182.840 123.830 184.220 ;
        RECT 123.630 182.520 123.890 182.840 ;
        RECT 123.630 181.500 123.890 181.820 ;
        RECT 123.690 176.915 123.830 181.500 ;
        RECT 124.090 180.820 124.350 181.140 ;
        RECT 120.400 176.545 120.680 176.915 ;
        RECT 123.620 176.545 123.900 176.915 ;
        RECT 124.150 176.720 124.290 180.820 ;
        RECT 120.470 171.620 120.610 176.545 ;
        RECT 124.090 176.400 124.350 176.720 ;
        RECT 121.790 175.720 122.050 176.040 ;
        RECT 121.850 174.340 121.990 175.720 ;
        RECT 122.710 175.380 122.970 175.700 ;
        RECT 121.790 174.020 122.050 174.340 ;
        RECT 120.410 171.530 120.670 171.620 ;
        RECT 120.410 171.390 121.530 171.530 ;
        RECT 120.410 171.300 120.670 171.390 ;
        RECT 120.410 170.620 120.670 170.940 ;
        RECT 121.390 170.680 121.530 171.390 ;
        RECT 121.850 171.360 121.990 174.020 ;
        RECT 121.850 171.220 122.450 171.360 ;
        RECT 122.310 170.940 122.450 171.220 ;
        RECT 120.470 168.560 120.610 170.620 ;
        RECT 121.390 170.540 121.990 170.680 ;
        RECT 122.250 170.620 122.510 170.940 ;
        RECT 121.330 169.940 121.590 170.260 ;
        RECT 120.410 168.240 120.670 168.560 ;
        RECT 120.470 165.500 120.610 168.240 ;
        RECT 121.390 167.960 121.530 169.940 ;
        RECT 120.930 167.820 121.530 167.960 ;
        RECT 120.410 165.180 120.670 165.500 ;
        RECT 120.400 162.265 120.680 162.635 ;
        RECT 120.470 157.680 120.610 162.265 ;
        RECT 120.410 157.360 120.670 157.680 ;
        RECT 120.930 155.300 121.070 167.820 ;
        RECT 121.330 167.395 121.590 167.540 ;
        RECT 121.320 167.025 121.600 167.395 ;
        RECT 121.390 163.120 121.530 167.025 ;
        RECT 121.330 162.800 121.590 163.120 ;
        RECT 121.390 162.440 121.530 162.800 ;
        RECT 121.330 162.120 121.590 162.440 ;
        RECT 121.390 157.875 121.530 162.120 ;
        RECT 121.850 160.060 121.990 170.540 ;
        RECT 122.250 162.800 122.510 163.120 ;
        RECT 121.790 159.740 122.050 160.060 ;
        RECT 122.310 159.235 122.450 162.800 ;
        RECT 122.770 161.840 122.910 175.380 ;
        RECT 123.630 174.360 123.890 174.680 ;
        RECT 123.170 173.680 123.430 174.000 ;
        RECT 123.230 170.260 123.370 173.680 ;
        RECT 123.690 171.620 123.830 174.360 ;
        RECT 124.150 172.980 124.290 176.400 ;
        RECT 124.610 175.700 124.750 197.820 ;
        RECT 125.070 193.720 125.210 197.820 ;
        RECT 126.850 197.480 127.110 197.800 ;
        RECT 125.470 195.440 125.730 195.760 ;
        RECT 125.010 193.400 125.270 193.720 ;
        RECT 125.530 193.020 125.670 195.440 ;
        RECT 125.070 192.880 125.670 193.020 ;
        RECT 124.550 175.380 124.810 175.700 ;
        RECT 124.090 172.660 124.350 172.980 ;
        RECT 123.630 171.300 123.890 171.620 ;
        RECT 123.170 169.940 123.430 170.260 ;
        RECT 123.230 168.900 123.370 169.940 ;
        RECT 123.170 168.580 123.430 168.900 ;
        RECT 123.690 167.540 123.830 171.300 ;
        RECT 124.080 171.105 124.360 171.475 ;
        RECT 124.610 171.280 124.750 175.380 ;
        RECT 124.150 170.940 124.290 171.105 ;
        RECT 124.550 170.960 124.810 171.280 ;
        RECT 124.090 170.620 124.350 170.940 ;
        RECT 124.610 168.220 124.750 170.960 ;
        RECT 124.550 167.900 124.810 168.220 ;
        RECT 123.630 167.220 123.890 167.540 ;
        RECT 124.090 166.200 124.350 166.520 ;
        RECT 123.630 165.180 123.890 165.500 ;
        RECT 123.690 163.120 123.830 165.180 ;
        RECT 123.630 162.800 123.890 163.120 ;
        RECT 123.690 162.100 123.830 162.800 ;
        RECT 122.770 161.700 123.370 161.840 ;
        RECT 123.630 161.780 123.890 162.100 ;
        RECT 122.240 158.865 122.520 159.235 ;
        RECT 122.710 159.060 122.970 159.380 ;
        RECT 121.320 157.505 121.600 157.875 ;
        RECT 122.770 157.760 122.910 159.060 ;
        RECT 123.230 158.360 123.370 161.700 ;
        RECT 124.150 160.400 124.290 166.200 ;
        RECT 124.610 165.160 124.750 167.900 ;
        RECT 124.550 164.840 124.810 165.160 ;
        RECT 124.550 161.780 124.810 162.100 ;
        RECT 124.090 160.080 124.350 160.400 ;
        RECT 124.150 159.380 124.290 160.080 ;
        RECT 124.090 159.060 124.350 159.380 ;
        RECT 123.170 158.040 123.430 158.360 ;
        RECT 122.310 157.620 122.910 157.760 ;
        RECT 123.230 157.760 123.370 158.040 ;
        RECT 123.230 157.680 124.290 157.760 ;
        RECT 123.230 157.620 124.350 157.680 ;
        RECT 120.870 154.980 121.130 155.300 ;
        RECT 120.930 154.360 121.070 154.980 ;
        RECT 120.470 154.220 121.070 154.360 ;
        RECT 120.470 151.900 120.610 154.220 ;
        RECT 120.870 153.620 121.130 153.940 ;
        RECT 120.410 151.580 120.670 151.900 ;
        RECT 120.410 146.480 120.670 146.800 ;
        RECT 120.470 142.040 120.610 146.480 ;
        RECT 120.410 141.720 120.670 142.040 ;
        RECT 119.950 139.000 120.210 139.320 ;
        RECT 120.930 138.980 121.070 153.620 ;
        RECT 121.390 152.240 121.530 157.505 ;
        RECT 122.310 156.660 122.450 157.620 ;
        RECT 124.090 157.360 124.350 157.620 ;
        RECT 122.710 156.680 122.970 157.000 ;
        RECT 122.250 156.340 122.510 156.660 ;
        RECT 121.330 151.920 121.590 152.240 ;
        RECT 122.250 151.920 122.510 152.240 ;
        RECT 121.390 149.180 121.530 151.920 ;
        RECT 121.330 148.860 121.590 149.180 ;
        RECT 121.790 148.860 122.050 149.180 ;
        RECT 121.850 143.740 121.990 148.860 ;
        RECT 121.790 143.420 122.050 143.740 ;
        RECT 122.310 143.060 122.450 151.920 ;
        RECT 122.770 149.520 122.910 156.680 ;
        RECT 124.090 156.340 124.350 156.660 ;
        RECT 124.150 155.300 124.290 156.340 ;
        RECT 124.090 154.980 124.350 155.300 ;
        RECT 123.630 152.150 123.890 152.240 ;
        RECT 124.610 152.150 124.750 161.780 ;
        RECT 123.630 152.010 124.750 152.150 ;
        RECT 123.630 151.920 123.890 152.010 ;
        RECT 122.710 149.200 122.970 149.520 ;
        RECT 123.170 149.090 123.430 149.180 ;
        RECT 123.690 149.090 123.830 151.920 ;
        RECT 124.090 149.090 124.350 149.180 ;
        RECT 123.170 148.950 124.350 149.090 ;
        RECT 123.170 148.860 123.430 148.950 ;
        RECT 124.090 148.860 124.350 148.950 ;
        RECT 124.550 144.720 124.810 144.760 ;
        RECT 125.070 144.720 125.210 192.880 ;
        RECT 126.910 188.280 127.050 197.480 ;
        RECT 131.910 197.140 132.170 197.460 ;
        RECT 127.310 196.120 127.570 196.440 ;
        RECT 127.370 193.040 127.510 196.120 ;
        RECT 131.970 193.720 132.110 197.140 ;
        RECT 132.370 195.440 132.630 195.760 ;
        RECT 134.210 195.440 134.470 195.760 ;
        RECT 132.430 193.720 132.570 195.440 ;
        RECT 132.830 194.760 133.090 195.080 ;
        RECT 131.910 193.400 132.170 193.720 ;
        RECT 132.370 193.400 132.630 193.720 ;
        RECT 127.310 192.720 127.570 193.040 ;
        RECT 132.370 192.720 132.630 193.040 ;
        RECT 130.990 192.380 131.250 192.700 ;
        RECT 127.770 191.700 128.030 192.020 ;
        RECT 130.070 191.700 130.330 192.020 ;
        RECT 127.830 191.000 127.970 191.700 ;
        RECT 127.770 190.680 128.030 191.000 ;
        RECT 128.690 190.340 128.950 190.660 ;
        RECT 128.230 188.980 128.490 189.300 ;
        RECT 126.850 187.960 127.110 188.280 ;
        RECT 126.390 187.620 126.650 187.940 ;
        RECT 125.470 186.600 125.730 186.920 ;
        RECT 125.930 186.600 126.190 186.920 ;
        RECT 125.530 181.480 125.670 186.600 ;
        RECT 125.990 185.560 126.130 186.600 ;
        RECT 125.930 185.240 126.190 185.560 ;
        RECT 126.450 185.220 126.590 187.620 ;
        RECT 127.310 187.280 127.570 187.600 ;
        RECT 126.390 184.900 126.650 185.220 ;
        RECT 125.470 181.160 125.730 181.480 ;
        RECT 126.450 181.140 126.590 184.900 ;
        RECT 126.850 183.540 127.110 183.860 ;
        RECT 126.390 180.820 126.650 181.140 ;
        RECT 126.450 180.120 126.590 180.820 ;
        RECT 126.390 179.800 126.650 180.120 ;
        RECT 126.390 179.120 126.650 179.440 ;
        RECT 125.920 177.225 126.200 177.595 ;
        RECT 125.930 177.080 126.190 177.225 ;
        RECT 125.470 176.740 125.730 177.060 ;
        RECT 125.530 176.380 125.670 176.740 ;
        RECT 125.470 176.060 125.730 176.380 ;
        RECT 125.530 174.340 125.670 176.060 ;
        RECT 126.450 174.680 126.590 179.120 ;
        RECT 126.910 176.040 127.050 183.540 ;
        RECT 126.850 175.720 127.110 176.040 ;
        RECT 126.390 174.360 126.650 174.680 ;
        RECT 127.370 174.340 127.510 187.280 ;
        RECT 128.290 187.260 128.430 188.980 ;
        RECT 128.750 187.680 128.890 190.340 ;
        RECT 128.750 187.540 129.350 187.680 ;
        RECT 129.610 187.620 129.870 187.940 ;
        RECT 128.230 186.940 128.490 187.260 ;
        RECT 127.770 186.600 128.030 186.920 ;
        RECT 127.830 183.860 127.970 186.600 ;
        RECT 128.750 184.960 128.890 187.540 ;
        RECT 129.210 187.260 129.350 187.540 ;
        RECT 129.670 187.260 129.810 187.620 ;
        RECT 129.150 186.940 129.410 187.260 ;
        RECT 129.610 186.940 129.870 187.260 ;
        RECT 129.150 186.260 129.410 186.580 ;
        RECT 129.210 185.220 129.350 186.260 ;
        RECT 129.610 185.240 129.870 185.560 ;
        RECT 128.290 184.820 128.890 184.960 ;
        RECT 129.150 184.900 129.410 185.220 ;
        RECT 128.290 184.540 128.430 184.820 ;
        RECT 128.230 184.220 128.490 184.540 ;
        RECT 127.770 183.540 128.030 183.860 ;
        RECT 127.830 177.480 127.970 183.540 ;
        RECT 129.210 182.840 129.350 184.900 ;
        RECT 129.150 182.520 129.410 182.840 ;
        RECT 128.230 181.500 128.490 181.820 ;
        RECT 128.290 181.140 128.430 181.500 ;
        RECT 128.680 181.305 128.960 181.675 ;
        RECT 128.750 181.140 128.890 181.305 ;
        RECT 128.230 180.820 128.490 181.140 ;
        RECT 128.690 180.820 128.950 181.140 ;
        RECT 128.290 179.440 128.430 180.820 ;
        RECT 128.750 179.520 128.890 180.820 ;
        RECT 129.210 180.120 129.350 182.520 ;
        RECT 129.670 180.120 129.810 185.240 ;
        RECT 130.130 184.200 130.270 191.700 ;
        RECT 130.530 186.600 130.790 186.920 ;
        RECT 130.590 184.540 130.730 186.600 ;
        RECT 130.530 184.220 130.790 184.540 ;
        RECT 130.070 183.880 130.330 184.200 ;
        RECT 129.150 179.800 129.410 180.120 ;
        RECT 129.610 179.800 129.870 180.120 ;
        RECT 128.230 179.120 128.490 179.440 ;
        RECT 128.750 179.380 129.350 179.520 ;
        RECT 127.830 177.340 128.430 177.480 ;
        RECT 127.770 176.740 128.030 177.060 ;
        RECT 127.830 176.380 127.970 176.740 ;
        RECT 127.770 176.060 128.030 176.380 ;
        RECT 128.290 176.120 128.430 177.340 ;
        RECT 125.470 174.020 125.730 174.340 ;
        RECT 127.310 174.020 127.570 174.340 ;
        RECT 125.930 173.340 126.190 173.660 ;
        RECT 125.990 169.240 126.130 173.340 ;
        RECT 127.370 170.680 127.510 174.020 ;
        RECT 127.830 171.475 127.970 176.060 ;
        RECT 128.290 175.980 128.890 176.120 ;
        RECT 128.750 175.700 128.890 175.980 ;
        RECT 128.230 175.380 128.490 175.700 ;
        RECT 128.690 175.380 128.950 175.700 ;
        RECT 127.760 171.105 128.040 171.475 ;
        RECT 128.290 171.280 128.430 175.380 ;
        RECT 129.210 174.760 129.350 179.380 ;
        RECT 130.130 179.220 130.270 183.880 ;
        RECT 130.590 180.995 130.730 184.220 ;
        RECT 130.520 180.625 130.800 180.995 ;
        RECT 130.590 179.780 130.730 180.625 ;
        RECT 130.530 179.460 130.790 179.780 ;
        RECT 130.130 179.080 130.730 179.220 ;
        RECT 129.610 178.440 129.870 178.760 ;
        RECT 130.070 178.440 130.330 178.760 ;
        RECT 129.670 178.275 129.810 178.440 ;
        RECT 129.600 177.905 129.880 178.275 ;
        RECT 130.130 177.400 130.270 178.440 ;
        RECT 130.070 177.080 130.330 177.400 ;
        RECT 130.070 175.720 130.330 176.040 ;
        RECT 129.210 174.620 129.810 174.760 ;
        RECT 129.150 173.680 129.410 174.000 ;
        RECT 128.690 172.660 128.950 172.980 ;
        RECT 128.750 171.620 128.890 172.660 ;
        RECT 128.690 171.300 128.950 171.620 ;
        RECT 127.770 170.960 128.030 171.105 ;
        RECT 128.230 170.960 128.490 171.280 ;
        RECT 126.910 170.600 127.510 170.680 ;
        RECT 126.850 170.540 127.510 170.600 ;
        RECT 126.850 170.280 127.110 170.540 ;
        RECT 127.770 170.280 128.030 170.600 ;
        RECT 125.930 168.920 126.190 169.240 ;
        RECT 127.830 166.520 127.970 170.280 ;
        RECT 129.210 170.260 129.350 173.680 ;
        RECT 129.150 169.940 129.410 170.260 ;
        RECT 128.690 168.470 128.950 168.560 ;
        RECT 129.210 168.470 129.350 169.940 ;
        RECT 128.690 168.330 129.350 168.470 ;
        RECT 128.690 168.240 128.950 168.330 ;
        RECT 129.150 167.560 129.410 167.880 ;
        RECT 127.770 166.200 128.030 166.520 ;
        RECT 125.920 165.665 126.200 166.035 ;
        RECT 125.990 160.400 126.130 165.665 ;
        RECT 127.770 165.520 128.030 165.840 ;
        RECT 127.830 163.460 127.970 165.520 ;
        RECT 128.690 165.410 128.950 165.500 ;
        RECT 129.210 165.410 129.350 167.560 ;
        RECT 129.670 165.840 129.810 174.620 ;
        RECT 130.130 173.320 130.270 175.720 ;
        RECT 130.590 174.340 130.730 179.080 ;
        RECT 131.050 178.955 131.190 192.380 ;
        RECT 131.910 190.000 132.170 190.320 ;
        RECT 131.450 187.620 131.710 187.940 ;
        RECT 131.510 184.880 131.650 187.620 ;
        RECT 131.970 187.260 132.110 190.000 ;
        RECT 131.910 186.940 132.170 187.260 ;
        RECT 131.970 185.560 132.110 186.940 ;
        RECT 132.430 186.920 132.570 192.720 ;
        RECT 132.890 188.280 133.030 194.760 ;
        RECT 133.750 192.380 134.010 192.700 ;
        RECT 133.810 191.000 133.950 192.380 ;
        RECT 134.270 191.000 134.410 195.440 ;
        RECT 133.750 190.680 134.010 191.000 ;
        RECT 134.210 190.680 134.470 191.000 ;
        RECT 132.830 187.960 133.090 188.280 ;
        RECT 132.370 186.600 132.630 186.920 ;
        RECT 131.910 185.240 132.170 185.560 ;
        RECT 131.970 185.075 132.110 185.240 ;
        RECT 131.450 184.560 131.710 184.880 ;
        RECT 131.900 184.705 132.180 185.075 ;
        RECT 131.510 179.100 131.650 184.560 ;
        RECT 132.430 184.200 132.570 186.600 ;
        RECT 132.890 185.560 133.030 187.960 ;
        RECT 132.830 185.240 133.090 185.560 ;
        RECT 132.890 184.880 133.950 184.960 ;
        RECT 132.890 184.820 134.010 184.880 ;
        RECT 132.370 183.880 132.630 184.200 ;
        RECT 131.910 183.540 132.170 183.860 ;
        RECT 131.970 181.820 132.110 183.540 ;
        RECT 131.910 181.500 132.170 181.820 ;
        RECT 132.430 180.880 132.570 183.880 ;
        RECT 132.890 181.140 133.030 184.820 ;
        RECT 133.750 184.560 134.010 184.820 ;
        RECT 133.290 184.220 133.550 184.540 ;
        RECT 134.270 184.280 134.410 190.680 ;
        RECT 140.650 190.000 140.910 190.320 ;
        RECT 137.430 188.980 137.690 189.300 ;
        RECT 137.490 187.260 137.630 188.980 ;
        RECT 140.710 188.280 140.850 190.000 ;
        RECT 140.650 187.960 140.910 188.280 ;
        RECT 137.430 186.940 137.690 187.260 ;
        RECT 142.030 186.940 142.290 187.260 ;
        RECT 143.870 186.940 144.130 187.260 ;
        RECT 135.590 186.600 135.850 186.920 ;
        RECT 135.650 185.560 135.790 186.600 ;
        RECT 135.590 185.240 135.850 185.560 ;
        RECT 134.660 184.705 134.940 185.075 ;
        RECT 137.490 184.880 137.630 186.940 ;
        RECT 140.650 186.260 140.910 186.580 ;
        RECT 134.670 184.560 134.930 184.705 ;
        RECT 136.510 184.560 136.770 184.880 ;
        RECT 137.430 184.560 137.690 184.880 ;
        RECT 137.890 184.560 138.150 184.880 ;
        RECT 138.810 184.560 139.070 184.880 ;
        RECT 133.350 182.500 133.490 184.220 ;
        RECT 134.270 184.140 134.870 184.280 ;
        RECT 133.290 182.180 133.550 182.500 ;
        RECT 133.290 181.500 133.550 181.820 ;
        RECT 133.750 181.500 134.010 181.820 ;
        RECT 134.210 181.500 134.470 181.820 ;
        RECT 131.970 180.740 132.570 180.880 ;
        RECT 132.830 180.820 133.090 181.140 ;
        RECT 130.980 178.585 131.260 178.955 ;
        RECT 131.450 178.780 131.710 179.100 ;
        RECT 130.990 178.100 131.250 178.420 ;
        RECT 131.050 177.060 131.190 178.100 ;
        RECT 130.990 176.740 131.250 177.060 ;
        RECT 131.450 176.060 131.710 176.380 ;
        RECT 130.530 174.020 130.790 174.340 ;
        RECT 130.980 173.825 131.260 174.195 ;
        RECT 130.990 173.680 131.250 173.825 ;
        RECT 130.070 173.000 130.330 173.320 ;
        RECT 130.130 170.940 130.270 173.000 ;
        RECT 130.990 171.300 131.250 171.620 ;
        RECT 130.070 170.620 130.330 170.940 ;
        RECT 130.130 168.560 130.270 170.620 ;
        RECT 131.050 170.260 131.190 171.300 ;
        RECT 130.530 169.940 130.790 170.260 ;
        RECT 130.990 169.940 131.250 170.260 ;
        RECT 130.070 168.240 130.330 168.560 ;
        RECT 130.130 167.540 130.270 168.240 ;
        RECT 130.070 167.220 130.330 167.540 ;
        RECT 129.610 165.520 129.870 165.840 ;
        RECT 130.590 165.500 130.730 169.940 ;
        RECT 128.690 165.270 129.350 165.410 ;
        RECT 128.690 165.180 128.950 165.270 ;
        RECT 130.530 165.180 130.790 165.500 ;
        RECT 130.990 165.180 131.250 165.500 ;
        RECT 128.230 164.840 128.490 165.160 ;
        RECT 129.610 164.840 129.870 165.160 ;
        RECT 127.770 163.140 128.030 163.460 ;
        RECT 127.770 162.460 128.030 162.780 ;
        RECT 127.830 161.080 127.970 162.460 ;
        RECT 127.770 160.760 128.030 161.080 ;
        RECT 126.390 160.480 126.650 160.740 ;
        RECT 128.290 160.480 128.430 164.840 ;
        RECT 128.690 164.560 128.950 164.820 ;
        RECT 128.690 164.500 129.350 164.560 ;
        RECT 128.750 164.420 129.350 164.500 ;
        RECT 126.390 160.420 128.430 160.480 ;
        RECT 125.930 160.080 126.190 160.400 ;
        RECT 126.450 160.340 128.430 160.420 ;
        RECT 125.470 159.400 125.730 159.720 ;
        RECT 125.530 157.680 125.670 159.400 ;
        RECT 125.470 157.360 125.730 157.680 ;
        RECT 125.530 154.360 125.670 157.360 ;
        RECT 125.990 157.340 126.130 160.080 ;
        RECT 126.390 159.740 126.650 160.060 ;
        RECT 127.770 159.740 128.030 160.060 ;
        RECT 125.930 157.020 126.190 157.340 ;
        RECT 126.450 154.960 126.590 159.740 ;
        RECT 127.830 159.380 127.970 159.740 ;
        RECT 127.770 159.060 128.030 159.380 ;
        RECT 128.290 157.680 128.430 160.340 ;
        RECT 128.230 157.360 128.490 157.680 ;
        RECT 127.310 157.020 127.570 157.340 ;
        RECT 126.390 154.640 126.650 154.960 ;
        RECT 125.530 154.220 126.130 154.360 ;
        RECT 125.470 153.620 125.730 153.940 ;
        RECT 125.530 152.240 125.670 153.620 ;
        RECT 125.470 151.920 125.730 152.240 ;
        RECT 125.990 149.180 126.130 154.220 ;
        RECT 126.850 153.620 127.110 153.940 ;
        RECT 126.910 150.200 127.050 153.620 ;
        RECT 127.370 152.920 127.510 157.020 ;
        RECT 127.310 152.600 127.570 152.920 ;
        RECT 126.850 149.880 127.110 150.200 ;
        RECT 128.690 149.200 128.950 149.520 ;
        RECT 125.930 148.860 126.190 149.180 ;
        RECT 128.750 147.140 128.890 149.200 ;
        RECT 128.690 146.820 128.950 147.140 ;
        RECT 129.210 146.800 129.350 164.420 ;
        RECT 129.670 163.800 129.810 164.840 ;
        RECT 129.610 163.480 129.870 163.800 ;
        RECT 130.520 162.945 130.800 163.315 ;
        RECT 130.590 162.440 130.730 162.945 ;
        RECT 131.050 162.635 131.190 165.180 ;
        RECT 130.530 162.120 130.790 162.440 ;
        RECT 130.980 162.265 131.260 162.635 ;
        RECT 131.050 160.400 131.190 162.265 ;
        RECT 130.990 160.080 131.250 160.400 ;
        RECT 131.510 160.060 131.650 176.060 ;
        RECT 131.970 173.515 132.110 180.740 ;
        RECT 132.890 179.440 133.030 180.820 ;
        RECT 133.350 180.120 133.490 181.500 ;
        RECT 133.290 179.800 133.550 180.120 ;
        RECT 133.350 179.635 133.490 179.800 ;
        RECT 132.830 179.120 133.090 179.440 ;
        RECT 133.280 179.265 133.560 179.635 ;
        RECT 133.810 179.440 133.950 181.500 ;
        RECT 134.270 179.440 134.410 181.500 ;
        RECT 134.730 179.440 134.870 184.140 ;
        RECT 135.590 183.880 135.850 184.200 ;
        RECT 135.650 181.820 135.790 183.880 ;
        RECT 136.570 183.860 136.710 184.560 ;
        RECT 136.050 183.540 136.310 183.860 ;
        RECT 136.510 183.540 136.770 183.860 ;
        RECT 136.110 182.500 136.250 183.540 ;
        RECT 136.050 182.180 136.310 182.500 ;
        RECT 135.590 181.500 135.850 181.820 ;
        RECT 132.370 178.440 132.630 178.760 ;
        RECT 132.830 178.440 133.090 178.760 ;
        RECT 132.430 178.275 132.570 178.440 ;
        RECT 132.360 177.905 132.640 178.275 ;
        RECT 131.900 173.145 132.180 173.515 ;
        RECT 131.910 172.660 132.170 172.980 ;
        RECT 131.970 168.560 132.110 172.660 ;
        RECT 132.430 171.960 132.570 177.905 ;
        RECT 132.890 176.915 133.030 178.440 ;
        RECT 132.820 176.545 133.100 176.915 ;
        RECT 132.890 176.040 133.030 176.545 ;
        RECT 132.830 175.720 133.090 176.040 ;
        RECT 133.350 174.195 133.490 179.265 ;
        RECT 133.750 179.120 134.010 179.440 ;
        RECT 134.210 179.120 134.470 179.440 ;
        RECT 134.670 179.120 134.930 179.440 ;
        RECT 134.210 177.080 134.470 177.400 ;
        RECT 134.270 176.120 134.410 177.080 ;
        RECT 134.730 177.060 134.870 179.120 ;
        RECT 135.130 178.780 135.390 179.100 ;
        RECT 135.190 178.420 135.330 178.780 ;
        RECT 135.130 178.100 135.390 178.420 ;
        RECT 135.590 178.100 135.850 178.420 ;
        RECT 134.670 176.740 134.930 177.060 ;
        RECT 135.650 176.720 135.790 178.100 ;
        RECT 136.570 177.595 136.710 183.540 ;
        RECT 136.970 178.440 137.230 178.760 ;
        RECT 136.050 177.080 136.310 177.400 ;
        RECT 136.500 177.225 136.780 177.595 ;
        RECT 135.590 176.400 135.850 176.720 ;
        RECT 136.110 176.120 136.250 177.080 ;
        RECT 137.030 176.380 137.170 178.440 ;
        RECT 134.270 175.980 134.870 176.120 ;
        RECT 133.750 175.380 134.010 175.700 ;
        RECT 134.210 175.380 134.470 175.700 ;
        RECT 133.280 173.825 133.560 174.195 ;
        RECT 132.370 171.640 132.630 171.960 ;
        RECT 133.810 170.940 133.950 175.380 ;
        RECT 133.750 170.620 134.010 170.940 ;
        RECT 132.370 170.280 132.630 170.600 ;
        RECT 133.290 170.280 133.550 170.600 ;
        RECT 132.430 169.240 132.570 170.280 ;
        RECT 132.370 169.150 132.630 169.240 ;
        RECT 132.370 169.010 133.030 169.150 ;
        RECT 132.370 168.920 132.630 169.010 ;
        RECT 131.910 168.240 132.170 168.560 ;
        RECT 132.370 168.240 132.630 168.560 ;
        RECT 132.430 167.395 132.570 168.240 ;
        RECT 132.890 167.960 133.030 169.010 ;
        RECT 133.350 168.560 133.490 170.280 ;
        RECT 133.750 168.920 134.010 169.240 ;
        RECT 133.810 168.560 133.950 168.920 ;
        RECT 133.290 168.240 133.550 168.560 ;
        RECT 133.750 168.240 134.010 168.560 ;
        RECT 132.890 167.820 133.490 167.960 ;
        RECT 132.360 167.025 132.640 167.395 ;
        RECT 132.830 167.220 133.090 167.540 ;
        RECT 132.360 165.665 132.640 166.035 ;
        RECT 132.370 165.520 132.630 165.665 ;
        RECT 132.890 163.800 133.030 167.220 ;
        RECT 132.830 163.480 133.090 163.800 ;
        RECT 132.370 162.800 132.630 163.120 ;
        RECT 132.430 161.080 132.570 162.800 ;
        RECT 133.350 162.100 133.490 167.820 ;
        RECT 133.750 167.560 134.010 167.880 ;
        RECT 133.290 161.780 133.550 162.100 ;
        RECT 132.370 160.760 132.630 161.080 ;
        RECT 129.610 159.740 129.870 160.060 ;
        RECT 131.450 159.740 131.710 160.060 ;
        RECT 129.670 158.360 129.810 159.740 ;
        RECT 129.610 158.040 129.870 158.360 ;
        RECT 129.610 157.360 129.870 157.680 ;
        RECT 130.060 157.590 130.340 157.875 ;
        RECT 131.450 157.700 131.710 158.020 ;
        RECT 130.060 157.505 130.730 157.590 ;
        RECT 130.070 157.450 130.730 157.505 ;
        RECT 130.070 157.360 130.330 157.450 ;
        RECT 129.670 149.860 129.810 157.360 ;
        RECT 130.070 156.340 130.330 156.660 ;
        RECT 129.610 149.540 129.870 149.860 ;
        RECT 130.130 149.180 130.270 156.340 ;
        RECT 130.590 149.180 130.730 157.450 ;
        RECT 130.990 154.640 131.250 154.960 ;
        RECT 131.050 152.920 131.190 154.640 ;
        RECT 130.990 152.600 131.250 152.920 ;
        RECT 130.070 148.860 130.330 149.180 ;
        RECT 130.530 148.860 130.790 149.180 ;
        RECT 130.070 148.180 130.330 148.500 ;
        RECT 129.150 146.480 129.410 146.800 ;
        RECT 124.550 144.580 125.210 144.720 ;
        RECT 124.550 144.440 124.810 144.580 ;
        RECT 125.070 143.740 125.210 144.580 ;
        RECT 125.010 143.420 125.270 143.740 ;
        RECT 128.230 143.080 128.490 143.400 ;
        RECT 122.250 142.740 122.510 143.060 ;
        RECT 128.290 142.040 128.430 143.080 ;
        RECT 128.230 141.720 128.490 142.040 ;
        RECT 129.150 141.040 129.410 141.360 ;
        RECT 122.250 140.700 122.510 141.020 ;
        RECT 120.870 138.890 121.130 138.980 ;
        RECT 120.870 138.750 121.530 138.890 ;
        RECT 120.870 138.660 121.130 138.750 ;
        RECT 120.870 137.980 121.130 138.300 ;
        RECT 119.490 134.580 119.750 134.900 ;
        RECT 118.570 132.880 118.830 133.200 ;
        RECT 119.550 130.920 119.690 134.580 ;
        RECT 119.550 130.780 120.150 130.920 ;
        RECT 117.650 128.120 117.910 128.440 ;
        RECT 120.010 127.420 120.150 130.780 ;
        RECT 120.930 127.420 121.070 137.980 ;
        RECT 121.390 136.260 121.530 138.750 ;
        RECT 122.310 136.600 122.450 140.700 ;
        RECT 129.210 139.320 129.350 141.040 ;
        RECT 127.310 139.000 127.570 139.320 ;
        RECT 129.150 139.000 129.410 139.320 ;
        RECT 122.710 137.640 122.970 137.960 ;
        RECT 122.250 136.280 122.510 136.600 ;
        RECT 121.330 135.940 121.590 136.260 ;
        RECT 122.770 133.880 122.910 137.640 ;
        RECT 127.370 135.920 127.510 139.000 ;
        RECT 130.130 138.640 130.270 148.180 ;
        RECT 130.590 147.140 130.730 148.860 ;
        RECT 130.530 146.820 130.790 147.140 ;
        RECT 131.510 144.720 131.650 157.700 ;
        RECT 133.350 157.680 133.490 161.780 ;
        RECT 133.810 160.400 133.950 167.560 ;
        RECT 134.270 165.500 134.410 175.380 ;
        RECT 134.730 170.940 134.870 175.980 ;
        RECT 135.650 175.980 136.250 176.120 ;
        RECT 136.970 176.060 137.230 176.380 ;
        RECT 135.130 173.680 135.390 174.000 ;
        RECT 134.670 170.620 134.930 170.940 ;
        RECT 134.670 169.940 134.930 170.260 ;
        RECT 134.210 165.180 134.470 165.500 ;
        RECT 134.210 162.800 134.470 163.120 ;
        RECT 133.750 160.080 134.010 160.400 ;
        RECT 133.810 157.680 133.950 160.080 ;
        RECT 133.290 157.360 133.550 157.680 ;
        RECT 133.750 157.360 134.010 157.680 ;
        RECT 133.810 154.960 133.950 157.360 ;
        RECT 133.750 154.640 134.010 154.960 ;
        RECT 133.810 152.580 133.950 154.640 ;
        RECT 133.750 152.260 134.010 152.580 ;
        RECT 131.910 148.180 132.170 148.500 ;
        RECT 131.050 144.580 131.650 144.720 ;
        RECT 130.530 142.740 130.790 143.060 ;
        RECT 130.590 141.360 130.730 142.740 ;
        RECT 130.530 141.040 130.790 141.360 ;
        RECT 130.070 138.320 130.330 138.640 ;
        RECT 127.310 135.600 127.570 135.920 ;
        RECT 123.170 134.580 123.430 134.900 ;
        RECT 122.710 133.560 122.970 133.880 ;
        RECT 123.230 133.200 123.370 134.580 ;
        RECT 128.230 133.220 128.490 133.540 ;
        RECT 123.170 132.880 123.430 133.200 ;
        RECT 126.390 129.820 126.650 130.140 ;
        RECT 121.330 129.140 121.590 129.460 ;
        RECT 118.110 127.100 118.370 127.420 ;
        RECT 119.950 127.100 120.210 127.420 ;
        RECT 120.870 127.100 121.130 127.420 ;
        RECT 115.810 125.400 116.070 125.720 ;
        RECT 118.170 125.380 118.310 127.100 ;
        RECT 119.490 126.760 119.750 127.080 ;
        RECT 118.110 125.060 118.370 125.380 ;
        RECT 114.890 124.720 115.150 125.040 ;
        RECT 114.030 124.300 114.630 124.440 ;
        RECT 116.270 124.380 116.530 124.700 ;
        RECT 113.970 123.700 114.230 124.020 ;
        RECT 113.110 122.260 113.710 122.400 ;
        RECT 110.750 121.660 111.010 121.980 ;
        RECT 108.910 119.850 109.170 119.940 ;
        RECT 108.910 119.710 109.570 119.850 ;
        RECT 108.910 119.620 109.170 119.710 ;
        RECT 108.910 118.940 109.170 119.260 ;
        RECT 108.450 116.560 108.710 116.880 ;
        RECT 107.990 116.220 108.250 116.540 ;
        RECT 108.050 114.500 108.190 116.220 ;
        RECT 107.990 114.180 108.250 114.500 ;
        RECT 108.050 113.140 108.190 114.180 ;
        RECT 108.510 113.480 108.650 116.560 ;
        RECT 108.970 115.860 109.110 118.940 ;
        RECT 108.910 115.540 109.170 115.860 ;
        RECT 108.450 113.160 108.710 113.480 ;
        RECT 107.990 112.820 108.250 113.140 ;
        RECT 107.070 102.620 107.330 102.940 ;
        RECT 106.610 100.920 106.870 101.240 ;
        RECT 105.230 100.580 105.490 100.900 ;
        RECT 107.130 100.220 107.270 102.620 ;
        RECT 104.310 99.900 104.570 100.220 ;
        RECT 107.070 99.900 107.330 100.220 ;
        RECT 104.370 94.780 104.510 99.900 ;
        RECT 104.770 99.560 105.030 99.880 ;
        RECT 107.530 99.560 107.790 99.880 ;
        RECT 104.830 96.820 104.970 99.560 ;
        RECT 107.590 98.520 107.730 99.560 ;
        RECT 107.530 98.200 107.790 98.520 ;
        RECT 104.770 96.500 105.030 96.820 ;
        RECT 97.410 94.460 97.670 94.780 ;
        RECT 102.930 94.460 103.190 94.780 ;
        RECT 104.310 94.460 104.570 94.780 ;
        RECT 98.790 93.780 99.050 94.100 ;
        RECT 102.010 93.780 102.270 94.100 ;
        RECT 98.850 86.550 98.990 93.780 ;
        RECT 102.070 86.550 102.210 93.780 ;
        RECT 104.830 92.740 104.970 96.500 ;
        RECT 108.050 94.780 108.190 112.820 ;
        RECT 108.510 106.000 108.650 113.160 ;
        RECT 109.430 111.100 109.570 119.710 ;
        RECT 109.830 118.260 110.090 118.580 ;
        RECT 109.890 111.780 110.030 118.260 ;
        RECT 110.290 115.880 110.550 116.200 ;
        RECT 110.350 112.120 110.490 115.880 ;
        RECT 110.290 111.800 110.550 112.120 ;
        RECT 109.830 111.460 110.090 111.780 ;
        RECT 109.370 110.780 109.630 111.100 ;
        RECT 109.430 109.060 109.570 110.780 ;
        RECT 109.370 108.740 109.630 109.060 ;
        RECT 108.910 107.720 109.170 108.040 ;
        RECT 108.450 105.680 108.710 106.000 ;
        RECT 108.450 104.660 108.710 104.980 ;
        RECT 108.510 97.160 108.650 104.660 ;
        RECT 108.970 103.960 109.110 107.720 ;
        RECT 109.370 107.380 109.630 107.700 ;
        RECT 108.910 103.640 109.170 103.960 ;
        RECT 109.430 103.620 109.570 107.380 ;
        RECT 110.290 104.660 110.550 104.980 ;
        RECT 110.350 103.620 110.490 104.660 ;
        RECT 109.370 103.300 109.630 103.620 ;
        RECT 110.290 103.300 110.550 103.620 ;
        RECT 110.810 98.180 110.950 121.660 ;
        RECT 111.210 115.540 111.470 115.860 ;
        RECT 111.270 114.160 111.410 115.540 ;
        RECT 111.210 113.840 111.470 114.160 ;
        RECT 110.750 97.860 111.010 98.180 ;
        RECT 108.450 96.840 108.710 97.160 ;
        RECT 111.270 94.780 111.410 113.840 ;
        RECT 112.590 108.740 112.850 109.060 ;
        RECT 111.670 107.380 111.930 107.700 ;
        RECT 111.730 106.340 111.870 107.380 ;
        RECT 111.670 106.020 111.930 106.340 ;
        RECT 112.650 98.180 112.790 108.740 ;
        RECT 113.110 105.320 113.250 122.260 ;
        RECT 113.510 121.660 113.770 121.980 ;
        RECT 113.570 117.560 113.710 121.660 ;
        RECT 114.030 118.920 114.170 123.700 ;
        RECT 113.970 118.600 114.230 118.920 ;
        RECT 113.510 117.240 113.770 117.560 ;
        RECT 114.490 111.100 114.630 124.300 ;
        RECT 115.350 122.680 115.610 123.000 ;
        RECT 114.890 121.320 115.150 121.640 ;
        RECT 114.950 120.280 115.090 121.320 ;
        RECT 115.410 121.300 115.550 122.680 ;
        RECT 116.330 121.980 116.470 124.380 ;
        RECT 116.270 121.660 116.530 121.980 ;
        RECT 115.350 120.980 115.610 121.300 ;
        RECT 114.890 119.960 115.150 120.280 ;
        RECT 119.030 118.260 119.290 118.580 ;
        RECT 114.890 114.180 115.150 114.500 ;
        RECT 114.430 111.010 114.690 111.100 ;
        RECT 114.030 110.870 114.690 111.010 ;
        RECT 114.030 108.380 114.170 110.870 ;
        RECT 114.430 110.780 114.690 110.870 ;
        RECT 114.430 110.100 114.690 110.420 ;
        RECT 113.970 108.060 114.230 108.380 ;
        RECT 114.490 106.680 114.630 110.100 ;
        RECT 114.430 106.360 114.690 106.680 ;
        RECT 114.950 106.340 115.090 114.180 ;
        RECT 116.730 113.500 116.990 113.820 ;
        RECT 116.790 108.720 116.930 113.500 ;
        RECT 118.570 110.440 118.830 110.760 ;
        RECT 117.650 110.100 117.910 110.420 ;
        RECT 116.730 108.400 116.990 108.720 ;
        RECT 114.890 106.020 115.150 106.340 ;
        RECT 116.790 105.660 116.930 108.400 ;
        RECT 117.710 108.040 117.850 110.100 ;
        RECT 118.630 109.400 118.770 110.440 ;
        RECT 118.110 109.080 118.370 109.400 ;
        RECT 118.570 109.080 118.830 109.400 ;
        RECT 117.650 107.720 117.910 108.040 ;
        RECT 117.190 106.020 117.450 106.340 ;
        RECT 114.890 105.340 115.150 105.660 ;
        RECT 116.730 105.340 116.990 105.660 ;
        RECT 113.050 105.000 113.310 105.320 ;
        RECT 114.950 99.540 115.090 105.340 ;
        RECT 115.350 104.660 115.610 104.980 ;
        RECT 116.730 104.660 116.990 104.980 ;
        RECT 113.050 99.220 113.310 99.540 ;
        RECT 114.890 99.220 115.150 99.540 ;
        RECT 112.590 97.860 112.850 98.180 ;
        RECT 113.110 94.780 113.250 99.220 ;
        RECT 113.510 97.180 113.770 97.500 ;
        RECT 113.570 95.460 113.710 97.180 ;
        RECT 115.410 95.800 115.550 104.660 ;
        RECT 116.790 103.280 116.930 104.660 ;
        RECT 117.250 103.620 117.390 106.020 ;
        RECT 118.170 106.000 118.310 109.080 ;
        RECT 118.110 105.680 118.370 106.000 ;
        RECT 117.650 103.640 117.910 103.960 ;
        RECT 117.190 103.300 117.450 103.620 ;
        RECT 116.730 102.960 116.990 103.280 ;
        RECT 116.790 102.600 116.930 102.960 ;
        RECT 116.730 102.280 116.990 102.600 ;
        RECT 116.270 101.940 116.530 102.260 ;
        RECT 115.810 99.560 116.070 99.880 ;
        RECT 115.870 98.520 116.010 99.560 ;
        RECT 115.810 98.200 116.070 98.520 ;
        RECT 115.350 95.480 115.610 95.800 ;
        RECT 116.330 95.460 116.470 101.940 ;
        RECT 117.710 98.520 117.850 103.640 ;
        RECT 118.110 99.220 118.370 99.540 ;
        RECT 118.170 98.520 118.310 99.220 ;
        RECT 117.650 98.200 117.910 98.520 ;
        RECT 118.110 98.200 118.370 98.520 ;
        RECT 118.170 96.420 118.310 98.200 ;
        RECT 119.090 97.500 119.230 118.260 ;
        RECT 119.550 106.680 119.690 126.760 ;
        RECT 120.410 125.060 120.670 125.380 ;
        RECT 119.950 122.340 120.210 122.660 ;
        RECT 119.490 106.360 119.750 106.680 ;
        RECT 119.030 97.180 119.290 97.500 ;
        RECT 120.010 96.420 120.150 122.340 ;
        RECT 120.470 121.980 120.610 125.060 ;
        RECT 120.410 121.660 120.670 121.980 ;
        RECT 120.930 119.600 121.070 127.100 ;
        RECT 121.390 127.080 121.530 129.140 ;
        RECT 125.010 127.100 125.270 127.420 ;
        RECT 121.330 126.760 121.590 127.080 ;
        RECT 125.070 125.380 125.210 127.100 ;
        RECT 125.010 125.060 125.270 125.380 ;
        RECT 124.550 121.320 124.810 121.640 ;
        RECT 123.630 119.620 123.890 119.940 ;
        RECT 120.870 119.280 121.130 119.600 ;
        RECT 123.690 117.560 123.830 119.620 ;
        RECT 123.630 117.240 123.890 117.560 ;
        RECT 124.610 116.880 124.750 121.320 ;
        RECT 125.010 116.900 125.270 117.220 ;
        RECT 122.250 116.560 122.510 116.880 ;
        RECT 124.550 116.560 124.810 116.880 ;
        RECT 122.310 113.820 122.450 116.560 ;
        RECT 124.090 115.540 124.350 115.860 ;
        RECT 124.150 114.500 124.290 115.540 ;
        RECT 125.070 114.840 125.210 116.900 ;
        RECT 126.450 116.880 126.590 129.820 ;
        RECT 126.850 129.480 127.110 129.800 ;
        RECT 126.910 125.720 127.050 129.480 ;
        RECT 128.290 125.720 128.430 133.220 ;
        RECT 128.690 132.540 128.950 132.860 ;
        RECT 128.750 128.440 128.890 132.540 ;
        RECT 129.150 130.840 129.410 131.160 ;
        RECT 129.210 130.675 129.350 130.840 ;
        RECT 129.140 130.305 129.420 130.675 ;
        RECT 130.130 130.480 130.270 138.320 ;
        RECT 131.050 133.540 131.190 144.580 ;
        RECT 131.450 135.600 131.710 135.920 ;
        RECT 130.990 133.220 131.250 133.540 ;
        RECT 130.530 132.200 130.790 132.520 ;
        RECT 130.070 130.160 130.330 130.480 ;
        RECT 130.590 130.140 130.730 132.200 ;
        RECT 130.530 129.820 130.790 130.140 ;
        RECT 128.690 128.120 128.950 128.440 ;
        RECT 130.590 127.760 130.730 129.820 ;
        RECT 130.530 127.440 130.790 127.760 ;
        RECT 129.150 126.420 129.410 126.740 ;
        RECT 126.850 125.400 127.110 125.720 ;
        RECT 128.230 125.400 128.490 125.720 ;
        RECT 126.390 116.560 126.650 116.880 ;
        RECT 125.010 114.520 125.270 114.840 ;
        RECT 124.090 114.180 124.350 114.500 ;
        RECT 122.250 113.500 122.510 113.820 ;
        RECT 122.310 111.100 122.450 113.500 ;
        RECT 124.550 111.800 124.810 112.120 ;
        RECT 122.250 110.780 122.510 111.100 ;
        RECT 120.870 102.960 121.130 103.280 ;
        RECT 118.170 96.280 118.770 96.420 ;
        RECT 113.510 95.140 113.770 95.460 ;
        RECT 116.270 95.140 116.530 95.460 ;
        RECT 118.110 95.140 118.370 95.460 ;
        RECT 107.990 94.460 108.250 94.780 ;
        RECT 111.210 94.460 111.470 94.780 ;
        RECT 113.050 94.460 113.310 94.780 ;
        RECT 114.890 94.120 115.150 94.440 ;
        RECT 105.230 93.780 105.490 94.100 ;
        RECT 108.450 93.780 108.710 94.100 ;
        RECT 111.670 93.780 111.930 94.100 ;
        RECT 104.770 92.420 105.030 92.740 ;
        RECT 105.290 86.550 105.430 93.780 ;
        RECT 108.510 86.550 108.650 93.780 ;
        RECT 111.730 86.550 111.870 93.780 ;
        RECT 114.950 86.550 115.090 94.120 ;
        RECT 116.270 93.780 116.530 94.100 ;
        RECT 116.330 93.080 116.470 93.780 ;
        RECT 116.270 92.760 116.530 93.080 ;
        RECT 118.170 86.550 118.310 95.140 ;
        RECT 118.630 95.120 118.770 96.280 ;
        RECT 119.550 96.280 120.150 96.420 ;
        RECT 118.570 94.800 118.830 95.120 ;
        RECT 118.630 94.440 118.770 94.800 ;
        RECT 119.550 94.780 119.690 96.280 ;
        RECT 119.950 95.480 120.210 95.800 ;
        RECT 120.010 94.780 120.150 95.480 ;
        RECT 120.930 94.780 121.070 102.960 ;
        RECT 124.610 102.940 124.750 111.800 ;
        RECT 126.450 111.440 126.590 116.560 ;
        RECT 126.390 111.120 126.650 111.440 ;
        RECT 126.450 106.000 126.590 111.120 ;
        RECT 126.390 105.680 126.650 106.000 ;
        RECT 128.290 104.040 128.430 125.400 ;
        RECT 129.210 125.040 129.350 126.420 ;
        RECT 129.150 124.720 129.410 125.040 ;
        RECT 130.990 123.700 131.250 124.020 ;
        RECT 129.150 121.660 129.410 121.980 ;
        RECT 130.530 121.660 130.790 121.980 ;
        RECT 128.690 118.260 128.950 118.580 ;
        RECT 128.750 117.560 128.890 118.260 ;
        RECT 128.690 117.240 128.950 117.560 ;
        RECT 129.210 114.500 129.350 121.660 ;
        RECT 129.610 120.980 129.870 121.300 ;
        RECT 129.150 114.180 129.410 114.500 ;
        RECT 129.670 113.560 129.810 120.980 ;
        RECT 130.590 120.280 130.730 121.660 ;
        RECT 131.050 121.640 131.190 123.700 ;
        RECT 131.510 123.000 131.650 135.600 ;
        RECT 131.970 131.160 132.110 148.180 ;
        RECT 132.830 146.820 133.090 147.140 ;
        RECT 132.370 145.460 132.630 145.780 ;
        RECT 132.430 141.020 132.570 145.460 ;
        RECT 132.890 144.720 133.030 146.820 ;
        RECT 133.810 146.800 133.950 152.260 ;
        RECT 134.270 150.200 134.410 162.800 ;
        RECT 134.730 157.760 134.870 169.940 ;
        RECT 135.190 165.500 135.330 173.680 ;
        RECT 135.130 165.180 135.390 165.500 ;
        RECT 135.190 164.820 135.330 165.180 ;
        RECT 135.130 164.500 135.390 164.820 ;
        RECT 135.650 163.315 135.790 175.980 ;
        RECT 137.490 174.340 137.630 184.560 ;
        RECT 137.950 182.500 138.090 184.560 ;
        RECT 138.870 182.840 139.010 184.560 ;
        RECT 138.810 182.520 139.070 182.840 ;
        RECT 137.890 182.180 138.150 182.500 ;
        RECT 140.710 181.820 140.850 186.260 ;
        RECT 137.890 181.500 138.150 181.820 ;
        RECT 140.650 181.500 140.910 181.820 ;
        RECT 142.090 181.675 142.230 186.940 ;
        RECT 143.930 185.220 144.070 186.940 ;
        RECT 143.870 184.900 144.130 185.220 ;
        RECT 137.950 180.995 138.090 181.500 ;
        RECT 138.350 181.160 138.610 181.480 ;
        RECT 137.880 180.625 138.160 180.995 ;
        RECT 138.410 179.440 138.550 181.160 ;
        RECT 140.710 179.440 140.850 181.500 ;
        RECT 142.020 181.305 142.300 181.675 ;
        RECT 143.930 179.780 144.070 184.900 ;
        RECT 143.870 179.460 144.130 179.780 ;
        RECT 138.350 179.120 138.610 179.440 ;
        RECT 140.650 179.120 140.910 179.440 ;
        RECT 145.250 176.060 145.510 176.380 ;
        RECT 145.310 174.875 145.450 176.060 ;
        RECT 145.240 174.505 145.520 174.875 ;
        RECT 137.430 174.020 137.690 174.340 ;
        RECT 137.890 173.680 138.150 174.000 ;
        RECT 143.870 173.680 144.130 174.000 ;
        RECT 136.510 173.000 136.770 173.320 ;
        RECT 136.570 171.280 136.710 173.000 ;
        RECT 137.950 171.960 138.090 173.680 ;
        RECT 143.410 172.660 143.670 172.980 ;
        RECT 137.890 171.640 138.150 171.960 ;
        RECT 136.510 170.960 136.770 171.280 ;
        RECT 143.470 170.940 143.610 172.660 ;
        RECT 143.410 170.620 143.670 170.940 ;
        RECT 138.810 170.280 139.070 170.600 ;
        RECT 136.050 169.940 136.310 170.260 ;
        RECT 135.580 162.945 135.860 163.315 ;
        RECT 135.130 161.780 135.390 162.100 ;
        RECT 135.190 160.060 135.330 161.780 ;
        RECT 135.130 159.740 135.390 160.060 ;
        RECT 134.730 157.620 135.330 157.760 ;
        RECT 134.210 149.880 134.470 150.200 ;
        RECT 134.670 148.180 134.930 148.500 ;
        RECT 134.730 147.140 134.870 148.180 ;
        RECT 134.670 146.820 134.930 147.140 ;
        RECT 133.750 146.480 134.010 146.800 ;
        RECT 132.890 144.580 133.490 144.720 ;
        RECT 132.370 140.700 132.630 141.020 ;
        RECT 132.370 140.020 132.630 140.340 ;
        RECT 132.430 138.980 132.570 140.020 ;
        RECT 132.370 138.660 132.630 138.980 ;
        RECT 133.350 135.830 133.490 144.580 ;
        RECT 134.210 143.080 134.470 143.400 ;
        RECT 134.270 142.040 134.410 143.080 ;
        RECT 134.210 141.720 134.470 142.040 ;
        RECT 135.190 140.680 135.330 157.620 ;
        RECT 136.110 149.520 136.250 169.940 ;
        RECT 136.970 168.240 137.230 168.560 ;
        RECT 137.030 166.520 137.170 168.240 ;
        RECT 136.970 166.200 137.230 166.520 ;
        RECT 137.890 164.500 138.150 164.820 ;
        RECT 136.510 162.800 136.770 163.120 ;
        RECT 136.570 158.360 136.710 162.800 ;
        RECT 137.950 162.100 138.090 164.500 ;
        RECT 137.890 161.780 138.150 162.100 ;
        RECT 138.870 161.840 139.010 170.280 ;
        RECT 139.730 169.940 139.990 170.260 ;
        RECT 139.790 169.240 139.930 169.940 ;
        RECT 139.730 168.920 139.990 169.240 ;
        RECT 142.490 167.220 142.750 167.540 ;
        RECT 142.550 165.840 142.690 167.220 ;
        RECT 142.490 165.520 142.750 165.840 ;
        RECT 140.650 163.140 140.910 163.460 ;
        RECT 138.870 161.700 139.470 161.840 ;
        RECT 138.810 160.760 139.070 161.080 ;
        RECT 136.510 158.040 136.770 158.360 ;
        RECT 137.430 156.340 137.690 156.660 ;
        RECT 137.490 154.280 137.630 156.340 ;
        RECT 137.430 153.960 137.690 154.280 ;
        RECT 137.490 152.240 137.630 153.960 ;
        RECT 138.870 152.920 139.010 160.760 ;
        RECT 138.810 152.600 139.070 152.920 ;
        RECT 137.430 151.920 137.690 152.240 ;
        RECT 136.050 149.200 136.310 149.520 ;
        RECT 136.050 143.080 136.310 143.400 ;
        RECT 136.110 141.700 136.250 143.080 ;
        RECT 139.330 141.700 139.470 161.700 ;
        RECT 140.710 161.080 140.850 163.140 ;
        RECT 143.470 163.120 143.610 170.620 ;
        RECT 143.930 163.800 144.070 173.680 ;
        RECT 144.790 172.660 145.050 172.980 ;
        RECT 144.850 171.475 144.990 172.660 ;
        RECT 144.780 171.105 145.060 171.475 ;
        RECT 144.330 168.580 144.590 168.900 ;
        RECT 143.870 163.480 144.130 163.800 ;
        RECT 144.390 163.200 144.530 168.580 ;
        RECT 144.780 167.705 145.060 168.075 ;
        RECT 144.790 167.560 145.050 167.705 ;
        RECT 144.780 164.305 145.060 164.675 ;
        RECT 144.850 163.800 144.990 164.305 ;
        RECT 144.790 163.480 145.050 163.800 ;
        RECT 143.410 162.800 143.670 163.120 ;
        RECT 143.930 163.060 144.530 163.200 ;
        RECT 142.950 162.120 143.210 162.440 ;
        RECT 143.010 161.275 143.150 162.120 ;
        RECT 140.650 160.760 140.910 161.080 ;
        RECT 142.940 160.905 143.220 161.275 ;
        RECT 143.400 160.225 143.680 160.595 ;
        RECT 143.930 160.400 144.070 163.060 ;
        RECT 144.780 162.945 145.060 163.315 ;
        RECT 145.250 163.140 145.510 163.460 ;
        RECT 143.410 160.080 143.670 160.225 ;
        RECT 143.870 160.080 144.130 160.400 ;
        RECT 141.110 159.060 141.370 159.380 ;
        RECT 142.950 159.060 143.210 159.380 ;
        RECT 141.170 158.020 141.310 159.060 ;
        RECT 141.110 157.700 141.370 158.020 ;
        RECT 141.570 156.340 141.830 156.660 ;
        RECT 141.630 154.620 141.770 156.340 ;
        RECT 143.010 155.640 143.150 159.060 ;
        RECT 144.850 157.340 144.990 162.945 ;
        RECT 145.310 157.875 145.450 163.140 ;
        RECT 145.240 157.505 145.520 157.875 ;
        RECT 143.870 157.020 144.130 157.340 ;
        RECT 144.790 157.020 145.050 157.340 ;
        RECT 142.950 155.320 143.210 155.640 ;
        RECT 143.410 154.980 143.670 155.300 ;
        RECT 141.570 154.300 141.830 154.620 ;
        RECT 142.030 153.620 142.290 153.940 ;
        RECT 142.090 152.240 142.230 153.620 ;
        RECT 142.950 152.600 143.210 152.920 ;
        RECT 140.190 152.150 140.450 152.240 ;
        RECT 139.790 152.010 140.450 152.150 ;
        RECT 139.790 147.480 139.930 152.010 ;
        RECT 140.190 151.920 140.450 152.010 ;
        RECT 142.030 151.920 142.290 152.240 ;
        RECT 143.010 151.075 143.150 152.600 ;
        RECT 142.940 150.705 143.220 151.075 ;
        RECT 143.470 149.180 143.610 154.980 ;
        RECT 143.930 152.920 144.070 157.020 ;
        RECT 144.780 154.105 145.060 154.475 ;
        RECT 143.870 152.600 144.130 152.920 ;
        RECT 143.870 151.580 144.130 151.900 ;
        RECT 143.930 149.180 144.070 151.580 ;
        RECT 144.850 150.200 144.990 154.105 ;
        RECT 144.790 149.880 145.050 150.200 ;
        RECT 140.190 148.860 140.450 149.180 ;
        RECT 143.410 148.860 143.670 149.180 ;
        RECT 143.870 148.860 144.130 149.180 ;
        RECT 140.250 147.480 140.390 148.860 ;
        RECT 139.730 147.160 139.990 147.480 ;
        RECT 140.190 147.160 140.450 147.480 ;
        RECT 144.780 147.305 145.060 147.675 ;
        RECT 144.790 147.160 145.050 147.305 ;
        RECT 142.950 145.460 143.210 145.780 ;
        RECT 143.010 144.275 143.150 145.460 ;
        RECT 142.030 143.760 142.290 144.080 ;
        RECT 142.940 143.905 143.220 144.275 ;
        RECT 141.110 142.740 141.370 143.060 ;
        RECT 141.170 142.040 141.310 142.740 ;
        RECT 141.110 141.720 141.370 142.040 ;
        RECT 136.050 141.380 136.310 141.700 ;
        RECT 139.270 141.380 139.530 141.700 ;
        RECT 135.590 141.040 135.850 141.360 ;
        RECT 135.130 140.360 135.390 140.680 ;
        RECT 135.650 138.300 135.790 141.040 ;
        RECT 134.670 137.980 134.930 138.300 ;
        RECT 135.590 137.980 135.850 138.300 ;
        RECT 134.730 136.600 134.870 137.980 ;
        RECT 136.110 137.620 136.250 141.380 ;
        RECT 136.510 138.660 136.770 138.980 ;
        RECT 136.050 137.300 136.310 137.620 ;
        RECT 136.570 137.360 136.710 138.660 ;
        RECT 136.970 138.210 137.230 138.300 ;
        RECT 136.970 138.070 139.010 138.210 ;
        RECT 136.970 137.980 137.230 138.070 ;
        RECT 134.670 136.280 134.930 136.600 ;
        RECT 133.750 135.830 134.010 135.920 ;
        RECT 133.350 135.690 134.010 135.830 ;
        RECT 131.910 130.840 132.170 131.160 ;
        RECT 131.910 129.140 132.170 129.460 ;
        RECT 132.370 129.140 132.630 129.460 ;
        RECT 131.970 125.720 132.110 129.140 ;
        RECT 132.430 128.100 132.570 129.140 ;
        RECT 132.370 127.780 132.630 128.100 ;
        RECT 131.910 125.400 132.170 125.720 ;
        RECT 131.450 122.680 131.710 123.000 ;
        RECT 133.350 122.320 133.490 135.690 ;
        RECT 133.750 135.600 134.010 135.690 ;
        RECT 134.210 130.160 134.470 130.480 ;
        RECT 133.750 129.480 134.010 129.800 ;
        RECT 133.810 123.000 133.950 129.480 ;
        RECT 133.750 122.680 134.010 123.000 ;
        RECT 133.290 122.000 133.550 122.320 ;
        RECT 130.990 121.320 131.250 121.640 ;
        RECT 130.530 119.960 130.790 120.280 ;
        RECT 133.350 119.600 133.490 122.000 ;
        RECT 134.270 119.940 134.410 130.160 ;
        RECT 134.730 127.420 134.870 136.280 ;
        RECT 136.110 135.580 136.250 137.300 ;
        RECT 136.570 137.220 137.170 137.360 ;
        RECT 136.510 135.600 136.770 135.920 ;
        RECT 136.050 135.260 136.310 135.580 ;
        RECT 135.590 134.580 135.850 134.900 ;
        RECT 135.650 133.540 135.790 134.580 ;
        RECT 135.590 133.220 135.850 133.540 ;
        RECT 135.130 129.480 135.390 129.800 ;
        RECT 135.190 127.420 135.330 129.480 ;
        RECT 136.110 128.100 136.250 135.260 ;
        RECT 136.570 133.880 136.710 135.600 ;
        RECT 136.510 133.560 136.770 133.880 ;
        RECT 136.510 131.860 136.770 132.180 ;
        RECT 136.050 127.780 136.310 128.100 ;
        RECT 134.670 127.100 134.930 127.420 ;
        RECT 135.130 127.100 135.390 127.420 ;
        RECT 135.190 126.740 135.330 127.100 ;
        RECT 135.130 126.420 135.390 126.740 ;
        RECT 136.050 122.000 136.310 122.320 ;
        RECT 136.110 120.280 136.250 122.000 ;
        RECT 136.050 119.960 136.310 120.280 ;
        RECT 134.210 119.620 134.470 119.940 ;
        RECT 133.290 119.280 133.550 119.600 ;
        RECT 132.830 118.940 133.090 119.260 ;
        RECT 131.450 116.220 131.710 116.540 ;
        RECT 129.210 113.420 129.810 113.560 ;
        RECT 128.690 104.660 128.950 104.980 ;
        RECT 126.910 103.960 128.430 104.040 ;
        RECT 126.850 103.900 128.430 103.960 ;
        RECT 126.850 103.640 127.110 103.900 ;
        RECT 128.750 103.620 128.890 104.660 ;
        RECT 128.690 103.300 128.950 103.620 ;
        RECT 123.630 102.620 123.890 102.940 ;
        RECT 124.550 102.620 124.810 102.940 ;
        RECT 123.690 101.240 123.830 102.620 ;
        RECT 123.630 100.920 123.890 101.240 ;
        RECT 122.710 99.900 122.970 100.220 ;
        RECT 122.770 98.180 122.910 99.900 ;
        RECT 124.090 99.560 124.350 99.880 ;
        RECT 122.710 97.860 122.970 98.180 ;
        RECT 119.490 94.460 119.750 94.780 ;
        RECT 119.950 94.460 120.210 94.780 ;
        RECT 120.870 94.460 121.130 94.780 ;
        RECT 118.570 94.120 118.830 94.440 ;
        RECT 119.030 94.120 119.290 94.440 ;
        RECT 121.330 94.120 121.590 94.440 ;
        RECT 119.090 92.740 119.230 94.120 ;
        RECT 119.030 92.420 119.290 92.740 ;
        RECT 121.390 86.550 121.530 94.120 ;
        RECT 124.150 93.080 124.290 99.560 ;
        RECT 124.610 95.120 124.750 102.620 ;
        RECT 125.930 100.920 126.190 101.240 ;
        RECT 125.990 95.800 126.130 100.920 ;
        RECT 129.210 97.160 129.350 113.420 ;
        RECT 130.990 107.720 131.250 108.040 ;
        RECT 129.610 107.380 129.870 107.700 ;
        RECT 129.670 105.320 129.810 107.380 ;
        RECT 131.050 106.340 131.190 107.720 ;
        RECT 130.530 106.020 130.790 106.340 ;
        RECT 130.990 106.020 131.250 106.340 ;
        RECT 129.610 105.000 129.870 105.320 ;
        RECT 129.150 96.840 129.410 97.160 ;
        RECT 129.670 96.820 129.810 105.000 ;
        RECT 130.070 99.220 130.330 99.540 ;
        RECT 130.130 97.840 130.270 99.220 ;
        RECT 130.590 98.520 130.730 106.020 ;
        RECT 131.050 103.620 131.190 106.020 ;
        RECT 131.510 105.660 131.650 116.220 ;
        RECT 132.890 113.820 133.030 118.940 ;
        RECT 134.270 116.540 134.410 119.620 ;
        RECT 136.570 119.510 136.710 131.860 ;
        RECT 137.030 127.760 137.170 137.220 ;
        RECT 137.430 130.840 137.690 131.160 ;
        RECT 136.970 127.440 137.230 127.760 ;
        RECT 137.030 124.555 137.170 127.440 ;
        RECT 136.960 124.185 137.240 124.555 ;
        RECT 136.570 119.370 137.170 119.510 ;
        RECT 136.050 118.940 136.310 119.260 ;
        RECT 136.110 117.220 136.250 118.940 ;
        RECT 136.510 118.600 136.770 118.920 ;
        RECT 136.570 117.560 136.710 118.600 ;
        RECT 136.510 117.240 136.770 117.560 ;
        RECT 136.050 116.900 136.310 117.220 ;
        RECT 134.210 116.220 134.470 116.540 ;
        RECT 132.830 113.500 133.090 113.820 ;
        RECT 132.890 112.120 133.030 113.500 ;
        RECT 133.290 112.820 133.550 113.140 ;
        RECT 132.830 111.800 133.090 112.120 ;
        RECT 133.350 111.780 133.490 112.820 ;
        RECT 133.290 111.460 133.550 111.780 ;
        RECT 136.110 111.440 136.250 116.900 ;
        RECT 136.510 112.820 136.770 113.140 ;
        RECT 136.050 111.120 136.310 111.440 ;
        RECT 136.110 108.720 136.250 111.120 ;
        RECT 132.370 108.400 132.630 108.720 ;
        RECT 135.590 108.400 135.850 108.720 ;
        RECT 136.050 108.400 136.310 108.720 ;
        RECT 131.450 105.340 131.710 105.660 ;
        RECT 130.990 103.300 131.250 103.620 ;
        RECT 130.990 100.580 131.250 100.900 ;
        RECT 130.530 98.200 130.790 98.520 ;
        RECT 130.070 97.520 130.330 97.840 ;
        RECT 130.070 96.840 130.330 97.160 ;
        RECT 129.610 96.500 129.870 96.820 ;
        RECT 130.130 96.420 130.270 96.840 ;
        RECT 130.130 96.280 130.730 96.420 ;
        RECT 125.930 95.480 126.190 95.800 ;
        RECT 125.010 95.140 125.270 95.460 ;
        RECT 124.550 94.800 124.810 95.120 ;
        RECT 124.090 92.760 124.350 93.080 ;
        RECT 125.070 88.400 125.210 95.140 ;
        RECT 125.990 94.780 126.130 95.480 ;
        RECT 130.590 94.780 130.730 96.280 ;
        RECT 131.050 95.800 131.190 100.580 ;
        RECT 131.450 96.840 131.710 97.160 ;
        RECT 131.510 96.675 131.650 96.840 ;
        RECT 131.440 96.305 131.720 96.675 ;
        RECT 130.990 95.480 131.250 95.800 ;
        RECT 130.990 95.030 131.250 95.120 ;
        RECT 131.510 95.030 131.650 96.305 ;
        RECT 130.990 94.890 131.650 95.030 ;
        RECT 130.990 94.800 131.250 94.890 ;
        RECT 132.430 94.780 132.570 108.400 ;
        RECT 133.750 108.060 134.010 108.380 ;
        RECT 133.810 106.000 133.950 108.060 ;
        RECT 133.750 105.680 134.010 106.000 ;
        RECT 133.810 102.940 133.950 105.680 ;
        RECT 135.650 105.660 135.790 108.400 ;
        RECT 135.590 105.340 135.850 105.660 ;
        RECT 133.750 102.620 134.010 102.940 ;
        RECT 133.290 101.940 133.550 102.260 ;
        RECT 132.830 99.220 133.090 99.540 ;
        RECT 132.890 98.520 133.030 99.220 ;
        RECT 133.350 98.520 133.490 101.940 ;
        RECT 133.810 100.560 133.950 102.620 ;
        RECT 136.110 102.600 136.250 108.400 ;
        RECT 136.570 108.040 136.710 112.820 ;
        RECT 136.510 107.720 136.770 108.040 ;
        RECT 137.030 106.760 137.170 119.370 ;
        RECT 137.490 116.540 137.630 130.840 ;
        RECT 138.350 129.820 138.610 130.140 ;
        RECT 138.410 124.360 138.550 129.820 ;
        RECT 138.350 124.040 138.610 124.360 ;
        RECT 137.430 116.220 137.690 116.540 ;
        RECT 137.490 114.840 137.630 116.220 ;
        RECT 137.430 114.520 137.690 114.840 ;
        RECT 137.490 114.160 137.630 114.520 ;
        RECT 137.430 113.840 137.690 114.160 ;
        RECT 137.890 113.500 138.150 113.820 ;
        RECT 137.950 110.420 138.090 113.500 ;
        RECT 137.890 110.100 138.150 110.420 ;
        RECT 137.030 106.620 137.630 106.760 ;
        RECT 136.510 106.020 136.770 106.340 ;
        RECT 136.570 103.960 136.710 106.020 ;
        RECT 136.970 105.680 137.230 106.000 ;
        RECT 136.510 103.640 136.770 103.960 ;
        RECT 136.050 102.280 136.310 102.600 ;
        RECT 136.110 101.240 136.250 102.280 ;
        RECT 136.050 100.920 136.310 101.240 ;
        RECT 136.110 100.640 136.250 100.920 ;
        RECT 133.750 100.240 134.010 100.560 ;
        RECT 136.110 100.500 136.710 100.640 ;
        RECT 132.830 98.200 133.090 98.520 ;
        RECT 133.290 98.200 133.550 98.520 ;
        RECT 125.930 94.460 126.190 94.780 ;
        RECT 130.530 94.460 130.790 94.780 ;
        RECT 132.370 94.460 132.630 94.780 ;
        RECT 130.990 94.120 131.250 94.440 ;
        RECT 127.770 89.020 128.030 89.340 ;
        RECT 124.610 88.260 125.210 88.400 ;
        RECT 124.610 86.550 124.750 88.260 ;
        RECT 127.830 86.550 127.970 89.020 ;
        RECT 131.050 86.550 131.190 94.120 ;
        RECT 132.890 94.100 133.030 98.200 ;
        RECT 133.810 97.160 133.950 100.240 ;
        RECT 135.130 98.200 135.390 98.520 ;
        RECT 133.750 96.840 134.010 97.160 ;
        RECT 135.190 94.780 135.330 98.200 ;
        RECT 136.570 97.840 136.710 100.500 ;
        RECT 137.030 100.220 137.170 105.680 ;
        RECT 137.490 103.960 137.630 106.620 ;
        RECT 137.950 105.660 138.090 110.100 ;
        RECT 137.890 105.340 138.150 105.660 ;
        RECT 138.350 105.000 138.610 105.320 ;
        RECT 138.410 103.960 138.550 105.000 ;
        RECT 137.430 103.640 137.690 103.960 ;
        RECT 138.350 103.640 138.610 103.960 ;
        RECT 137.490 102.680 137.630 103.640 ;
        RECT 137.490 102.540 138.090 102.680 ;
        RECT 137.430 101.940 137.690 102.260 ;
        RECT 136.970 99.900 137.230 100.220 ;
        RECT 136.050 97.520 136.310 97.840 ;
        RECT 136.510 97.520 136.770 97.840 ;
        RECT 135.130 94.635 135.390 94.780 ;
        RECT 135.120 94.265 135.400 94.635 ;
        RECT 135.590 94.460 135.850 94.780 ;
        RECT 132.830 93.780 133.090 94.100 ;
        RECT 135.650 92.740 135.790 94.460 ;
        RECT 135.590 92.420 135.850 92.740 ;
        RECT 136.110 89.340 136.250 97.520 ;
        RECT 136.510 97.070 136.770 97.160 ;
        RECT 136.510 96.930 137.170 97.070 ;
        RECT 136.510 96.840 136.770 96.930 ;
        RECT 136.500 96.305 136.780 96.675 ;
        RECT 136.570 94.780 136.710 96.305 ;
        RECT 136.510 94.460 136.770 94.780 ;
        RECT 137.030 94.690 137.170 96.930 ;
        RECT 137.490 95.460 137.630 101.940 ;
        RECT 137.950 99.540 138.090 102.540 ;
        RECT 137.890 99.220 138.150 99.540 ;
        RECT 138.870 95.800 139.010 138.070 ;
        RECT 139.330 132.180 139.470 141.380 ;
        RECT 142.090 141.360 142.230 143.760 ;
        RECT 142.030 141.040 142.290 141.360 ;
        RECT 140.650 140.700 140.910 141.020 ;
        RECT 140.710 134.900 140.850 140.700 ;
        RECT 144.330 140.360 144.590 140.680 ;
        RECT 144.780 140.505 145.060 140.875 ;
        RECT 144.790 140.360 145.050 140.505 ;
        RECT 144.390 139.320 144.530 140.360 ;
        RECT 144.330 139.000 144.590 139.320 ;
        RECT 144.390 135.920 144.530 139.000 ;
        RECT 144.780 137.105 145.060 137.475 ;
        RECT 144.850 136.600 144.990 137.105 ;
        RECT 144.790 136.280 145.050 136.600 ;
        RECT 144.330 135.600 144.590 135.920 ;
        RECT 143.870 134.920 144.130 135.240 ;
        RECT 140.650 134.580 140.910 134.900 ;
        RECT 139.270 131.860 139.530 132.180 ;
        RECT 140.710 130.140 140.850 134.580 ;
        RECT 143.930 132.860 144.070 134.920 ;
        RECT 144.780 133.705 145.060 134.075 ;
        RECT 144.790 133.560 145.050 133.705 ;
        RECT 142.030 132.540 142.290 132.860 ;
        RECT 143.870 132.540 144.130 132.860 ;
        RECT 142.090 130.820 142.230 132.540 ;
        RECT 142.950 131.860 143.210 132.180 ;
        RECT 142.030 130.500 142.290 130.820 ;
        RECT 143.010 130.675 143.150 131.860 ;
        RECT 142.940 130.305 143.220 130.675 ;
        RECT 140.650 129.820 140.910 130.140 ;
        RECT 140.650 127.100 140.910 127.420 ;
        RECT 139.270 124.040 139.530 124.360 ;
        RECT 139.330 121.640 139.470 124.040 ;
        RECT 139.730 122.000 139.990 122.320 ;
        RECT 139.270 121.320 139.530 121.640 ;
        RECT 139.270 118.320 139.530 118.580 ;
        RECT 139.790 118.320 139.930 122.000 ;
        RECT 139.270 118.260 139.930 118.320 ;
        RECT 139.330 118.180 139.930 118.260 ;
        RECT 139.790 116.880 139.930 118.180 ;
        RECT 139.730 116.560 139.990 116.880 ;
        RECT 139.790 114.840 139.930 116.560 ;
        RECT 140.710 115.860 140.850 127.100 ;
        RECT 144.780 126.905 145.060 127.275 ;
        RECT 143.870 126.420 144.130 126.740 ;
        RECT 142.950 124.040 143.210 124.360 ;
        RECT 143.010 123.875 143.150 124.040 ;
        RECT 142.940 123.505 143.220 123.875 ;
        RECT 141.570 122.340 141.830 122.660 ;
        RECT 141.630 116.540 141.770 122.340 ;
        RECT 143.930 121.980 144.070 126.420 ;
        RECT 144.850 125.720 144.990 126.905 ;
        RECT 144.790 125.400 145.050 125.720 ;
        RECT 147.430 124.640 147.570 221.710 ;
        RECT 150.390 174.360 150.990 175.020 ;
        RECT 151.220 170.940 151.930 171.630 ;
        RECT 148.730 167.540 149.410 168.190 ;
        RECT 148.950 165.245 149.160 167.540 ;
        RECT 148.535 165.035 149.160 165.245 ;
        RECT 147.800 143.850 148.310 144.300 ;
        RECT 147.430 124.500 147.820 124.640 ;
        RECT 143.870 121.660 144.130 121.980 ;
        RECT 142.490 120.980 142.750 121.300 ;
        RECT 142.950 120.980 143.210 121.300 ;
        RECT 144.790 120.980 145.050 121.300 ;
        RECT 142.550 116.540 142.690 120.980 ;
        RECT 143.010 117.075 143.150 120.980 ;
        RECT 144.850 120.475 144.990 120.980 ;
        RECT 144.780 120.105 145.060 120.475 ;
        RECT 144.330 118.260 144.590 118.580 ;
        RECT 142.940 116.705 143.220 117.075 ;
        RECT 144.390 116.880 144.530 118.260 ;
        RECT 144.330 116.560 144.590 116.880 ;
        RECT 141.570 116.220 141.830 116.540 ;
        RECT 142.490 116.220 142.750 116.540 ;
        RECT 143.410 116.220 143.670 116.540 ;
        RECT 140.650 115.540 140.910 115.860 ;
        RECT 141.110 115.540 141.370 115.860 ;
        RECT 139.730 114.520 139.990 114.840 ;
        RECT 139.730 113.500 139.990 113.820 ;
        RECT 139.270 113.160 139.530 113.480 ;
        RECT 139.330 102.940 139.470 113.160 ;
        RECT 139.270 102.620 139.530 102.940 ;
        RECT 139.790 102.600 139.930 113.500 ;
        RECT 141.170 104.980 141.310 115.540 ;
        RECT 141.110 104.660 141.370 104.980 ;
        RECT 141.630 103.190 141.770 116.220 ;
        RECT 143.470 114.500 143.610 116.220 ;
        RECT 143.410 114.180 143.670 114.500 ;
        RECT 142.030 113.500 142.290 113.820 ;
        RECT 142.090 109.400 142.230 113.500 ;
        RECT 142.490 110.840 142.750 111.100 ;
        RECT 142.490 110.780 143.150 110.840 ;
        RECT 142.550 110.700 143.150 110.780 ;
        RECT 142.030 109.080 142.290 109.400 ;
        RECT 142.090 105.660 142.230 109.080 ;
        RECT 142.030 105.340 142.290 105.660 ;
        RECT 142.030 103.190 142.290 103.280 ;
        RECT 141.630 103.050 142.290 103.190 ;
        RECT 142.030 102.960 142.290 103.050 ;
        RECT 139.730 102.280 139.990 102.600 ;
        RECT 141.110 102.280 141.370 102.600 ;
        RECT 139.790 98.520 139.930 102.280 ;
        RECT 141.170 101.240 141.310 102.280 ;
        RECT 141.110 100.920 141.370 101.240 ;
        RECT 139.730 98.200 139.990 98.520 ;
        RECT 141.170 98.180 141.310 100.920 ;
        RECT 141.570 99.220 141.830 99.540 ;
        RECT 141.110 97.860 141.370 98.180 ;
        RECT 139.730 97.520 139.990 97.840 ;
        RECT 139.790 95.800 139.930 97.520 ;
        RECT 140.180 96.305 140.460 96.675 ;
        RECT 138.810 95.480 139.070 95.800 ;
        RECT 139.730 95.480 139.990 95.800 ;
        RECT 137.430 95.140 137.690 95.460 ;
        RECT 138.350 94.800 138.610 95.120 ;
        RECT 137.430 94.690 137.690 94.780 ;
        RECT 137.030 94.550 137.690 94.690 ;
        RECT 137.430 94.460 137.690 94.550 ;
        RECT 136.050 89.020 136.310 89.340 ;
        RECT 138.410 88.400 138.550 94.800 ;
        RECT 140.250 94.780 140.390 96.305 ;
        RECT 141.630 95.460 141.770 99.220 ;
        RECT 141.570 95.140 141.830 95.460 ;
        RECT 143.010 94.780 143.150 110.700 ;
        RECT 143.470 108.720 143.610 114.180 ;
        RECT 144.390 114.160 144.530 116.560 ;
        RECT 145.250 114.520 145.510 114.840 ;
        RECT 144.330 113.840 144.590 114.160 ;
        RECT 144.780 113.305 145.060 113.675 ;
        RECT 144.790 113.160 145.050 113.305 ;
        RECT 144.790 110.275 145.050 110.420 ;
        RECT 144.780 109.905 145.060 110.275 ;
        RECT 143.410 108.400 143.670 108.720 ;
        RECT 144.790 107.380 145.050 107.700 ;
        RECT 144.850 106.875 144.990 107.380 ;
        RECT 144.780 106.505 145.060 106.875 ;
        RECT 143.870 102.960 144.130 103.280 ;
        RECT 143.930 99.540 144.070 102.960 ;
        RECT 144.330 101.940 144.590 102.260 ;
        RECT 143.870 99.220 144.130 99.540 ;
        RECT 143.930 98.520 144.070 99.220 ;
        RECT 143.870 98.200 144.130 98.520 ;
        RECT 144.390 96.420 144.530 101.940 ;
        RECT 145.310 100.560 145.450 114.520 ;
        RECT 147.090 105.000 147.350 105.320 ;
        RECT 145.250 100.240 145.510 100.560 ;
        RECT 144.790 96.500 145.050 96.820 ;
        RECT 143.930 96.280 144.530 96.420 ;
        RECT 140.190 94.460 140.450 94.780 ;
        RECT 142.030 94.635 142.290 94.780 ;
        RECT 142.020 94.265 142.300 94.635 ;
        RECT 142.950 94.460 143.210 94.780 ;
        RECT 142.950 93.780 143.210 94.100 ;
        RECT 140.650 88.680 140.910 89.000 ;
        RECT 134.210 88.000 134.470 88.320 ;
        RECT 137.490 88.260 138.550 88.400 ;
        RECT 134.270 86.550 134.410 88.000 ;
        RECT 137.490 86.550 137.630 88.260 ;
        RECT 140.710 86.550 140.850 88.680 ;
        RECT 143.010 88.320 143.150 93.780 ;
        RECT 142.950 88.000 143.210 88.320 ;
        RECT 143.930 86.550 144.070 96.280 ;
        RECT 144.850 89.000 144.990 96.500 ;
        RECT 144.790 88.680 145.050 89.000 ;
        RECT 147.150 86.550 147.290 105.000 ;
        RECT 147.680 104.310 147.820 124.500 ;
        RECT 147.975 104.770 148.130 143.850 ;
        RECT 147.975 104.615 148.285 104.770 ;
        RECT 147.620 103.990 147.880 104.310 ;
        RECT 147.510 103.060 147.900 103.540 ;
        RECT 50.480 82.550 50.760 86.550 ;
        RECT 53.700 82.930 53.980 86.550 ;
        RECT 56.920 83.660 57.200 86.550 ;
        RECT 56.880 83.290 57.250 83.660 ;
        RECT 53.670 82.650 54.010 82.930 ;
        RECT 53.700 82.550 53.980 82.650 ;
        RECT 56.920 82.550 57.200 83.290 ;
        RECT 60.140 82.550 60.420 86.550 ;
        RECT 63.360 82.550 63.640 86.550 ;
        RECT 66.580 82.550 66.860 86.550 ;
        RECT 69.800 82.550 70.080 86.550 ;
        RECT 73.020 82.550 73.300 86.550 ;
        RECT 76.240 82.550 76.520 86.550 ;
        RECT 79.460 82.550 79.740 86.550 ;
        RECT 82.680 82.550 82.960 86.550 ;
        RECT 85.900 82.550 86.180 86.550 ;
        RECT 89.120 82.550 89.400 86.550 ;
        RECT 92.340 82.550 92.620 86.550 ;
        RECT 95.560 82.550 95.840 86.550 ;
        RECT 98.780 82.550 99.060 86.550 ;
        RECT 102.000 82.550 102.280 86.550 ;
        RECT 105.220 82.550 105.500 86.550 ;
        RECT 108.440 82.550 108.720 86.550 ;
        RECT 111.660 82.550 111.940 86.550 ;
        RECT 114.880 82.550 115.160 86.550 ;
        RECT 118.100 82.550 118.380 86.550 ;
        RECT 121.320 82.550 121.600 86.550 ;
        RECT 124.540 82.550 124.820 86.550 ;
        RECT 127.760 82.550 128.040 86.550 ;
        RECT 130.980 82.550 131.260 86.550 ;
        RECT 134.200 82.550 134.480 86.550 ;
        RECT 137.420 82.550 137.700 86.550 ;
        RECT 140.640 82.550 140.920 86.550 ;
        RECT 143.860 82.550 144.140 86.550 ;
        RECT 147.080 82.550 147.360 86.550 ;
        RECT 147.625 85.690 147.775 103.060 ;
        RECT 147.570 85.370 147.830 85.690 ;
        RECT 148.130 85.065 148.285 104.615 ;
        RECT 147.935 84.855 148.285 85.065 ;
        RECT 147.935 84.805 148.255 84.855 ;
        RECT 148.535 84.450 148.745 165.035 ;
        RECT 149.160 164.160 149.840 164.810 ;
        RECT 148.510 84.130 148.770 84.450 ;
        RECT 149.370 83.690 149.630 164.160 ;
        RECT 151.465 162.195 151.695 170.940 ;
        RECT 151.465 161.965 152.705 162.195 ;
        RECT 151.090 161.230 151.770 161.420 ;
        RECT 151.090 160.950 152.200 161.230 ;
        RECT 151.090 160.770 151.770 160.950 ;
        RECT 151.235 157.840 151.735 158.010 ;
        RECT 150.120 157.540 151.735 157.840 ;
        RECT 150.120 152.170 150.420 157.540 ;
        RECT 151.235 157.370 151.735 157.540 ;
        RECT 150.690 153.970 151.370 154.620 ;
        RECT 150.170 105.780 150.370 152.170 ;
        RECT 148.790 83.430 149.630 83.690 ;
        RECT 149.830 105.580 150.370 105.780 ;
        RECT 149.830 83.100 150.030 105.580 ;
        RECT 150.310 104.660 150.570 104.980 ;
        RECT 150.370 86.550 150.510 104.660 ;
        RECT 149.660 82.960 150.030 83.100 ;
        RECT 149.410 82.730 150.030 82.960 ;
        RECT 149.410 82.700 149.730 82.730 ;
        RECT 150.300 82.550 150.580 86.550 ;
        RECT 150.950 82.370 151.130 153.970 ;
        RECT 151.920 141.850 152.200 160.950 ;
        RECT 152.475 142.560 152.705 161.965 ;
        RECT 152.460 142.240 152.720 142.560 ;
        RECT 151.920 141.570 152.390 141.850 ;
        RECT 151.505 140.370 151.785 141.010 ;
        RECT 55.590 82.190 151.130 82.370 ;
        RECT 31.160 81.710 54.180 81.990 ;
        RECT 11.840 81.000 36.790 81.280 ;
        RECT 37.570 81.110 53.520 81.390 ;
        RECT 36.510 80.800 36.790 81.000 ;
        RECT 36.510 80.520 52.790 80.800 ;
        RECT 52.510 28.470 52.790 80.520 ;
        RECT 53.240 29.080 53.520 81.110 ;
        RECT 53.900 29.630 54.180 81.710 ;
        RECT 54.720 75.210 55.380 75.920 ;
        RECT 55.590 67.550 55.770 82.190 ;
        RECT 151.555 82.000 151.735 140.370 ;
        RECT 57.130 81.820 151.735 82.000 ;
        RECT 55.550 67.230 55.810 67.550 ;
        RECT 57.130 67.510 57.310 81.820 ;
        RECT 152.110 81.570 152.390 141.570 ;
        RECT 148.310 81.545 152.390 81.570 ;
        RECT 58.660 81.320 152.390 81.545 ;
        RECT 58.660 67.535 58.885 81.320 ;
        RECT 148.310 81.290 152.390 81.320 ;
        RECT 149.410 81.000 149.730 81.030 ;
        RECT 60.190 80.800 149.730 81.000 ;
        RECT 60.190 67.590 60.390 80.800 ;
        RECT 149.410 80.770 149.730 80.800 ;
        RECT 148.820 80.510 149.080 80.540 ;
        RECT 61.770 80.250 149.080 80.510 ;
        RECT 57.090 67.190 57.350 67.510 ;
        RECT 58.645 67.215 58.905 67.535 ;
        RECT 60.160 67.270 60.420 67.590 ;
        RECT 61.770 67.180 62.030 80.250 ;
        RECT 148.820 80.220 149.080 80.250 ;
        RECT 148.270 79.965 148.590 79.990 ;
        RECT 63.385 79.755 148.590 79.965 ;
        RECT 63.385 67.550 63.595 79.755 ;
        RECT 148.270 79.730 148.590 79.755 ;
        RECT 147.785 79.355 148.105 79.395 ;
        RECT 64.975 79.180 148.105 79.355 ;
        RECT 63.360 67.230 63.620 67.550 ;
        RECT 64.975 67.515 65.150 79.180 ;
        RECT 147.785 79.135 148.105 79.180 ;
        RECT 152.430 78.815 152.750 78.830 ;
        RECT 66.515 78.585 152.750 78.815 ;
        RECT 64.935 67.195 65.195 67.515 ;
        RECT 66.515 67.510 66.745 78.585 ;
        RECT 152.430 78.570 152.750 78.585 ;
        RECT 151.770 78.145 152.090 78.155 ;
        RECT 67.745 77.910 152.090 78.145 ;
        RECT 66.500 67.190 66.760 67.510 ;
        RECT 54.840 65.000 55.160 65.870 ;
        RECT 54.830 63.970 55.160 65.000 ;
        RECT 56.510 64.980 56.830 65.860 ;
        RECT 54.830 62.210 55.140 63.970 ;
        RECT 56.490 63.960 56.830 64.980 ;
        RECT 58.070 63.960 58.390 65.860 ;
        RECT 59.610 64.970 59.930 65.870 ;
        RECT 59.590 63.970 59.930 64.970 ;
        RECT 61.200 64.780 61.520 65.890 ;
        RECT 56.490 62.320 56.800 63.960 ;
        RECT 54.830 62.050 55.050 62.210 ;
        RECT 55.300 62.050 55.840 62.190 ;
        RECT 54.830 59.960 55.840 62.050 ;
        RECT 54.870 59.940 55.840 59.960 ;
        RECT 56.490 62.000 57.300 62.320 ;
        RECT 58.070 62.190 58.380 63.960 ;
        RECT 56.490 59.940 57.220 62.000 ;
        RECT 55.230 59.850 55.840 59.940 ;
        RECT 56.770 59.910 57.220 59.940 ;
        RECT 56.800 59.880 57.170 59.910 ;
        RECT 58.070 59.900 58.740 62.190 ;
        RECT 59.590 62.170 59.900 63.970 ;
        RECT 61.160 63.540 61.530 64.780 ;
        RECT 62.760 64.770 63.080 65.860 ;
        RECT 64.350 64.810 64.670 65.880 ;
        RECT 65.950 65.120 66.230 65.870 ;
        RECT 62.740 63.540 63.110 64.770 ;
        RECT 61.160 62.530 63.130 63.540 ;
        RECT 61.160 62.200 61.530 62.530 ;
        RECT 62.740 62.230 63.110 62.530 ;
        RECT 59.590 59.930 60.250 62.170 ;
        RECT 58.190 59.840 58.740 59.900 ;
        RECT 59.700 59.820 60.250 59.930 ;
        RECT 61.160 59.850 61.710 62.200 ;
        RECT 62.640 59.880 63.190 62.230 ;
        RECT 64.350 62.220 64.700 64.810 ;
        RECT 65.930 62.230 66.230 65.120 ;
        RECT 64.090 59.970 64.700 62.220 ;
        RECT 64.090 59.870 64.640 59.970 ;
        RECT 65.590 59.940 66.230 62.230 ;
        RECT 65.590 59.880 66.140 59.940 ;
        RECT 54.840 47.520 56.480 48.440 ;
        RECT 60.060 43.960 60.450 46.750 ;
        RECT 62.295 46.195 62.665 49.555 ;
        RECT 63.510 43.960 63.960 46.740 ;
        RECT 60.060 41.300 63.960 43.960 ;
        RECT 58.760 38.320 59.280 39.870 ;
        RECT 60.060 38.760 60.450 41.300 ;
        RECT 63.510 38.800 63.960 41.300 ;
        RECT 65.980 39.110 66.370 39.145 ;
        RECT 67.745 39.110 67.980 77.910 ;
        RECT 151.770 77.895 152.090 77.910 ;
        RECT 147.360 77.555 147.680 77.610 ;
        RECT 68.345 77.405 147.680 77.555 ;
        RECT 68.345 76.500 68.495 77.405 ;
        RECT 147.360 77.350 147.680 77.405 ;
        RECT 68.290 76.180 68.550 76.500 ;
        RECT 88.610 76.490 89.830 76.580 ;
        RECT 82.370 76.000 143.470 76.490 ;
        RECT 82.360 75.500 143.470 76.000 ;
        RECT 82.360 75.230 83.300 75.500 ;
        RECT 80.420 71.980 80.810 74.770 ;
        RECT 82.340 74.300 83.310 75.230 ;
        RECT 83.870 71.980 84.320 74.760 ;
        RECT 87.810 74.490 88.440 75.330 ;
        RECT 73.540 71.020 79.680 71.900 ;
        RECT 80.420 69.320 84.320 71.980 ;
        RECT 80.420 66.780 80.810 69.320 ;
        RECT 83.870 66.820 84.320 69.320 ;
        RECT 73.390 65.430 74.340 66.540 ;
        RECT 75.120 65.720 75.860 65.740 ;
        RECT 75.120 65.430 76.720 65.720 ;
        RECT 85.290 65.430 86.080 65.500 ;
        RECT 75.110 64.730 86.080 65.430 ;
        RECT 75.120 64.420 76.720 64.730 ;
        RECT 85.290 64.640 86.080 64.730 ;
        RECT 75.120 64.390 75.860 64.420 ;
        RECT 77.870 63.020 78.540 63.370 ;
        RECT 77.870 61.470 83.450 63.020 ;
        RECT 77.870 60.990 78.550 61.470 ;
        RECT 72.920 58.850 73.780 59.530 ;
        RECT 77.870 59.490 78.540 60.990 ;
        RECT 85.930 60.570 86.690 61.300 ;
        RECT 77.870 59.460 78.270 59.490 ;
        RECT 78.440 57.960 79.970 58.710 ;
        RECT 88.610 58.110 89.830 75.500 ;
        RECT 97.330 75.240 98.270 75.500 ;
        RECT 95.400 71.960 95.790 74.750 ;
        RECT 97.310 74.310 98.280 75.240 ;
        RECT 98.850 71.960 99.300 74.740 ;
        RECT 93.840 69.110 94.790 70.220 ;
        RECT 95.400 69.300 99.300 71.960 ;
        RECT 95.400 66.760 95.790 69.300 ;
        RECT 98.850 66.800 99.300 69.300 ;
        RECT 90.100 65.700 90.840 65.720 ;
        RECT 90.100 65.410 91.700 65.700 ;
        RECT 100.270 65.410 101.060 65.480 ;
        RECT 90.090 64.710 101.060 65.410 ;
        RECT 90.100 64.400 91.700 64.710 ;
        RECT 100.270 64.620 101.060 64.710 ;
        RECT 90.100 64.370 90.840 64.400 ;
        RECT 92.850 63.000 93.520 63.350 ;
        RECT 92.850 61.450 98.430 63.000 ;
        RECT 92.850 60.970 93.530 61.450 ;
        RECT 92.850 59.470 93.520 60.970 ;
        RECT 100.790 60.420 101.550 61.150 ;
        RECT 92.850 59.440 93.250 59.470 ;
        RECT 103.680 58.110 104.900 75.500 ;
        RECT 112.290 75.260 113.230 75.500 ;
        RECT 110.410 71.960 110.800 74.750 ;
        RECT 112.240 74.270 113.270 75.260 ;
        RECT 113.860 71.960 114.310 74.740 ;
        RECT 108.870 68.840 109.820 69.950 ;
        RECT 110.410 69.300 114.310 71.960 ;
        RECT 110.410 66.760 110.800 69.300 ;
        RECT 113.860 66.800 114.310 69.300 ;
        RECT 105.110 65.700 105.850 65.720 ;
        RECT 105.110 65.410 106.710 65.700 ;
        RECT 115.280 65.410 116.070 65.480 ;
        RECT 105.100 64.710 116.070 65.410 ;
        RECT 105.110 64.400 106.710 64.710 ;
        RECT 115.280 64.620 116.070 64.710 ;
        RECT 105.110 64.370 105.850 64.400 ;
        RECT 107.860 63.000 108.530 63.350 ;
        RECT 107.860 61.450 113.440 63.000 ;
        RECT 107.860 60.970 108.540 61.450 ;
        RECT 107.860 59.470 108.530 60.970 ;
        RECT 115.710 60.460 116.470 61.190 ;
        RECT 107.860 59.440 108.260 59.470 ;
        RECT 118.710 58.110 119.930 75.500 ;
        RECT 127.380 75.230 128.320 75.500 ;
        RECT 125.420 71.960 125.810 74.750 ;
        RECT 127.350 74.380 128.320 75.230 ;
        RECT 128.870 71.960 129.320 74.740 ;
        RECT 123.720 69.010 124.920 70.310 ;
        RECT 125.420 69.300 129.320 71.960 ;
        RECT 125.420 66.760 125.810 69.300 ;
        RECT 128.870 66.800 129.320 69.300 ;
        RECT 120.120 65.700 120.860 65.720 ;
        RECT 120.120 65.410 121.720 65.700 ;
        RECT 130.290 65.410 131.080 65.480 ;
        RECT 120.110 64.710 131.080 65.410 ;
        RECT 120.120 64.400 121.720 64.710 ;
        RECT 130.290 64.620 131.080 64.710 ;
        RECT 120.120 64.370 120.860 64.400 ;
        RECT 122.870 63.000 123.540 63.350 ;
        RECT 122.870 61.450 128.450 63.000 ;
        RECT 122.870 60.970 123.550 61.450 ;
        RECT 122.870 59.470 123.540 60.970 ;
        RECT 130.800 60.450 131.560 61.180 ;
        RECT 122.870 59.440 123.270 59.470 ;
        RECT 133.570 58.110 134.790 75.500 ;
        RECT 142.330 75.230 143.270 75.500 ;
        RECT 140.410 71.960 140.800 74.750 ;
        RECT 142.330 74.380 143.300 75.230 ;
        RECT 143.860 71.960 144.310 74.740 ;
        RECT 138.850 69.210 139.790 70.290 ;
        RECT 140.410 69.300 144.310 71.960 ;
        RECT 140.410 66.760 140.800 69.300 ;
        RECT 143.860 66.800 144.310 69.300 ;
        RECT 135.110 65.700 135.850 65.720 ;
        RECT 135.110 65.410 136.710 65.700 ;
        RECT 145.280 65.410 146.070 65.480 ;
        RECT 135.100 64.710 146.070 65.410 ;
        RECT 135.110 64.400 136.710 64.710 ;
        RECT 145.280 64.620 146.070 64.710 ;
        RECT 135.110 64.370 135.850 64.400 ;
        RECT 137.860 63.000 138.530 63.350 ;
        RECT 137.860 61.450 143.440 63.000 ;
        RECT 137.860 60.970 138.540 61.450 ;
        RECT 137.860 59.470 138.530 60.970 ;
        RECT 145.810 60.500 146.620 61.150 ;
        RECT 137.860 59.440 138.260 59.470 ;
        RECT 82.300 57.170 143.280 58.110 ;
        RECT 73.220 56.420 74.080 57.100 ;
        RECT 82.300 57.010 143.390 57.170 ;
        RECT 82.340 56.190 83.200 57.010 ;
        RECT 73.520 52.480 74.380 53.160 ;
        RECT 80.420 52.970 80.810 55.760 ;
        RECT 82.340 55.270 83.320 56.190 ;
        RECT 82.350 55.260 83.320 55.270 ;
        RECT 83.870 52.970 84.320 55.750 ;
        RECT 87.810 55.510 88.440 56.580 ;
        RECT 73.220 50.860 74.080 50.920 ;
        RECT 78.850 50.860 79.830 50.970 ;
        RECT 73.220 50.410 79.830 50.860 ;
        RECT 73.220 50.240 74.080 50.410 ;
        RECT 78.850 50.240 79.830 50.410 ;
        RECT 80.420 50.310 84.320 52.970 ;
        RECT 80.420 47.770 80.810 50.310 ;
        RECT 83.870 47.810 84.320 50.310 ;
        RECT 73.530 46.940 74.490 47.750 ;
        RECT 75.120 46.710 75.860 46.730 ;
        RECT 75.120 46.420 76.720 46.710 ;
        RECT 85.290 46.420 86.080 46.490 ;
        RECT 75.110 45.720 86.080 46.420 ;
        RECT 75.120 45.410 76.720 45.720 ;
        RECT 85.290 45.630 86.080 45.720 ;
        RECT 75.120 45.380 75.860 45.410 ;
        RECT 73.450 44.210 74.410 45.020 ;
        RECT 77.870 44.010 78.540 44.360 ;
        RECT 77.870 42.460 83.450 44.010 ;
        RECT 73.400 41.250 74.040 42.230 ;
        RECT 77.870 41.980 78.550 42.460 ;
        RECT 77.870 40.480 78.540 41.980 ;
        RECT 85.790 41.490 86.550 42.220 ;
        RECT 77.870 40.450 78.270 40.480 ;
        RECT 65.980 38.875 67.980 39.110 ;
        RECT 65.980 38.845 66.370 38.875 ;
        RECT 58.760 37.800 69.300 38.320 ;
        RECT 73.410 38.070 74.070 39.000 ;
        RECT 78.240 38.970 79.770 39.720 ;
        RECT 88.610 39.150 89.830 57.010 ;
        RECT 97.390 56.110 98.250 57.010 ;
        RECT 95.400 52.960 95.790 55.750 ;
        RECT 97.370 55.370 98.250 56.110 ;
        RECT 97.370 55.360 98.140 55.370 ;
        RECT 98.850 52.960 99.300 55.740 ;
        RECT 93.910 49.700 94.660 50.630 ;
        RECT 95.400 50.300 99.300 52.960 ;
        RECT 95.400 47.760 95.790 50.300 ;
        RECT 98.850 47.800 99.300 50.300 ;
        RECT 90.100 46.700 90.840 46.720 ;
        RECT 90.100 46.410 91.700 46.700 ;
        RECT 100.270 46.410 101.060 46.480 ;
        RECT 90.090 45.710 101.060 46.410 ;
        RECT 90.100 45.400 91.700 45.710 ;
        RECT 100.270 45.620 101.060 45.710 ;
        RECT 90.100 45.370 90.840 45.400 ;
        RECT 92.850 44.000 93.520 44.350 ;
        RECT 92.850 42.450 98.430 44.000 ;
        RECT 92.850 41.970 93.530 42.450 ;
        RECT 92.850 40.470 93.520 41.970 ;
        RECT 100.810 41.550 101.570 42.280 ;
        RECT 92.850 40.440 93.250 40.470 ;
        RECT 103.680 39.150 104.900 57.010 ;
        RECT 110.440 52.960 110.830 55.750 ;
        RECT 112.510 55.390 113.370 57.010 ;
        RECT 112.510 55.380 113.280 55.390 ;
        RECT 113.890 52.960 114.340 55.740 ;
        RECT 109.000 49.780 109.750 50.710 ;
        RECT 110.440 50.300 114.340 52.960 ;
        RECT 110.440 47.760 110.830 50.300 ;
        RECT 113.890 47.800 114.340 50.300 ;
        RECT 105.140 46.700 105.880 46.720 ;
        RECT 105.140 46.410 106.740 46.700 ;
        RECT 115.310 46.410 116.100 46.480 ;
        RECT 105.130 45.710 116.100 46.410 ;
        RECT 105.140 45.400 106.740 45.710 ;
        RECT 115.310 45.620 116.100 45.710 ;
        RECT 105.140 45.370 105.880 45.400 ;
        RECT 107.890 44.000 108.560 44.350 ;
        RECT 107.890 42.450 113.470 44.000 ;
        RECT 107.890 41.970 108.570 42.450 ;
        RECT 107.890 40.470 108.560 41.970 ;
        RECT 115.860 41.550 116.620 42.280 ;
        RECT 107.890 40.440 108.290 40.470 ;
        RECT 118.710 39.150 119.930 57.010 ;
        RECT 125.420 52.960 125.810 55.750 ;
        RECT 127.420 55.370 128.280 57.010 ;
        RECT 127.420 55.340 128.260 55.370 ;
        RECT 128.870 52.960 129.320 55.740 ;
        RECT 123.970 49.790 124.720 50.720 ;
        RECT 125.420 50.300 129.320 52.960 ;
        RECT 125.420 47.760 125.810 50.300 ;
        RECT 128.870 47.800 129.320 50.300 ;
        RECT 120.120 46.700 120.860 46.720 ;
        RECT 120.120 46.410 121.720 46.700 ;
        RECT 130.290 46.410 131.080 46.480 ;
        RECT 120.110 45.710 131.080 46.410 ;
        RECT 120.120 45.400 121.720 45.710 ;
        RECT 130.290 45.620 131.080 45.710 ;
        RECT 120.120 45.370 120.860 45.400 ;
        RECT 122.870 44.000 123.540 44.350 ;
        RECT 122.870 42.450 128.450 44.000 ;
        RECT 122.870 41.970 123.550 42.450 ;
        RECT 122.870 40.470 123.540 41.970 ;
        RECT 130.880 41.540 131.640 42.270 ;
        RECT 122.870 40.440 123.270 40.470 ;
        RECT 133.570 39.150 134.790 57.010 ;
        RECT 142.450 56.180 143.390 57.010 ;
        RECT 140.430 52.990 140.820 55.780 ;
        RECT 142.440 55.500 143.390 56.180 ;
        RECT 142.440 55.460 143.210 55.500 ;
        RECT 143.880 52.990 144.330 55.770 ;
        RECT 138.960 49.690 139.710 50.620 ;
        RECT 140.430 50.330 144.330 52.990 ;
        RECT 140.430 47.790 140.820 50.330 ;
        RECT 143.880 47.830 144.330 50.330 ;
        RECT 135.130 46.730 135.870 46.750 ;
        RECT 135.130 46.440 136.730 46.730 ;
        RECT 145.300 46.440 146.090 46.510 ;
        RECT 135.120 45.740 146.090 46.440 ;
        RECT 135.130 45.430 136.730 45.740 ;
        RECT 145.300 45.650 146.090 45.740 ;
        RECT 135.130 45.400 135.870 45.430 ;
        RECT 137.880 44.030 138.550 44.380 ;
        RECT 137.880 42.480 143.460 44.030 ;
        RECT 137.880 42.000 138.560 42.480 ;
        RECT 137.880 40.500 138.550 42.000 ;
        RECT 146.050 41.520 146.510 42.000 ;
        RECT 137.880 40.470 138.280 40.500 ;
        RECT 54.760 37.410 55.500 37.720 ;
        RECT 64.930 37.410 65.720 37.480 ;
        RECT 54.750 36.710 65.720 37.410 ;
        RECT 54.760 36.370 55.500 36.710 ;
        RECT 64.930 36.620 65.720 36.710 ;
        RECT 65.995 33.020 66.355 33.030 ;
        RECT 65.990 32.740 66.360 33.020 ;
        RECT 65.995 32.730 66.355 32.740 ;
        RECT 61.450 29.920 63.100 30.760 ;
        RECT 53.900 29.350 61.000 29.630 ;
        RECT 53.240 28.800 60.250 29.080 ;
        RECT 52.510 28.190 59.540 28.470 ;
        RECT 59.260 16.820 59.540 28.190 ;
        RECT 59.970 17.360 60.250 28.800 ;
        RECT 60.720 17.940 61.000 29.350 ;
        RECT 61.440 28.210 62.560 28.980 ;
        RECT 62.950 27.660 65.580 28.010 ;
        RECT 62.950 27.460 63.220 27.660 ;
        RECT 62.540 23.580 63.220 27.460 ;
        RECT 62.930 23.360 63.210 23.580 ;
        RECT 62.930 23.040 66.070 23.360 ;
        RECT 63.810 23.030 64.140 23.040 ;
        RECT 64.770 23.030 65.100 23.040 ;
        RECT 65.730 23.030 66.060 23.040 ;
        RECT 61.490 22.050 62.670 22.710 ;
        RECT 68.780 22.520 69.300 37.800 ;
        RECT 82.440 37.680 143.290 39.150 ;
        RECT 82.520 37.120 83.260 37.680 ;
        RECT 73.430 35.870 74.170 36.000 ;
        RECT 78.990 35.870 79.730 36.010 ;
        RECT 73.430 35.340 79.730 35.870 ;
        RECT 73.430 35.220 74.170 35.340 ;
        RECT 78.990 35.230 79.730 35.340 ;
        RECT 80.460 33.960 80.850 36.750 ;
        RECT 82.510 36.470 83.260 37.120 ;
        RECT 88.370 36.880 89.700 37.330 ;
        RECT 97.450 37.110 98.190 37.680 ;
        RECT 112.420 37.110 113.160 37.680 ;
        RECT 82.510 36.430 83.250 36.470 ;
        RECT 83.910 33.960 84.360 36.740 ;
        RECT 93.840 34.020 94.620 35.010 ;
        RECT 73.250 32.130 73.920 33.000 ;
        RECT 80.460 31.300 84.360 33.960 ;
        RECT 73.390 28.900 74.060 29.770 ;
        RECT 80.460 28.760 80.850 31.300 ;
        RECT 83.910 28.800 84.360 31.300 ;
        RECT 95.400 33.960 95.790 36.750 ;
        RECT 97.450 36.460 98.210 37.110 ;
        RECT 97.470 36.420 98.210 36.460 ;
        RECT 98.850 33.960 99.300 36.740 ;
        RECT 110.410 33.960 110.800 36.750 ;
        RECT 112.390 36.350 113.220 37.110 ;
        RECT 127.460 37.100 128.200 37.680 ;
        RECT 113.860 33.960 114.310 36.740 ;
        RECT 95.400 31.300 99.300 33.960 ;
        RECT 108.990 32.970 109.770 33.960 ;
        RECT 95.400 28.760 95.790 31.300 ;
        RECT 98.850 28.800 99.300 31.300 ;
        RECT 110.410 31.300 114.310 33.960 ;
        RECT 125.450 33.960 125.840 36.750 ;
        RECT 127.460 36.390 128.250 37.100 ;
        RECT 127.480 36.380 128.250 36.390 ;
        RECT 128.900 33.960 129.350 36.740 ;
        RECT 123.860 31.790 124.640 32.780 ;
        RECT 110.410 28.760 110.800 31.300 ;
        RECT 113.860 28.800 114.310 31.300 ;
        RECT 125.450 31.300 129.350 33.960 ;
        RECT 125.450 28.760 125.840 31.300 ;
        RECT 128.900 28.800 129.350 31.300 ;
        RECT 75.160 27.700 75.900 27.720 ;
        RECT 90.100 27.700 90.840 27.720 ;
        RECT 105.110 27.700 105.850 27.720 ;
        RECT 120.150 27.700 120.890 27.720 ;
        RECT 71.660 26.460 72.560 27.360 ;
        RECT 73.230 26.610 73.900 27.480 ;
        RECT 75.160 27.410 76.760 27.700 ;
        RECT 85.330 27.410 86.120 27.480 ;
        RECT 90.100 27.410 91.700 27.700 ;
        RECT 100.270 27.410 101.060 27.480 ;
        RECT 105.110 27.410 106.710 27.700 ;
        RECT 115.280 27.410 116.070 27.480 ;
        RECT 120.150 27.410 121.750 27.700 ;
        RECT 130.320 27.410 131.110 27.480 ;
        RECT 75.150 26.710 86.120 27.410 ;
        RECT 90.090 26.710 101.060 27.410 ;
        RECT 105.100 26.710 116.070 27.410 ;
        RECT 120.140 26.710 131.110 27.410 ;
        RECT 75.160 26.400 76.760 26.710 ;
        RECT 85.330 26.620 86.120 26.710 ;
        RECT 90.100 26.400 91.700 26.710 ;
        RECT 100.270 26.620 101.060 26.710 ;
        RECT 105.110 26.400 106.710 26.710 ;
        RECT 115.280 26.620 116.070 26.710 ;
        RECT 120.150 26.400 121.750 26.710 ;
        RECT 130.320 26.620 131.110 26.710 ;
        RECT 75.160 26.370 75.900 26.400 ;
        RECT 90.100 26.370 90.840 26.400 ;
        RECT 105.110 26.370 105.850 26.400 ;
        RECT 120.150 26.370 120.890 26.400 ;
        RECT 61.490 21.710 63.330 22.050 ;
        RECT 64.050 22.000 69.300 22.520 ;
        RECT 61.490 21.700 62.670 21.710 ;
        RECT 63.060 21.500 63.290 21.710 ;
        RECT 63.060 21.180 65.570 21.500 ;
        RECT 63.060 19.860 63.290 21.180 ;
        RECT 64.280 21.170 64.610 21.180 ;
        RECT 65.240 21.170 65.570 21.180 ;
        RECT 63.060 19.520 66.060 19.860 ;
        RECT 68.780 19.750 69.300 22.000 ;
        RECT 77.910 25.000 78.580 25.350 ;
        RECT 92.850 25.000 93.520 25.350 ;
        RECT 107.860 25.000 108.530 25.350 ;
        RECT 122.900 25.000 123.570 25.350 ;
        RECT 77.910 23.450 83.490 25.000 ;
        RECT 92.850 23.450 98.430 25.000 ;
        RECT 107.860 23.450 113.440 25.000 ;
        RECT 122.900 23.450 128.480 25.000 ;
        RECT 77.910 22.970 78.590 23.450 ;
        RECT 77.910 21.470 78.580 22.970 ;
        RECT 85.870 22.650 86.300 23.060 ;
        RECT 92.850 22.970 93.530 23.450 ;
        RECT 92.850 21.470 93.520 22.970 ;
        RECT 100.870 22.600 101.300 23.010 ;
        RECT 107.860 22.970 108.540 23.450 ;
        RECT 107.860 21.470 108.530 22.970 ;
        RECT 115.990 22.570 116.420 22.980 ;
        RECT 122.900 22.970 123.580 23.450 ;
        RECT 122.900 21.470 123.570 22.970 ;
        RECT 130.980 22.580 131.410 22.990 ;
        RECT 77.910 21.440 78.310 21.470 ;
        RECT 92.850 21.440 93.250 21.470 ;
        RECT 107.860 21.440 108.260 21.470 ;
        RECT 122.900 21.440 123.300 21.470 ;
        RECT 78.230 20.010 79.810 20.710 ;
        RECT 133.975 19.750 134.790 37.680 ;
        RECT 142.440 37.140 143.180 37.680 ;
        RECT 140.410 33.960 140.800 36.750 ;
        RECT 142.420 36.420 143.190 37.140 ;
        RECT 143.860 33.960 144.310 36.740 ;
        RECT 140.410 31.300 144.310 33.960 ;
        RECT 139.010 30.260 139.790 31.250 ;
        RECT 140.410 28.760 140.800 31.300 ;
        RECT 143.860 28.800 144.310 31.300 ;
        RECT 135.110 27.700 135.850 27.720 ;
        RECT 135.110 27.410 136.710 27.700 ;
        RECT 145.280 27.410 146.070 27.480 ;
        RECT 135.100 26.710 146.070 27.410 ;
        RECT 135.110 26.400 136.710 26.710 ;
        RECT 145.280 26.620 146.070 26.710 ;
        RECT 135.110 26.370 135.850 26.400 ;
        RECT 137.860 25.000 138.530 25.350 ;
        RECT 137.860 23.450 143.440 25.000 ;
        RECT 137.860 22.970 138.540 23.450 ;
        RECT 137.860 21.470 138.530 22.970 ;
        RECT 137.860 21.440 138.260 21.470 ;
        RECT 68.780 19.725 152.585 19.750 ;
        RECT 61.560 18.380 63.320 19.020 ;
        RECT 68.550 18.960 152.585 19.725 ;
        RECT 68.835 18.935 152.585 18.960 ;
        RECT 85.895 17.940 86.285 17.950 ;
        RECT 60.720 17.660 86.285 17.940 ;
        RECT 116.010 17.780 116.410 18.180 ;
        RECT 85.895 17.650 86.285 17.660 ;
        RECT 100.885 17.360 101.275 17.370 ;
        RECT 59.970 17.080 101.275 17.360 ;
        RECT 100.885 17.070 101.275 17.080 ;
        RECT 130.985 16.820 131.375 16.830 ;
        RECT 59.260 16.540 131.375 16.820 ;
        RECT 130.985 16.530 131.375 16.540 ;
        RECT 151.770 3.360 152.585 18.935 ;
        RECT 151.630 2.310 152.720 3.360 ;
      LAYER met3 ;
        RECT 33.300 224.810 33.870 225.380 ;
        RECT 63.670 225.040 64.140 225.560 ;
        RECT 71.910 224.880 72.380 225.650 ;
        RECT 74.640 224.940 75.350 225.590 ;
        RECT 77.450 224.860 78.030 225.470 ;
        RECT 80.190 224.880 80.730 225.500 ;
        RECT 82.970 224.880 83.500 225.440 ;
        RECT 85.640 224.780 86.400 225.570 ;
        RECT 88.520 225.060 89.040 225.620 ;
        RECT 91.220 224.940 91.850 225.620 ;
        RECT 94.150 225.040 94.450 225.340 ;
        RECT 126.980 224.850 127.530 225.540 ;
        RECT 95.920 224.500 96.240 224.540 ;
        RECT 97.940 224.500 98.320 224.510 ;
        RECT 95.920 224.200 98.320 224.500 ;
        RECT 95.920 224.160 96.240 224.200 ;
        RECT 97.940 224.190 98.320 224.200 ;
        RECT 74.550 223.720 83.690 224.020 ;
        RECT 125.800 223.980 126.280 224.400 ;
        RECT 74.550 223.430 74.850 223.720 ;
        RECT 61.740 223.200 74.850 223.430 ;
        RECT 83.390 223.430 83.690 223.720 ;
        RECT 125.880 223.430 126.180 223.980 ;
        RECT 61.740 223.130 74.830 223.200 ;
        RECT 61.740 222.800 62.040 223.130 ;
        RECT 79.420 222.970 80.080 223.360 ;
        RECT 83.390 223.130 126.180 223.430 ;
        RECT 16.015 222.500 62.040 222.800 ;
        RECT 127.140 222.630 127.440 224.850 ;
        RECT 129.900 224.680 130.460 225.340 ;
        RECT 132.450 224.710 133.340 225.530 ;
        RECT 135.310 224.910 136.020 225.580 ;
        RECT 137.900 224.820 138.550 225.640 ;
        RECT 140.930 224.920 141.430 225.440 ;
        RECT 143.830 224.860 144.150 225.240 ;
        RECT 16.015 220.645 16.315 222.500 ;
        RECT 62.800 222.330 127.440 222.630 ;
        RECT 32.180 221.930 35.010 222.050 ;
        RECT 62.800 221.930 63.100 222.330 ;
        RECT 63.845 222.000 64.195 222.330 ;
        RECT 130.010 222.000 130.310 224.680 ;
        RECT 136.550 224.335 137.150 224.410 ;
        RECT 143.840 224.335 144.140 224.860 ;
        RECT 136.550 224.035 144.140 224.335 ;
        RECT 136.550 223.930 137.150 224.035 ;
        RECT 63.845 221.985 130.310 222.000 ;
        RECT 16.650 221.740 63.100 221.930 ;
        RECT 16.650 221.630 32.500 221.740 ;
        RECT 34.680 221.630 63.100 221.740 ;
        RECT 63.870 221.700 130.310 221.985 ;
        RECT 15.990 220.295 16.340 220.645 ;
        RECT 11.750 198.640 15.750 198.790 ;
        RECT 16.650 198.640 16.950 221.630 ;
        RECT 32.800 221.105 34.380 221.435 ;
        RECT 36.100 218.385 37.680 218.715 ;
        RECT 32.800 215.665 34.380 215.995 ;
        RECT 36.100 212.945 37.680 213.275 ;
        RECT 32.800 210.225 34.380 210.555 ;
        RECT 36.100 207.505 37.680 207.835 ;
        RECT 32.800 204.785 34.380 205.115 ;
        RECT 36.100 202.065 37.680 202.395 ;
        RECT 96.915 201.360 97.245 201.375 ;
        RECT 102.435 201.360 102.765 201.375 ;
        RECT 96.915 201.060 102.765 201.360 ;
        RECT 96.915 201.045 97.245 201.060 ;
        RECT 102.435 201.045 102.765 201.060 ;
        RECT 38.955 200.000 39.285 200.015 ;
        RECT 52.295 200.000 52.625 200.015 ;
        RECT 65.635 200.000 65.965 200.015 ;
        RECT 38.955 199.700 65.965 200.000 ;
        RECT 38.955 199.685 39.285 199.700 ;
        RECT 52.295 199.685 52.625 199.700 ;
        RECT 65.635 199.685 65.965 199.700 ;
        RECT 32.800 199.345 34.380 199.675 ;
        RECT 18.715 198.640 19.045 198.655 ;
        RECT 11.750 198.340 19.045 198.640 ;
        RECT 11.750 198.190 15.750 198.340 ;
        RECT 18.715 198.325 19.045 198.340 ;
        RECT 90.475 198.640 90.805 198.655 ;
        RECT 101.055 198.640 101.385 198.655 ;
        RECT 105.655 198.640 105.985 198.655 ;
        RECT 90.475 198.340 105.985 198.640 ;
        RECT 90.475 198.325 90.805 198.340 ;
        RECT 101.055 198.325 101.385 198.340 ;
        RECT 105.655 198.325 105.985 198.340 ;
        RECT 95.995 197.960 96.325 197.975 ;
        RECT 105.195 197.960 105.525 197.975 ;
        RECT 95.995 197.660 105.525 197.960 ;
        RECT 95.995 197.645 96.325 197.660 ;
        RECT 105.195 197.645 105.525 197.660 ;
        RECT 36.100 196.625 37.680 196.955 ;
        RECT 32.800 193.905 34.380 194.235 ;
        RECT 36.100 191.185 37.680 191.515 ;
        RECT 32.800 188.465 34.380 188.795 ;
        RECT 36.100 185.745 37.680 186.075 ;
        RECT 131.875 185.040 132.205 185.055 ;
        RECT 134.635 185.040 134.965 185.055 ;
        RECT 131.875 184.740 134.965 185.040 ;
        RECT 131.875 184.725 132.205 184.740 ;
        RECT 134.635 184.725 134.965 184.740 ;
        RECT 32.800 183.025 34.380 183.355 ;
        RECT 128.655 181.640 128.985 181.655 ;
        RECT 141.995 181.640 142.325 181.655 ;
        RECT 128.655 181.340 142.325 181.640 ;
        RECT 128.655 181.325 128.985 181.340 ;
        RECT 141.995 181.325 142.325 181.340 ;
        RECT 130.495 180.960 130.825 180.975 ;
        RECT 137.855 180.960 138.185 180.975 ;
        RECT 130.495 180.660 138.185 180.960 ;
        RECT 130.495 180.645 130.825 180.660 ;
        RECT 137.855 180.645 138.185 180.660 ;
        RECT 36.100 180.305 37.680 180.635 ;
        RECT 118.535 179.600 118.865 179.615 ;
        RECT 133.255 179.600 133.585 179.615 ;
        RECT 118.535 179.300 133.585 179.600 ;
        RECT 118.535 179.285 118.865 179.300 ;
        RECT 133.255 179.285 133.585 179.300 ;
        RECT 119.455 178.920 119.785 178.935 ;
        RECT 130.955 178.920 131.285 178.935 ;
        RECT 119.455 178.620 131.285 178.920 ;
        RECT 119.455 178.605 119.785 178.620 ;
        RECT 130.955 178.605 131.285 178.620 ;
        RECT 107.495 178.250 107.825 178.255 ;
        RECT 107.495 178.240 108.080 178.250 ;
        RECT 129.575 178.240 129.905 178.255 ;
        RECT 132.335 178.240 132.665 178.255 ;
        RECT 107.495 177.940 108.280 178.240 ;
        RECT 129.575 177.940 132.665 178.240 ;
        RECT 107.495 177.930 108.080 177.940 ;
        RECT 107.495 177.925 107.825 177.930 ;
        RECT 129.575 177.925 129.905 177.940 ;
        RECT 132.335 177.925 132.665 177.940 ;
        RECT 32.800 177.585 34.380 177.915 ;
        RECT 107.955 177.560 108.285 177.575 ;
        RECT 107.740 177.245 108.285 177.560 ;
        RECT 125.895 177.560 126.225 177.575 ;
        RECT 136.475 177.560 136.805 177.575 ;
        RECT 125.895 177.260 136.805 177.560 ;
        RECT 125.895 177.245 126.225 177.260 ;
        RECT 136.475 177.245 136.805 177.260 ;
        RECT 107.740 176.215 108.040 177.245 ;
        RECT 120.375 176.880 120.705 176.895 ;
        RECT 123.595 176.880 123.925 176.895 ;
        RECT 132.795 176.880 133.125 176.895 ;
        RECT 120.375 176.580 133.125 176.880 ;
        RECT 120.375 176.565 120.705 176.580 ;
        RECT 123.595 176.565 123.925 176.580 ;
        RECT 132.795 176.565 133.125 176.580 ;
        RECT 107.740 175.900 108.285 176.215 ;
        RECT 107.955 175.885 108.285 175.900 ;
        RECT 105.195 175.520 105.525 175.535 ;
        RECT 110.255 175.520 110.585 175.535 ;
        RECT 105.195 175.220 110.585 175.520 ;
        RECT 105.195 175.205 105.525 175.220 ;
        RECT 110.255 175.205 110.585 175.220 ;
        RECT 36.100 174.865 37.680 175.195 ;
        RECT 145.215 174.840 145.545 174.855 ;
        RECT 148.755 174.840 152.755 174.990 ;
        RECT 145.215 174.540 152.755 174.840 ;
        RECT 145.215 174.525 145.545 174.540 ;
        RECT 148.755 174.390 152.755 174.540 ;
        RECT 130.955 174.160 131.285 174.175 ;
        RECT 133.255 174.160 133.585 174.175 ;
        RECT 130.955 173.860 133.585 174.160 ;
        RECT 130.955 173.845 131.285 173.860 ;
        RECT 133.255 173.845 133.585 173.860 ;
        RECT 131.875 173.480 132.205 173.495 ;
        RECT 132.540 173.480 132.920 173.490 ;
        RECT 131.875 173.180 132.920 173.480 ;
        RECT 131.875 173.165 132.205 173.180 ;
        RECT 132.540 173.170 132.920 173.180 ;
        RECT 32.800 172.145 34.380 172.475 ;
        RECT 151.220 171.590 151.930 171.630 ;
        RECT 124.055 171.440 124.385 171.455 ;
        RECT 127.735 171.440 128.065 171.455 ;
        RECT 124.055 171.140 128.065 171.440 ;
        RECT 124.055 171.125 124.385 171.140 ;
        RECT 127.735 171.125 128.065 171.140 ;
        RECT 144.755 171.440 145.085 171.455 ;
        RECT 148.755 171.440 152.755 171.590 ;
        RECT 144.755 171.140 152.755 171.440 ;
        RECT 144.755 171.125 145.085 171.140 ;
        RECT 148.755 170.990 152.755 171.140 ;
        RECT 151.220 170.940 151.930 170.990 ;
        RECT 36.100 169.425 37.680 169.755 ;
        RECT 88.175 168.720 88.505 168.735 ;
        RECT 99.675 168.720 100.005 168.735 ;
        RECT 88.175 168.420 100.005 168.720 ;
        RECT 88.175 168.405 88.505 168.420 ;
        RECT 99.675 168.405 100.005 168.420 ;
        RECT 144.755 168.040 145.085 168.055 ;
        RECT 148.730 168.040 152.755 168.190 ;
        RECT 144.755 167.740 152.755 168.040 ;
        RECT 144.755 167.725 145.085 167.740 ;
        RECT 148.730 167.590 152.755 167.740 ;
        RECT 148.730 167.540 149.410 167.590 ;
        RECT 121.295 167.360 121.625 167.375 ;
        RECT 132.335 167.360 132.665 167.375 ;
        RECT 121.295 167.060 132.665 167.360 ;
        RECT 121.295 167.045 121.625 167.060 ;
        RECT 132.335 167.045 132.665 167.060 ;
        RECT 32.800 166.705 34.380 167.035 ;
        RECT 112.555 166.000 112.885 166.015 ;
        RECT 118.995 166.000 119.325 166.015 ;
        RECT 125.895 166.000 126.225 166.015 ;
        RECT 132.335 166.010 132.665 166.015 ;
        RECT 132.335 166.000 132.920 166.010 ;
        RECT 112.555 165.700 132.920 166.000 ;
        RECT 112.555 165.685 112.885 165.700 ;
        RECT 118.995 165.685 119.325 165.700 ;
        RECT 125.895 165.685 126.225 165.700 ;
        RECT 132.335 165.690 132.920 165.700 ;
        RECT 132.335 165.685 132.665 165.690 ;
        RECT 149.160 164.790 149.840 164.810 ;
        RECT 116.235 164.650 116.565 164.655 ;
        RECT 115.980 164.640 116.565 164.650 ;
        RECT 115.780 164.340 116.565 164.640 ;
        RECT 115.980 164.330 116.565 164.340 ;
        RECT 116.235 164.325 116.565 164.330 ;
        RECT 144.755 164.640 145.085 164.655 ;
        RECT 148.755 164.640 152.755 164.790 ;
        RECT 144.755 164.340 152.755 164.640 ;
        RECT 144.755 164.325 145.085 164.340 ;
        RECT 36.100 163.985 37.680 164.315 ;
        RECT 148.755 164.190 152.755 164.340 ;
        RECT 149.160 164.160 149.840 164.190 ;
        RECT 130.495 163.280 130.825 163.295 ;
        RECT 135.555 163.280 135.885 163.295 ;
        RECT 144.755 163.280 145.085 163.295 ;
        RECT 130.495 162.980 145.085 163.280 ;
        RECT 130.495 162.965 130.825 162.980 ;
        RECT 135.555 162.965 135.885 162.980 ;
        RECT 144.755 162.965 145.085 162.980 ;
        RECT 116.235 162.600 116.565 162.615 ;
        RECT 120.375 162.600 120.705 162.615 ;
        RECT 130.955 162.600 131.285 162.615 ;
        RECT 116.235 162.300 131.285 162.600 ;
        RECT 116.235 162.285 116.565 162.300 ;
        RECT 120.375 162.285 120.705 162.300 ;
        RECT 130.955 162.285 131.285 162.300 ;
        RECT 15.955 161.920 16.285 161.935 ;
        RECT 15.740 161.605 16.285 161.920 ;
        RECT 15.740 161.390 16.040 161.605 ;
        RECT 11.750 160.940 16.040 161.390 ;
        RECT 32.800 161.265 34.380 161.595 ;
        RECT 151.090 161.390 151.770 161.420 ;
        RECT 107.955 161.250 108.285 161.255 ;
        RECT 107.700 161.240 108.285 161.250 ;
        RECT 107.500 160.940 108.285 161.240 ;
        RECT 11.750 160.790 15.750 160.940 ;
        RECT 107.700 160.930 108.285 160.940 ;
        RECT 107.955 160.925 108.285 160.930 ;
        RECT 142.915 161.240 143.245 161.255 ;
        RECT 148.755 161.240 152.755 161.390 ;
        RECT 142.915 160.940 152.755 161.240 ;
        RECT 142.915 160.925 143.245 160.940 ;
        RECT 148.755 160.790 152.755 160.940 ;
        RECT 151.090 160.770 151.770 160.790 ;
        RECT 118.995 160.560 119.325 160.575 ;
        RECT 143.375 160.560 143.705 160.575 ;
        RECT 118.995 160.260 143.705 160.560 ;
        RECT 118.995 160.245 119.325 160.260 ;
        RECT 143.375 160.245 143.705 160.260 ;
        RECT 122.215 159.210 122.545 159.215 ;
        RECT 122.215 159.200 122.800 159.210 ;
        RECT 122.215 158.900 123.000 159.200 ;
        RECT 122.215 158.890 122.800 158.900 ;
        RECT 122.215 158.885 122.545 158.890 ;
        RECT 11.730 158.430 15.730 158.560 ;
        RECT 36.100 158.545 37.680 158.875 ;
        RECT 11.730 157.960 16.280 158.430 ;
        RECT 14.940 157.930 16.280 157.960 ;
        RECT 121.295 157.840 121.625 157.855 ;
        RECT 130.035 157.840 130.365 157.855 ;
        RECT 121.295 157.540 130.365 157.840 ;
        RECT 121.295 157.525 121.625 157.540 ;
        RECT 130.035 157.525 130.365 157.540 ;
        RECT 145.215 157.840 145.545 157.855 ;
        RECT 148.755 157.840 152.755 157.990 ;
        RECT 145.215 157.540 152.755 157.840 ;
        RECT 145.215 157.525 145.545 157.540 ;
        RECT 148.755 157.390 152.755 157.540 ;
        RECT 32.800 155.825 34.380 156.155 ;
        RECT 150.690 154.590 151.370 154.620 ;
        RECT 144.755 154.440 145.085 154.455 ;
        RECT 148.755 154.440 152.755 154.590 ;
        RECT 144.755 154.140 152.755 154.440 ;
        RECT 144.755 154.125 145.085 154.140 ;
        RECT 148.755 153.990 152.755 154.140 ;
        RECT 150.690 153.970 151.370 153.990 ;
        RECT 36.100 153.105 37.680 153.435 ;
        RECT 115.775 151.730 116.105 151.735 ;
        RECT 115.775 151.720 116.360 151.730 ;
        RECT 115.550 151.420 116.360 151.720 ;
        RECT 115.775 151.410 116.360 151.420 ;
        RECT 115.775 151.405 116.105 151.410 ;
        RECT 142.915 151.040 143.245 151.055 ;
        RECT 148.755 151.040 152.755 151.190 ;
        RECT 142.915 150.740 152.755 151.040 ;
        RECT 142.915 150.725 143.245 150.740 ;
        RECT 32.800 150.385 34.380 150.715 ;
        RECT 148.755 150.590 152.755 150.740 ;
        RECT 36.100 147.665 37.680 147.995 ;
        RECT 144.755 147.640 145.085 147.655 ;
        RECT 148.755 147.640 152.755 147.790 ;
        RECT 144.755 147.340 152.755 147.640 ;
        RECT 144.755 147.325 145.085 147.340 ;
        RECT 148.755 147.190 152.755 147.340 ;
        RECT 32.800 144.945 34.380 145.275 ;
        RECT 13.480 144.390 14.180 144.420 ;
        RECT 11.750 144.240 15.750 144.390 ;
        RECT 19.175 144.240 19.505 144.255 ;
        RECT 11.750 143.940 19.505 144.240 ;
        RECT 11.750 143.790 15.750 143.940 ;
        RECT 19.175 143.925 19.505 143.940 ;
        RECT 142.915 144.240 143.245 144.255 ;
        RECT 147.800 144.240 148.310 144.300 ;
        RECT 148.755 144.240 152.755 144.390 ;
        RECT 142.915 143.940 152.755 144.240 ;
        RECT 142.915 143.925 143.245 143.940 ;
        RECT 147.800 143.850 148.310 143.940 ;
        RECT 148.755 143.790 152.755 143.940 ;
        RECT 13.480 143.750 14.180 143.790 ;
        RECT 36.100 142.225 37.680 142.555 ;
        RECT 15.955 141.520 16.285 141.535 ;
        RECT 15.740 141.205 16.285 141.520 ;
        RECT 15.740 140.990 16.040 141.205 ;
        RECT 11.750 140.540 16.040 140.990 ;
        RECT 144.755 140.840 145.085 140.855 ;
        RECT 148.755 140.840 152.755 140.990 ;
        RECT 144.755 140.540 152.755 140.840 ;
        RECT 11.750 140.390 15.750 140.540 ;
        RECT 144.755 140.525 145.085 140.540 ;
        RECT 148.755 140.390 152.755 140.540 ;
        RECT 32.800 139.505 34.380 139.835 ;
        RECT 15.460 137.590 16.060 137.620 ;
        RECT 11.750 136.990 16.900 137.590 ;
        RECT 144.755 137.440 145.085 137.455 ;
        RECT 148.755 137.440 152.755 137.590 ;
        RECT 144.755 137.140 152.755 137.440 ;
        RECT 144.755 137.125 145.085 137.140 ;
        RECT 15.460 136.960 16.060 136.990 ;
        RECT 12.230 135.630 12.700 136.200 ;
        RECT 16.450 135.645 16.755 136.990 ;
        RECT 36.100 136.785 37.680 137.115 ;
        RECT 148.755 136.990 152.755 137.140 ;
        RECT 16.450 135.340 16.960 135.645 ;
        RECT 15.955 134.720 16.285 134.735 ;
        RECT 15.740 134.405 16.285 134.720 ;
        RECT 14.805 134.190 15.395 134.195 ;
        RECT 15.740 134.190 16.040 134.405 ;
        RECT 11.750 133.740 16.040 134.190 ;
        RECT 11.750 133.590 15.750 133.740 ;
        RECT 14.805 133.545 15.395 133.590 ;
        RECT 11.750 130.640 15.750 130.790 ;
        RECT 11.750 130.190 16.040 130.640 ;
        RECT 15.740 129.975 16.040 130.190 ;
        RECT 15.740 129.660 16.285 129.975 ;
        RECT 15.955 129.645 16.285 129.660 ;
        RECT 15.955 127.920 16.285 127.935 ;
        RECT 15.740 127.605 16.285 127.920 ;
        RECT 15.740 127.390 16.040 127.605 ;
        RECT 11.750 126.940 16.040 127.390 ;
        RECT 11.750 126.790 15.750 126.940 ;
        RECT 15.465 125.295 15.845 125.305 ;
        RECT 16.655 125.295 16.960 135.340 ;
        RECT 32.800 134.065 34.380 134.395 ;
        RECT 144.755 134.040 145.085 134.055 ;
        RECT 148.755 134.040 152.755 134.190 ;
        RECT 144.755 133.740 152.755 134.040 ;
        RECT 144.755 133.725 145.085 133.740 ;
        RECT 148.755 133.590 152.755 133.740 ;
        RECT 36.100 131.345 37.680 131.675 ;
        RECT 111.175 130.640 111.505 130.655 ;
        RECT 129.115 130.640 129.445 130.655 ;
        RECT 111.175 130.340 129.445 130.640 ;
        RECT 111.175 130.325 111.505 130.340 ;
        RECT 129.115 130.325 129.445 130.340 ;
        RECT 142.915 130.640 143.245 130.655 ;
        RECT 148.755 130.640 152.755 130.790 ;
        RECT 142.915 130.340 152.755 130.640 ;
        RECT 142.915 130.325 143.245 130.340 ;
        RECT 148.755 130.190 152.755 130.340 ;
        RECT 32.800 128.625 34.380 128.955 ;
        RECT 113.475 127.240 113.805 127.255 ;
        RECT 122.420 127.240 122.800 127.250 ;
        RECT 113.475 126.940 122.800 127.240 ;
        RECT 113.475 126.925 113.805 126.940 ;
        RECT 122.420 126.930 122.800 126.940 ;
        RECT 144.755 127.240 145.085 127.255 ;
        RECT 148.755 127.240 152.755 127.390 ;
        RECT 144.755 126.940 152.755 127.240 ;
        RECT 144.755 126.925 145.085 126.940 ;
        RECT 148.755 126.790 152.755 126.940 ;
        RECT 36.100 125.905 37.680 126.235 ;
        RECT 15.465 124.990 16.960 125.295 ;
        RECT 15.465 124.985 15.845 124.990 ;
        RECT 108.415 124.520 108.745 124.535 ;
        RECT 136.935 124.520 137.265 124.535 ;
        RECT 108.415 124.220 137.265 124.520 ;
        RECT 108.415 124.205 108.745 124.220 ;
        RECT 136.935 124.205 137.265 124.220 ;
        RECT 11.750 123.980 15.750 123.990 ;
        RECT 11.750 123.840 16.180 123.980 ;
        RECT 21.015 123.840 21.345 123.855 ;
        RECT 11.750 123.540 21.345 123.840 ;
        RECT 11.750 123.390 16.180 123.540 ;
        RECT 21.015 123.525 21.345 123.540 ;
        RECT 142.915 123.840 143.245 123.855 ;
        RECT 148.755 123.840 152.755 123.990 ;
        RECT 142.915 123.540 152.755 123.840 ;
        RECT 142.915 123.525 143.245 123.540 ;
        RECT 15.480 123.380 16.180 123.390 ;
        RECT 32.800 123.185 34.380 123.515 ;
        RECT 148.755 123.390 152.755 123.540 ;
        RECT 11.750 120.440 15.750 120.590 ;
        RECT 36.100 120.465 37.680 120.795 ;
        RECT 144.755 120.440 145.085 120.455 ;
        RECT 148.755 120.440 152.755 120.590 ;
        RECT 11.750 119.990 16.040 120.440 ;
        RECT 144.755 120.140 152.755 120.440 ;
        RECT 144.755 120.125 145.085 120.140 ;
        RECT 148.755 119.990 152.755 120.140 ;
        RECT 15.590 119.775 16.040 119.990 ;
        RECT 15.590 119.680 16.285 119.775 ;
        RECT 15.590 119.440 16.300 119.680 ;
        RECT 15.760 119.280 16.300 119.440 ;
        RECT 32.800 117.745 34.380 118.075 ;
        RECT 12.100 117.190 12.780 117.210 ;
        RECT 11.750 117.040 15.750 117.190 ;
        RECT 20.095 117.040 20.425 117.055 ;
        RECT 11.750 116.740 20.425 117.040 ;
        RECT 11.750 116.590 15.750 116.740 ;
        RECT 20.095 116.725 20.425 116.740 ;
        RECT 142.915 117.040 143.245 117.055 ;
        RECT 148.755 117.040 152.755 117.190 ;
        RECT 142.915 116.740 152.755 117.040 ;
        RECT 142.915 116.725 143.245 116.740 ;
        RECT 148.755 116.590 152.755 116.740 ;
        RECT 12.100 116.560 12.780 116.590 ;
        RECT 36.100 115.025 37.680 115.355 ;
        RECT 11.750 113.640 15.750 113.790 ;
        RECT 144.755 113.640 145.085 113.655 ;
        RECT 148.755 113.640 152.755 113.790 ;
        RECT 11.750 113.190 16.040 113.640 ;
        RECT 144.755 113.340 152.755 113.640 ;
        RECT 144.755 113.325 145.085 113.340 ;
        RECT 148.755 113.190 152.755 113.340 ;
        RECT 15.740 112.975 16.040 113.190 ;
        RECT 15.740 112.660 16.285 112.975 ;
        RECT 15.955 112.645 16.285 112.660 ;
        RECT 32.800 112.305 34.380 112.635 ;
        RECT 14.700 110.390 15.750 110.490 ;
        RECT 11.750 110.240 15.750 110.390 ;
        RECT 18.255 110.240 18.585 110.255 ;
        RECT 11.750 109.940 18.585 110.240 ;
        RECT 11.750 109.790 15.750 109.940 ;
        RECT 18.255 109.925 18.585 109.940 ;
        RECT 144.755 110.240 145.085 110.255 ;
        RECT 148.755 110.240 152.755 110.390 ;
        RECT 144.755 109.940 152.755 110.240 ;
        RECT 144.755 109.925 145.085 109.940 ;
        RECT 14.700 109.720 15.750 109.790 ;
        RECT 36.100 109.585 37.680 109.915 ;
        RECT 148.755 109.790 152.755 109.940 ;
        RECT 11.750 106.840 15.750 106.990 ;
        RECT 32.800 106.865 34.380 107.195 ;
        RECT 18.255 106.840 18.585 106.855 ;
        RECT 11.750 106.540 18.585 106.840 ;
        RECT 11.750 106.390 15.750 106.540 ;
        RECT 18.255 106.525 18.585 106.540 ;
        RECT 144.755 106.840 145.085 106.855 ;
        RECT 148.755 106.840 152.755 106.990 ;
        RECT 144.755 106.540 152.755 106.840 ;
        RECT 144.755 106.525 145.085 106.540 ;
        RECT 148.755 106.390 152.755 106.540 ;
        RECT 36.100 104.145 37.680 104.475 ;
        RECT 11.750 103.440 15.750 103.590 ;
        RECT 16.875 103.440 17.205 103.455 ;
        RECT 70.695 103.450 71.025 103.455 ;
        RECT 70.695 103.440 71.280 103.450 ;
        RECT 71.615 103.440 71.945 103.455 ;
        RECT 11.750 103.140 17.205 103.440 ;
        RECT 70.470 103.140 71.945 103.440 ;
        RECT 11.750 102.990 15.750 103.140 ;
        RECT 16.875 103.125 17.205 103.140 ;
        RECT 70.695 103.130 71.280 103.140 ;
        RECT 70.695 103.125 71.025 103.130 ;
        RECT 71.615 103.125 71.945 103.140 ;
        RECT 147.400 102.720 147.900 103.540 ;
        RECT 32.800 101.425 34.380 101.755 ;
        RECT 36.100 98.705 37.680 99.035 ;
        RECT 90.015 98.000 90.345 98.015 ;
        RECT 92.775 98.000 93.105 98.015 ;
        RECT 94.155 98.000 94.485 98.015 ;
        RECT 90.015 97.700 94.485 98.000 ;
        RECT 90.015 97.685 90.345 97.700 ;
        RECT 92.775 97.685 93.105 97.700 ;
        RECT 94.155 97.685 94.485 97.700 ;
        RECT 131.415 96.640 131.745 96.655 ;
        RECT 136.475 96.640 136.805 96.655 ;
        RECT 140.155 96.640 140.485 96.655 ;
        RECT 131.415 96.340 140.485 96.640 ;
        RECT 131.415 96.325 131.745 96.340 ;
        RECT 136.475 96.325 136.805 96.340 ;
        RECT 140.155 96.325 140.485 96.340 ;
        RECT 32.800 95.985 34.380 96.315 ;
        RECT 71.155 95.290 71.485 95.295 ;
        RECT 70.900 95.280 71.485 95.290 ;
        RECT 70.900 94.980 71.710 95.280 ;
        RECT 70.900 94.970 71.485 94.980 ;
        RECT 71.155 94.965 71.485 94.970 ;
        RECT 135.095 94.600 135.425 94.615 ;
        RECT 141.995 94.600 142.325 94.615 ;
        RECT 135.095 94.300 142.325 94.600 ;
        RECT 135.095 94.285 135.425 94.300 ;
        RECT 141.995 94.285 142.325 94.300 ;
        RECT 36.100 93.265 37.680 93.595 ;
        RECT 12.910 91.970 13.390 92.520 ;
        RECT 47.170 91.730 47.890 92.230 ;
        RECT 34.845 91.170 35.195 91.195 ;
        RECT 38.940 91.170 39.320 91.180 ;
        RECT 34.845 90.870 39.320 91.170 ;
        RECT 34.845 90.845 35.195 90.870 ;
        RECT 38.940 90.860 39.320 90.870 ;
        RECT 43.920 89.980 45.010 90.620 ;
        RECT 40.730 89.320 41.420 89.770 ;
        RECT 24.685 88.940 25.035 88.965 ;
        RECT 38.980 88.940 39.360 88.950 ;
        RECT 24.685 88.640 39.360 88.940 ;
        RECT 24.685 88.615 25.035 88.640 ;
        RECT 38.980 88.630 39.360 88.640 ;
        RECT 16.450 88.310 16.830 88.320 ;
        RECT 38.900 88.310 39.280 88.320 ;
        RECT 16.450 88.010 39.280 88.310 ;
        RECT 16.450 88.000 16.830 88.010 ;
        RECT 38.900 88.000 39.280 88.010 ;
        RECT 50.360 87.680 51.620 88.180 ;
        RECT 15.025 87.220 15.375 87.245 ;
        RECT 38.980 87.220 39.300 87.260 ;
        RECT 15.025 86.920 39.300 87.220 ;
        RECT 15.025 86.895 15.375 86.920 ;
        RECT 38.980 86.880 39.300 86.920 ;
        RECT 15.740 86.590 16.120 86.595 ;
        RECT 15.740 86.285 38.380 86.590 ;
        RECT 15.740 86.275 16.120 86.285 ;
        RECT 38.075 86.135 38.380 86.285 ;
        RECT 38.930 86.135 39.310 86.145 ;
        RECT 18.180 85.850 18.640 85.910 ;
        RECT 18.180 85.550 35.890 85.850 ;
        RECT 38.075 85.830 39.310 86.135 ;
        RECT 38.930 85.825 39.310 85.830 ;
        RECT 18.180 85.490 18.640 85.550 ;
        RECT 35.590 85.240 35.890 85.550 ;
        RECT 38.730 85.240 39.110 85.250 ;
        RECT 35.590 84.940 39.110 85.240 ;
        RECT 38.730 84.930 39.110 84.940 ;
        RECT 32.750 75.210 55.380 75.920 ;
        RECT 53.360 48.450 54.180 75.210 ;
        RECT 87.730 74.420 89.710 75.370 ;
        RECT 93.840 70.090 94.790 70.220 ;
        RECT 73.580 70.030 94.790 70.090 ;
        RECT 73.400 69.110 94.790 70.030 ;
        RECT 73.400 69.090 94.700 69.110 ;
        RECT 73.400 66.540 74.370 69.090 ;
        RECT 108.870 69.030 109.820 69.950 ;
        RECT 108.740 68.840 109.820 69.030 ;
        RECT 123.720 69.010 124.920 70.310 ;
        RECT 138.850 69.210 139.790 70.290 ;
        RECT 74.740 68.780 78.950 68.790 ;
        RECT 108.740 68.780 109.810 68.840 ;
        RECT 74.740 68.750 109.810 68.780 ;
        RECT 73.390 65.430 74.370 66.540 ;
        RECT 73.400 65.420 74.370 65.430 ;
        RECT 74.730 67.820 109.810 68.750 ;
        RECT 74.730 67.810 78.950 67.820 ;
        RECT 74.730 65.380 75.870 67.810 ;
        RECT 93.390 67.640 109.810 67.820 ;
        RECT 123.850 67.420 124.790 69.010 ;
        RECT 78.680 67.410 92.800 67.420 ;
        RECT 76.490 67.160 92.800 67.410 ;
        RECT 112.200 67.160 124.790 67.420 ;
        RECT 76.490 66.310 124.790 67.160 ;
        RECT 61.480 62.530 63.130 63.540 ;
        RECT 74.730 59.550 75.900 65.380 ;
        RECT 72.960 59.530 75.900 59.550 ;
        RECT 72.920 58.900 75.900 59.530 ;
        RECT 72.920 58.850 73.780 58.900 ;
        RECT 75.100 58.860 75.900 58.900 ;
        RECT 76.510 58.270 76.930 66.310 ;
        RECT 78.680 66.190 124.790 66.310 ;
        RECT 123.850 66.150 124.790 66.190 ;
        RECT 139.020 65.790 139.710 69.210 ;
        RECT 77.570 65.770 139.710 65.790 ;
        RECT 77.560 65.210 139.710 65.770 ;
        RECT 73.270 57.890 76.940 58.270 ;
        RECT 73.290 57.100 74.000 57.890 ;
        RECT 73.220 56.420 74.080 57.100 ;
        RECT 73.520 53.050 74.380 53.160 ;
        RECT 77.560 53.050 78.090 65.210 ;
        RECT 85.930 60.570 86.690 61.300 ;
        RECT 100.790 60.420 101.550 61.150 ;
        RECT 115.710 60.460 116.470 61.190 ;
        RECT 130.800 60.450 131.560 61.180 ;
        RECT 145.810 60.500 146.620 61.150 ;
        RECT 88.940 58.830 90.130 59.010 ;
        RECT 78.440 57.960 79.970 58.710 ;
        RECT 88.860 58.040 90.130 58.830 ;
        RECT 88.940 57.950 90.130 58.040 ;
        RECT 89.040 56.480 90.020 57.950 ;
        RECT 87.740 55.550 90.020 56.480 ;
        RECT 87.740 55.530 89.320 55.550 ;
        RECT 73.520 52.520 78.090 53.050 ;
        RECT 73.520 52.480 74.380 52.520 ;
        RECT 77.560 52.500 78.090 52.520 ;
        RECT 73.220 50.240 74.080 50.920 ;
        RECT 93.910 49.980 94.660 50.630 ;
        RECT 74.300 49.700 94.660 49.980 ;
        RECT 109.000 49.780 109.750 50.710 ;
        RECT 123.970 49.790 124.720 50.720 ;
        RECT 74.300 49.570 94.570 49.700 ;
        RECT 53.360 47.510 56.500 48.450 ;
        RECT 74.320 47.750 74.730 49.570 ;
        RECT 94.040 49.560 94.560 49.570 ;
        RECT 109.020 49.130 109.740 49.780 ;
        RECT 73.530 47.720 74.730 47.750 ;
        RECT 75.080 48.610 109.750 49.130 ;
        RECT 54.070 29.220 55.010 47.510 ;
        RECT 73.530 46.980 74.740 47.720 ;
        RECT 73.530 46.960 74.730 46.980 ;
        RECT 73.530 46.940 74.490 46.960 ;
        RECT 73.450 44.980 74.410 45.020 ;
        RECT 75.080 44.980 75.710 48.610 ;
        RECT 124.080 48.060 124.650 49.790 ;
        RECT 138.960 49.690 139.710 50.620 ;
        RECT 76.330 48.040 124.720 48.060 ;
        RECT 76.310 47.450 124.720 48.040 ;
        RECT 73.450 44.430 75.740 44.980 ;
        RECT 73.450 44.210 74.410 44.430 ;
        RECT 75.080 44.420 75.710 44.430 ;
        RECT 73.400 42.170 74.040 42.230 ;
        RECT 76.310 42.170 76.880 47.450 ;
        RECT 139.140 46.930 139.570 49.690 ;
        RECT 73.400 41.560 76.880 42.170 ;
        RECT 77.340 46.550 139.570 46.930 ;
        RECT 77.340 46.440 139.550 46.550 ;
        RECT 73.400 41.250 74.040 41.560 ;
        RECT 66.000 38.820 66.350 39.170 ;
        RECT 73.410 38.970 74.070 39.000 ;
        RECT 77.340 38.970 77.860 46.440 ;
        RECT 85.790 41.490 86.550 42.220 ;
        RECT 100.810 41.550 101.570 42.280 ;
        RECT 115.860 41.550 116.620 42.280 ;
        RECT 130.880 41.540 131.640 42.270 ;
        RECT 145.850 41.470 146.610 42.200 ;
        RECT 78.240 38.970 79.770 39.720 ;
        RECT 66.025 33.045 66.325 38.820 ;
        RECT 73.410 38.510 77.860 38.970 ;
        RECT 73.410 38.500 77.850 38.510 ;
        RECT 73.410 38.070 74.070 38.500 ;
        RECT 88.910 37.430 90.160 38.780 ;
        RECT 88.320 37.090 90.160 37.430 ;
        RECT 88.320 36.870 89.820 37.090 ;
        RECT 93.840 34.850 94.620 35.010 ;
        RECT 73.290 34.790 94.620 34.850 ;
        RECT 73.270 34.350 94.620 34.790 ;
        RECT 66.010 32.715 66.340 33.045 ;
        RECT 73.270 33.000 73.790 34.350 ;
        RECT 93.840 34.020 94.620 34.350 ;
        RECT 108.990 33.610 109.770 33.960 ;
        RECT 74.370 33.530 109.770 33.610 ;
        RECT 73.250 32.130 73.920 33.000 ;
        RECT 74.350 32.970 109.770 33.530 ;
        RECT 74.350 32.950 109.690 32.970 ;
        RECT 61.450 29.920 63.100 30.760 ;
        RECT 73.390 29.580 74.060 29.770 ;
        RECT 74.370 29.580 74.910 32.950 ;
        RECT 123.860 32.460 124.640 32.780 ;
        RECT 75.580 31.810 124.640 32.460 ;
        RECT 54.070 28.980 62.450 29.220 ;
        RECT 73.390 29.010 74.910 29.580 ;
        RECT 54.070 28.280 62.560 28.980 ;
        RECT 73.390 28.900 74.060 29.010 ;
        RECT 74.370 28.980 74.910 29.010 ;
        RECT 75.600 28.360 76.250 31.810 ;
        RECT 123.860 31.790 124.640 31.810 ;
        RECT 139.010 30.970 139.790 31.250 ;
        RECT 61.440 28.210 62.560 28.280 ;
        RECT 71.710 27.800 76.250 28.360 ;
        RECT 76.780 30.490 139.790 30.970 ;
        RECT 71.730 27.360 72.340 27.800 ;
        RECT 73.230 27.400 73.900 27.480 ;
        RECT 76.780 27.400 77.330 30.490 ;
        RECT 139.010 30.260 139.790 30.490 ;
        RECT 71.660 26.460 72.560 27.360 ;
        RECT 73.230 26.710 77.330 27.400 ;
        RECT 73.230 26.610 73.900 26.710 ;
        RECT 76.780 26.620 77.330 26.710 ;
        RECT 85.925 22.685 86.255 23.015 ;
        RECT 78.230 20.010 79.810 20.710 ;
        RECT 61.480 18.310 63.520 19.170 ;
        RECT 85.940 17.975 86.240 22.685 ;
        RECT 100.915 22.635 101.245 22.965 ;
        RECT 85.915 17.625 86.265 17.975 ;
        RECT 100.930 17.395 101.230 22.635 ;
        RECT 116.045 22.615 116.375 22.945 ;
        RECT 116.060 18.180 116.360 22.615 ;
        RECT 131.015 22.595 131.345 22.925 ;
        RECT 116.010 17.780 116.410 18.180 ;
        RECT 100.905 17.045 101.255 17.395 ;
        RECT 131.030 16.855 131.330 22.595 ;
        RECT 131.005 16.505 131.355 16.855 ;
        RECT 151.630 2.310 152.720 3.360 ;
      LAYER met4 ;
        RECT 30.670 225.200 30.970 225.760 ;
        RECT 33.430 225.380 33.730 225.760 ;
        RECT 33.300 225.200 33.870 225.380 ;
        RECT 36.190 225.200 36.490 225.760 ;
        RECT 38.950 225.200 39.250 225.760 ;
        RECT 41.710 225.200 42.010 225.760 ;
        RECT 44.470 225.200 44.770 225.760 ;
        RECT 47.230 225.200 47.530 225.760 ;
        RECT 49.990 225.200 50.290 225.760 ;
        RECT 30.670 224.900 52.750 225.200 ;
        RECT 53.050 224.900 55.510 225.200 ;
        RECT 55.810 224.900 58.270 225.200 ;
        RECT 30.670 224.760 30.970 224.900 ;
        RECT 33.300 224.810 33.870 224.900 ;
        RECT 33.430 224.760 33.730 224.810 ;
        RECT 36.190 224.760 36.490 224.900 ;
        RECT 38.950 224.760 39.250 224.900 ;
        RECT 41.710 224.760 42.010 224.900 ;
        RECT 44.470 224.760 44.770 224.900 ;
        RECT 47.230 224.760 47.530 224.900 ;
        RECT 49.990 224.760 50.290 224.900 ;
        RECT 61.330 224.760 61.370 225.190 ;
        RECT 63.670 225.040 63.790 225.560 ;
        RECT 64.090 225.040 64.140 225.560 ;
        RECT 61.070 224.310 61.370 224.760 ;
        RECT 12.970 224.010 61.370 224.310 ;
        RECT 66.520 224.760 66.550 225.445 ;
        RECT 69.120 224.760 69.310 225.340 ;
        RECT 69.610 224.760 69.720 225.340 ;
        RECT 71.910 224.880 72.070 225.650 ;
        RECT 72.370 224.880 72.380 225.650 ;
        RECT 74.640 224.940 74.830 225.590 ;
        RECT 75.130 224.940 75.350 225.590 ;
        RECT 77.450 224.860 77.590 225.470 ;
        RECT 77.890 224.860 78.030 225.470 ;
        RECT 80.190 224.880 80.350 225.500 ;
        RECT 80.650 224.880 80.730 225.500 ;
        RECT 82.970 224.880 83.110 225.440 ;
        RECT 83.410 224.880 83.500 225.440 ;
        RECT 12.280 158.055 12.610 158.385 ;
        RECT 12.295 136.140 12.595 158.055 ;
        RECT 12.230 135.630 12.660 136.140 ;
        RECT 12.970 92.390 13.270 224.010 ;
        RECT 66.520 223.535 66.835 224.760 ;
        RECT 17.060 223.410 66.835 223.535 ;
        RECT 14.740 223.220 66.835 223.410 ;
        RECT 14.740 223.060 17.375 223.220 ;
        RECT 14.740 223.040 15.060 223.060 ;
        RECT 14.740 134.925 15.055 223.040 ;
        RECT 69.120 222.760 69.720 224.760 ;
        RECT 85.640 224.760 85.870 225.540 ;
        RECT 86.170 224.760 86.400 225.540 ;
        RECT 88.520 225.060 88.630 225.620 ;
        RECT 88.930 225.060 89.040 225.620 ;
        RECT 91.220 224.940 91.390 225.620 ;
        RECT 91.690 224.940 91.850 225.620 ;
        RECT 96.910 225.560 97.210 225.760 ;
        RECT 99.670 225.560 99.970 225.760 ;
        RECT 102.430 225.560 102.730 225.760 ;
        RECT 105.190 225.560 105.490 225.760 ;
        RECT 107.950 225.560 108.250 225.760 ;
        RECT 110.710 225.560 111.010 225.760 ;
        RECT 113.470 225.560 113.770 225.760 ;
        RECT 116.230 225.560 116.530 225.760 ;
        RECT 93.980 224.910 94.150 225.440 ;
        RECT 94.450 224.910 94.550 225.440 ;
        RECT 96.900 225.260 116.530 225.560 ;
        RECT 85.640 224.750 86.400 224.760 ;
        RECT 96.900 224.760 97.210 225.260 ;
        RECT 99.670 224.760 99.970 225.260 ;
        RECT 102.430 224.760 102.730 225.260 ;
        RECT 105.190 224.760 105.490 225.260 ;
        RECT 107.950 224.760 108.250 225.260 ;
        RECT 110.710 224.760 111.010 225.260 ;
        RECT 113.470 224.760 113.770 225.260 ;
        RECT 116.230 224.760 116.530 225.260 ;
        RECT 126.980 224.850 127.270 225.540 ;
        RECT 129.900 224.760 130.030 225.340 ;
        RECT 130.330 224.760 130.460 225.340 ;
        RECT 95.915 224.185 96.245 224.515 ;
        RECT 79.420 223.320 79.780 223.360 ;
        RECT 95.930 223.320 96.230 224.185 ;
        RECT 79.420 223.020 96.230 223.320 ;
        RECT 79.420 223.000 79.780 223.020 ;
        RECT 79.450 222.990 79.780 223.000 ;
        RECT 13.835 134.900 15.055 134.925 ;
        RECT 13.830 134.610 15.055 134.900 ;
        RECT 15.460 222.160 69.720 222.760 ;
        RECT 13.830 131.115 14.175 134.610 ;
        RECT 15.460 134.170 16.060 222.160 ;
        RECT 32.790 211.300 34.400 221.520 ;
        RECT 14.800 133.570 16.060 134.170 ;
        RECT 13.830 130.905 14.515 131.115 ;
        RECT 13.795 130.795 14.515 130.905 ;
        RECT 13.795 130.575 14.995 130.795 ;
        RECT 13.815 130.295 14.995 130.575 ;
        RECT 14.385 130.185 14.995 130.295 ;
        RECT 15.490 125.300 15.820 125.310 ;
        RECT 14.760 124.995 15.820 125.300 ;
        RECT 14.760 118.965 15.065 124.995 ;
        RECT 15.490 124.980 15.820 124.995 ;
        RECT 15.695 119.820 16.025 119.835 ;
        RECT 15.695 119.520 16.790 119.820 ;
        RECT 15.695 119.505 16.025 119.520 ;
        RECT 14.760 118.660 16.080 118.965 ;
        RECT 12.910 91.970 13.330 92.390 ;
        RECT 15.775 86.600 16.080 118.660 ;
        RECT 16.490 88.325 16.790 119.520 ;
        RECT 16.475 87.995 16.805 88.325 ;
        RECT 15.765 86.270 16.095 86.600 ;
        RECT 32.760 11.590 34.400 211.300 ;
        RECT 36.090 220.690 37.690 221.510 ;
        RECT 96.900 220.690 97.200 224.760 ;
        RECT 129.900 224.680 130.460 224.760 ;
        RECT 132.450 224.760 132.790 225.530 ;
        RECT 133.090 224.760 133.340 225.530 ;
        RECT 135.310 224.910 135.550 225.580 ;
        RECT 135.850 224.910 136.020 225.580 ;
        RECT 137.870 224.760 138.310 225.760 ;
        RECT 140.930 224.920 141.070 225.440 ;
        RECT 141.370 224.920 141.430 225.440 ;
        RECT 143.825 224.885 143.830 225.215 ;
        RECT 144.130 224.885 144.155 225.215 ;
        RECT 146.590 224.760 146.890 225.760 ;
        RECT 132.450 224.710 133.340 224.760 ;
        RECT 97.965 224.185 98.295 224.515 ;
        RECT 97.980 222.120 98.280 224.185 ;
        RECT 97.980 221.820 147.690 222.120 ;
        RECT 36.090 220.390 97.200 220.690 ;
        RECT 36.090 93.190 37.690 220.390 ;
        RECT 107.725 177.925 108.055 178.255 ;
        RECT 107.740 161.255 108.040 177.925 ;
        RECT 132.565 173.165 132.895 173.495 ;
        RECT 132.580 166.015 132.880 173.165 ;
        RECT 132.565 165.685 132.895 166.015 ;
        RECT 116.005 164.325 116.335 164.655 ;
        RECT 107.725 160.925 108.055 161.255 ;
        RECT 116.020 151.735 116.320 164.325 ;
        RECT 122.445 158.885 122.775 159.215 ;
        RECT 116.005 151.405 116.335 151.735 ;
        RECT 122.460 127.255 122.760 158.885 ;
        RECT 122.445 126.925 122.775 127.255 ;
        RECT 147.390 103.540 147.690 221.820 ;
        RECT 70.925 103.125 71.255 103.455 ;
        RECT 147.390 103.170 147.900 103.540 ;
        RECT 70.940 95.295 71.240 103.125 ;
        RECT 147.510 103.060 147.900 103.170 ;
        RECT 70.925 94.965 71.255 95.295 ;
        RECT 36.090 77.940 37.680 93.190 ;
        RECT 47.220 92.130 47.580 92.160 ;
        RECT 47.220 91.830 147.680 92.130 ;
        RECT 47.220 91.800 47.580 91.830 ;
        RECT 38.965 91.170 39.295 91.185 ;
        RECT 38.965 90.870 144.620 91.170 ;
        RECT 38.965 90.855 39.295 90.870 ;
        RECT 43.920 90.380 45.010 90.570 ;
        RECT 43.920 90.080 131.380 90.380 ;
        RECT 43.920 90.010 45.010 90.080 ;
        RECT 40.780 89.690 41.140 89.720 ;
        RECT 40.780 89.390 128.640 89.690 ;
        RECT 40.780 89.360 41.140 89.390 ;
        RECT 39.005 88.940 39.335 88.955 ;
        RECT 39.005 88.640 116.210 88.940 ;
        RECT 39.005 88.625 39.335 88.640 ;
        RECT 38.925 88.310 39.255 88.325 ;
        RECT 38.925 88.010 48.770 88.310 ;
        RECT 38.925 87.995 39.255 88.010 ;
        RECT 48.470 87.340 48.770 88.010 ;
        RECT 50.440 88.080 50.800 88.110 ;
        RECT 50.440 87.780 113.870 88.080 ;
        RECT 50.440 87.750 50.800 87.780 ;
        RECT 38.975 87.220 39.305 87.235 ;
        RECT 38.975 86.920 47.400 87.220 ;
        RECT 48.470 87.040 101.320 87.340 ;
        RECT 38.975 86.905 39.305 86.920 ;
        RECT 47.100 86.610 47.400 86.920 ;
        RECT 47.100 86.310 99.820 86.610 ;
        RECT 38.955 86.140 39.285 86.150 ;
        RECT 38.955 85.915 46.730 86.140 ;
        RECT 38.955 85.835 86.460 85.915 ;
        RECT 38.955 85.820 39.285 85.835 ;
        RECT 46.425 85.610 86.460 85.835 ;
        RECT 38.755 85.240 39.085 85.255 ;
        RECT 38.755 84.940 83.950 85.240 ;
        RECT 38.755 84.925 39.085 84.940 ;
        RECT 36.080 77.740 37.680 77.940 ;
        RECT 36.070 20.245 37.680 77.740 ;
        RECT 61.465 20.245 63.075 63.645 ;
        RECT 78.440 58.645 79.970 58.710 ;
        RECT 78.205 57.960 79.970 58.645 ;
        RECT 78.205 20.245 79.815 57.960 ;
        RECT 83.650 42.030 83.950 84.940 ;
        RECT 86.155 61.300 86.460 85.610 ;
        RECT 85.930 60.570 86.690 61.300 ;
        RECT 85.790 42.030 86.550 42.220 ;
        RECT 83.650 41.730 86.550 42.030 ;
        RECT 85.790 41.490 86.550 41.730 ;
        RECT 88.920 38.780 90.160 76.510 ;
        RECT 99.520 41.990 99.820 86.310 ;
        RECT 101.020 61.150 101.320 87.040 ;
        RECT 100.790 60.420 101.550 61.150 ;
        RECT 100.810 41.990 101.570 42.280 ;
        RECT 99.520 41.690 101.570 41.990 ;
        RECT 100.810 41.550 101.570 41.690 ;
        RECT 113.570 41.950 113.870 87.780 ;
        RECT 115.910 60.985 116.210 88.640 ;
        RECT 115.895 60.655 116.225 60.985 ;
        RECT 115.860 41.950 116.620 42.280 ;
        RECT 113.570 41.650 116.620 41.950 ;
        RECT 128.340 42.010 128.640 89.390 ;
        RECT 131.080 60.945 131.380 90.080 ;
        RECT 131.065 60.615 131.395 60.945 ;
        RECT 130.880 42.010 131.640 42.270 ;
        RECT 128.340 41.710 131.640 42.010 ;
        RECT 115.860 41.550 116.620 41.650 ;
        RECT 130.880 41.540 131.640 41.710 ;
        RECT 144.320 41.900 144.620 90.870 ;
        RECT 145.810 61.000 146.620 61.150 ;
        RECT 147.380 61.000 147.680 91.830 ;
        RECT 145.810 60.700 147.680 61.000 ;
        RECT 145.810 60.500 146.620 60.700 ;
        RECT 146.050 41.900 146.510 42.000 ;
        RECT 144.320 41.600 146.510 41.900 ;
        RECT 146.050 41.520 146.510 41.600 ;
        RECT 88.910 37.090 90.160 38.780 ;
        RECT 36.070 18.635 83.245 20.245 ;
        RECT 32.760 8.270 34.370 11.590 ;
        RECT 32.760 7.050 34.390 8.270 ;
        RECT 36.070 7.050 37.680 18.635 ;
        RECT 61.480 18.310 63.520 18.635 ;
        RECT 32.760 3.600 34.390 5.050 ;
        RECT 32.760 1.370 34.370 3.600 ;
        RECT 36.070 1.570 37.680 5.050 ;
        RECT 151.630 2.310 152.720 3.360 ;
        RECT 36.070 1.370 37.670 1.570 ;
        RECT 151.770 1.000 152.585 2.310 ;
        RECT 16.570 0.000 17.470 1.000 ;
        RECT 35.890 0.000 36.790 1.000 ;
        RECT 55.210 0.000 56.110 1.000 ;
        RECT 74.530 0.000 75.430 1.000 ;
        RECT 93.850 0.000 94.750 1.000 ;
        RECT 113.170 0.000 114.070 1.000 ;
        RECT 132.490 0.000 133.390 1.000 ;
        RECT 151.770 0.225 151.810 1.000 ;
  END
END top_dac_adc
END LIBRARY

