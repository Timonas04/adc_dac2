magic
tech sky130A
magscale 1 2
timestamp 1730493024
<< locali >>
rect 1416 1012 2480 1056
rect 1416 916 1472 1012
rect 2438 952 2480 1012
rect 1742 916 2480 952
rect 1416 904 2480 916
rect 1416 852 1742 904
rect 2458 852 2480 904
rect 1418 -962 2474 -920
rect 1418 -1078 1462 -962
rect 1764 -1012 2474 -962
rect 2436 -1078 2474 -1012
rect 1418 -1118 2474 -1078
<< viali >>
rect 1472 952 2438 1012
rect 1472 916 1742 952
rect 1462 -1012 1764 -962
rect 1462 -1078 2436 -1012
<< metal1 >>
rect 1416 1012 2480 1056
rect 1416 916 1472 1012
rect 2438 952 2480 1012
rect 1742 934 2480 952
rect 1742 918 1800 934
rect 1742 916 1766 918
rect 1416 852 1766 916
rect 1416 694 1486 852
rect 1916 848 2476 898
rect 1562 754 1626 804
rect 1416 -80 1566 694
rect 1620 678 1742 712
rect 1916 694 1948 848
rect 1976 814 2042 820
rect 1976 760 1982 814
rect 2036 760 2042 814
rect 2098 794 2140 848
rect 1976 754 2042 760
rect 2112 726 2140 794
rect 2168 814 2234 820
rect 2168 760 2174 814
rect 2228 760 2234 814
rect 2168 754 2234 760
rect 2328 752 2476 848
rect 2112 702 2170 726
rect 2112 696 2154 702
rect 2328 700 2362 752
rect 2398 736 2476 752
rect 1620 -30 1664 678
rect 1738 76 1742 678
rect 1738 -30 1744 76
rect 1620 -66 1744 -30
rect 1416 -82 1486 -80
rect 1516 -240 1652 -138
rect 1416 -270 1652 -240
rect 1416 -398 1450 -270
rect 1618 -398 1652 -270
rect 1416 -440 1652 -398
rect 1516 -538 1652 -440
rect 1416 -764 1564 -588
rect 1700 -590 1744 -66
rect 1800 -80 1858 -30
rect 2012 -78 2054 -42
rect 2210 -48 2244 -38
rect 2204 -78 2244 -48
rect 2330 -64 2362 700
rect 1800 -216 1852 -80
rect 1880 -114 1946 -108
rect 1880 -166 1888 -114
rect 1940 -166 1946 -114
rect 1880 -174 1946 -166
rect 2012 -210 2044 -78
rect 2072 -114 2138 -108
rect 2072 -168 2078 -114
rect 2132 -168 2138 -114
rect 2072 -174 2138 -168
rect 2204 -204 2236 -78
rect 2264 -114 2330 -108
rect 2264 -168 2270 -114
rect 2324 -168 2330 -114
rect 2264 -174 2330 -168
rect 1800 -218 1858 -216
rect 2012 -218 2054 -210
rect 2204 -218 2244 -204
rect 1800 -246 2244 -218
rect 2416 -228 2474 736
rect 1618 -646 1744 -590
rect 1798 -252 2244 -246
rect 1798 -348 2238 -252
rect 1798 -418 2292 -348
rect 1798 -436 2294 -418
rect 2322 -428 2522 -228
rect 1798 -626 1880 -436
rect 1974 -484 2040 -480
rect 1974 -540 1980 -484
rect 2034 -540 2040 -484
rect 1974 -546 2040 -540
rect 2070 -550 2104 -436
rect 2228 -438 2294 -436
rect 2166 -484 2232 -480
rect 2166 -540 2172 -484
rect 2226 -540 2232 -484
rect 2166 -546 2232 -540
rect 2264 -550 2294 -438
rect 2070 -596 2098 -550
rect 2074 -624 2098 -596
rect 2264 -622 2292 -550
rect 2416 -594 2474 -428
rect 1416 -808 1496 -764
rect 1618 -766 1738 -646
rect 1416 -916 1514 -808
rect 1556 -852 1626 -810
rect 1558 -864 1626 -852
rect 1878 -814 1944 -808
rect 1878 -870 1884 -814
rect 1938 -870 1944 -814
rect 1878 -874 1944 -870
rect 1974 -906 2002 -744
rect 2160 -778 2196 -732
rect 2330 -768 2474 -594
rect 2352 -778 2474 -768
rect 2164 -808 2196 -778
rect 2070 -814 2136 -808
rect 2070 -870 2076 -814
rect 2130 -870 2136 -814
rect 2070 -874 2136 -870
rect 2164 -906 2198 -808
rect 2262 -814 2328 -808
rect 2262 -870 2268 -814
rect 2322 -870 2328 -814
rect 2262 -874 2328 -870
rect 2356 -906 2474 -778
rect 1416 -920 1616 -916
rect 1416 -962 1776 -920
rect 1416 -1078 1462 -962
rect 1764 -1006 1776 -962
rect 1820 -946 2474 -906
rect 1820 -948 2386 -946
rect 1820 -978 2370 -948
rect 2422 -1006 2474 -998
rect 1764 -1012 2474 -1006
rect 2436 -1078 2474 -1012
rect 1416 -1116 2474 -1078
rect 1418 -1118 2474 -1116
<< via1 >>
rect 1982 760 2036 814
rect 2174 760 2228 814
rect 1664 -30 1738 678
rect 1450 -398 1618 -270
rect 1888 -166 1940 -114
rect 2078 -168 2132 -114
rect 2270 -168 2324 -114
rect 1980 -540 2034 -484
rect 2172 -540 2226 -484
rect 1884 -870 1938 -814
rect 2076 -870 2130 -814
rect 2268 -870 2322 -814
<< metal2 >>
rect 1708 814 2234 822
rect 1708 760 1982 814
rect 2036 760 2174 814
rect 2228 760 2234 814
rect 1708 752 2234 760
rect 1708 712 1762 752
rect 1626 678 1762 712
rect 1626 -30 1664 678
rect 1738 -30 1762 678
rect 1626 -64 1762 -30
rect 1704 -108 1760 -64
rect 1704 -114 2332 -108
rect 1704 -166 1888 -114
rect 1940 -166 2078 -114
rect 1704 -168 2078 -166
rect 2132 -168 2270 -114
rect 2324 -168 2332 -114
rect 1704 -172 2332 -168
rect 1880 -174 1946 -172
rect 2072 -174 2138 -172
rect 2264 -174 2330 -172
rect 1416 -270 1652 -238
rect 1416 -398 1450 -270
rect 1618 -370 1652 -270
rect 1618 -398 1784 -370
rect 1416 -438 1784 -398
rect 1416 -440 1652 -438
rect 1730 -480 1776 -438
rect 1730 -484 2232 -480
rect 1730 -540 1980 -484
rect 2034 -540 2172 -484
rect 2226 -540 2232 -484
rect 1730 -544 2232 -540
rect 1730 -808 1776 -544
rect 1974 -546 2040 -544
rect 2166 -546 2232 -544
rect 1730 -814 2330 -808
rect 1730 -870 1884 -814
rect 1938 -870 2076 -814
rect 2130 -870 2268 -814
rect 2322 -870 2330 -814
rect 1730 -876 2330 -870
use sky130_fd_pr__nfet_01v8_ATLS57  XM1
timestamp 1730493024
transform 1 0 2103 0 1 -678
box -407 -310 407 310
use sky130_fd_pr__pfet_01v8_XGSNAL  XM2
timestamp 1730493024
transform 1 0 2105 0 1 323
box -407 -619 407 619
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1730493024
transform 1 0 1591 0 1 -678
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGASDL  XM4
timestamp 1730493024
transform 1 0 1593 0 1 323
box -211 -619 211 619
<< labels >>
flabel metal1 1418 856 1618 1056 0 FreeSans 256 0 0 0 vdd
port 0 nsew
flabel metal1 1416 -1116 1616 -916 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 1416 -440 1616 -240 0 FreeSans 256 0 0 0 ctrl
port 1 nsew
flabel metal1 1896 -432 2096 -232 0 FreeSans 256 0 0 0 a
port 2 nsew
flabel metal1 2322 -428 2522 -228 0 FreeSans 256 0 0 0 b
port 3 nsew
<< end >>
